
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_NBIT32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_NBIT32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_0_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_0_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_0_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_14_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_14_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_14_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_13_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_13_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_13_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_12_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_12_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_12_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_11_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_11_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_11_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_10_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_10_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_10_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_9_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_9_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_9_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_8_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_8_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_8_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_7_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_7_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_7_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_6_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_6_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_6_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_5_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_5_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_5_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_4_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_4_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_4_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_3_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_3_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_3_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_2_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_2_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_2_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_1_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_GENERIC_NBIT64_1_DW01_add_0;

architecture SYN_rpl of RCA_GENERIC_NBIT64_1_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHMUL_NBIT32_DW01_inc_0 is

   port( A : in std_logic_vector (63 downto 0);  SUM : out std_logic_vector (63
         downto 0));

end BOOTHMUL_NBIT32_DW01_inc_0;

architecture SYN_rpl of BOOTHMUL_NBIT32_DW01_inc_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal SUM_62_port, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95
      , n96, n97, n98, n99, carry_31_port, carry_30_port, carry_29_port, 
      carry_28_port, carry_27_port, carry_26_port, carry_25_port, carry_24_port
      , carry_23_port, carry_22_port, carry_21_port, carry_20_port, 
      carry_19_port, carry_18_port, carry_17_port, carry_16_port, carry_15_port
      , carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, SUM_31_port, 
      n3, SUM_11_port, n5, SUM_12_port, n7, SUM_13_port, n9, SUM_14_port, n11, 
      SUM_15_port, n13, SUM_16_port, n15, SUM_17_port, n17, SUM_18_port, n19, 
      SUM_19_port, n21, SUM_20_port, n23, SUM_21_port, n25, SUM_22_port, n27, 
      SUM_23_port, n29, SUM_24_port, n31, SUM_25_port, n33, SUM_26_port, n35, 
      SUM_27_port, n37, SUM_28_port, n39, SUM_29_port, n41, SUM_30_port, n43, 
      SUM_9_port, n45, SUM_10_port, n47, SUM_7_port, n49, SUM_8_port, n51, 
      SUM_5_port, n53, SUM_6_port, n55, SUM_3_port, n57, SUM_4_port, n59, 
      SUM_1_port, n61, SUM_2_port, SUM_34_port, SUM_37_port, SUM_40_port, 
      SUM_45_port, SUM_51_port, n68, SUM_0_port : std_logic;

begin
   SUM <= ( SUM_51_port, SUM_51_port, SUM_51_port, SUM_51_port, SUM_51_port, 
      SUM_45_port, SUM_51_port, SUM_51_port, SUM_51_port, SUM_51_port, 
      SUM_40_port, SUM_34_port, SUM_51_port, SUM_45_port, SUM_45_port, 
      SUM_45_port, SUM_45_port, SUM_45_port, SUM_45_port, SUM_40_port, 
      SUM_37_port, SUM_40_port, SUM_40_port, SUM_40_port, SUM_37_port, 
      SUM_37_port, SUM_37_port, SUM_34_port, SUM_34_port, SUM_34_port, 
      SUM_51_port, SUM_51_port, SUM_31_port, SUM_30_port, SUM_29_port, 
      SUM_28_port, SUM_27_port, SUM_26_port, SUM_25_port, SUM_24_port, 
      SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, SUM_19_port, 
      SUM_18_port, SUM_17_port, SUM_16_port, SUM_15_port, SUM_14_port, 
      SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, SUM_6_port, SUM_5_port, SUM_4_port, SUM_3_port, 
      SUM_2_port, SUM_1_port, SUM_0_port );
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => n70);
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => n71);
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => n72);
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => n73);
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => n74);
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => n75);
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => n76);
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => n77);
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => n78);
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => n79);
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => n80);
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => n81);
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => n82);
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => n83);
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => n84);
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => n85);
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => n86);
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => n87);
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => n88);
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => n89);
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => n90);
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => n91);
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => n92);
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => n93);
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => n94);
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => n95);
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => n96);
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => n97);
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => n98);
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => n99)
                           ;
   U1 : BUF_X2 port map( A => SUM_62_port, Z => SUM_51_port);
   U2 : XNOR2_X1 port map( A => carry_31_port, B => A(62), ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => SUM_31_port);
   U4 : INV_X1 port map( A => n89, ZN => n3);
   U5 : INV_X1 port map( A => n3, ZN => SUM_11_port);
   U6 : INV_X1 port map( A => n88, ZN => n5);
   U7 : INV_X1 port map( A => n5, ZN => SUM_12_port);
   U8 : INV_X1 port map( A => n87, ZN => n7);
   U9 : INV_X1 port map( A => n7, ZN => SUM_13_port);
   U10 : INV_X1 port map( A => n86, ZN => n9);
   U11 : INV_X1 port map( A => n9, ZN => SUM_14_port);
   U12 : INV_X1 port map( A => n85, ZN => n11);
   U13 : INV_X1 port map( A => n11, ZN => SUM_15_port);
   U14 : INV_X1 port map( A => n84, ZN => n13);
   U15 : INV_X1 port map( A => n13, ZN => SUM_16_port);
   U16 : INV_X1 port map( A => n83, ZN => n15);
   U17 : INV_X1 port map( A => n15, ZN => SUM_17_port);
   U18 : INV_X1 port map( A => n82, ZN => n17);
   U19 : INV_X1 port map( A => n17, ZN => SUM_18_port);
   U20 : INV_X1 port map( A => n81, ZN => n19);
   U21 : INV_X1 port map( A => n19, ZN => SUM_19_port);
   U22 : INV_X1 port map( A => n80, ZN => n21);
   U23 : INV_X1 port map( A => n21, ZN => SUM_20_port);
   U24 : INV_X1 port map( A => n79, ZN => n23);
   U25 : INV_X1 port map( A => n23, ZN => SUM_21_port);
   U26 : INV_X1 port map( A => n78, ZN => n25);
   U27 : INV_X1 port map( A => n25, ZN => SUM_22_port);
   U28 : INV_X1 port map( A => n77, ZN => n27);
   U29 : INV_X1 port map( A => n27, ZN => SUM_23_port);
   U30 : INV_X1 port map( A => n76, ZN => n29);
   U31 : INV_X1 port map( A => n29, ZN => SUM_24_port);
   U32 : INV_X1 port map( A => n75, ZN => n31);
   U33 : INV_X1 port map( A => n31, ZN => SUM_25_port);
   U34 : INV_X1 port map( A => n74, ZN => n33);
   U35 : INV_X1 port map( A => n33, ZN => SUM_26_port);
   U36 : INV_X1 port map( A => n73, ZN => n35);
   U37 : INV_X1 port map( A => n35, ZN => SUM_27_port);
   U38 : INV_X1 port map( A => n72, ZN => n37);
   U39 : INV_X1 port map( A => n37, ZN => SUM_28_port);
   U40 : INV_X1 port map( A => n71, ZN => n39);
   U41 : INV_X1 port map( A => n39, ZN => SUM_29_port);
   U42 : INV_X1 port map( A => n70, ZN => n41);
   U43 : INV_X1 port map( A => n41, ZN => SUM_30_port);
   U44 : INV_X1 port map( A => n91, ZN => n43);
   U45 : INV_X1 port map( A => n43, ZN => SUM_9_port);
   U46 : INV_X1 port map( A => n90, ZN => n45);
   U47 : INV_X1 port map( A => n45, ZN => SUM_10_port);
   U48 : INV_X1 port map( A => n93, ZN => n47);
   U49 : INV_X1 port map( A => n47, ZN => SUM_7_port);
   U50 : INV_X1 port map( A => n92, ZN => n49);
   U51 : INV_X1 port map( A => n49, ZN => SUM_8_port);
   U52 : INV_X1 port map( A => n95, ZN => n51);
   U53 : INV_X1 port map( A => n51, ZN => SUM_5_port);
   U54 : INV_X1 port map( A => n94, ZN => n53);
   U55 : INV_X1 port map( A => n53, ZN => SUM_6_port);
   U56 : INV_X1 port map( A => n97, ZN => n55);
   U57 : INV_X1 port map( A => n55, ZN => SUM_3_port);
   U58 : INV_X1 port map( A => n96, ZN => n57);
   U59 : INV_X1 port map( A => n57, ZN => SUM_4_port);
   U60 : INV_X1 port map( A => n99, ZN => n59);
   U61 : INV_X1 port map( A => n59, ZN => SUM_1_port);
   U62 : INV_X1 port map( A => n98, ZN => n61);
   U63 : INV_X1 port map( A => n61, ZN => SUM_2_port);
   U64 : BUF_X4 port map( A => SUM_62_port, Z => SUM_45_port);
   U65 : INV_X1 port map( A => A(0), ZN => SUM_0_port);
   U66 : CLKBUF_X3 port map( A => SUM_62_port, Z => SUM_34_port);
   U67 : CLKBUF_X3 port map( A => SUM_62_port, Z => SUM_37_port);
   U68 : CLKBUF_X3 port map( A => SUM_62_port, Z => SUM_40_port);
   U69 : INV_X1 port map( A => A(62), ZN => n68);
   U70 : NOR2_X1 port map( A1 => carry_31_port, A2 => n68, ZN => SUM_62_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_63 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_63;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_63 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U11 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U12 : MUX2_X1 port map( A => A(63), B => B(63), S => n1, Z => Y(63));
   U13 : MUX2_X1 port map( A => A(62), B => B(62), S => n1, Z => Y(62));
   U14 : MUX2_X1 port map( A => A(61), B => B(61), S => n1, Z => Y(61));
   U15 : MUX2_X1 port map( A => A(60), B => B(60), S => n1, Z => Y(60));
   U16 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U17 : MUX2_X1 port map( A => A(59), B => B(59), S => n1, Z => Y(59));
   U18 : MUX2_X1 port map( A => A(58), B => B(58), S => n1, Z => Y(58));
   U19 : MUX2_X1 port map( A => A(57), B => B(57), S => n2, Z => Y(57));
   U20 : MUX2_X1 port map( A => A(56), B => B(56), S => n2, Z => Y(56));
   U21 : MUX2_X1 port map( A => A(55), B => B(55), S => n2, Z => Y(55));
   U22 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U25 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(4), B => B(4), S => n2, Z => Y(4));
   U28 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U29 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U30 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U31 : MUX2_X1 port map( A => A(46), B => B(46), S => n3, Z => Y(46));
   U32 : MUX2_X1 port map( A => A(45), B => B(45), S => n3, Z => Y(45));
   U33 : MUX2_X1 port map( A => A(44), B => B(44), S => n3, Z => Y(44));
   U34 : MUX2_X1 port map( A => A(43), B => B(43), S => n3, Z => Y(43));
   U35 : MUX2_X1 port map( A => A(42), B => B(42), S => n3, Z => Y(42));
   U36 : MUX2_X1 port map( A => A(41), B => B(41), S => n3, Z => Y(41));
   U37 : MUX2_X1 port map( A => A(40), B => B(40), S => n3, Z => Y(40));
   U38 : MUX2_X1 port map( A => A(3), B => B(3), S => n3, Z => Y(3));
   U39 : MUX2_X1 port map( A => A(39), B => B(39), S => n3, Z => Y(39));
   U40 : MUX2_X1 port map( A => A(38), B => B(38), S => n3, Z => Y(38));
   U41 : MUX2_X1 port map( A => A(37), B => B(37), S => n3, Z => Y(37));
   U42 : MUX2_X1 port map( A => A(36), B => B(36), S => n3, Z => Y(36));
   U43 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U44 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U45 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U46 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U47 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U48 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U49 : MUX2_X1 port map( A => A(2), B => B(2), S => n4, Z => Y(2));
   U50 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U51 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U52 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U53 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U54 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U55 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U56 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U57 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U58 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U59 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U60 : MUX2_X1 port map( A => A(1), B => B(1), S => n5, Z => Y(1));
   U61 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U62 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U63 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U64 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U65 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U66 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U67 : MUX2_X1 port map( A => A(13), B => B(13), S => n6, Z => Y(13));
   U68 : MUX2_X1 port map( A => A(12), B => B(12), S => n6, Z => Y(12));
   U69 : MUX2_X1 port map( A => A(11), B => B(11), S => n6, Z => Y(11));
   U70 : MUX2_X1 port map( A => A(10), B => B(10), S => n6, Z => Y(10));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_62 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_62;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_62 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U3 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U4 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U5 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U6 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U7 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U8 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U9 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U10 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U11 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U12 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U13 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U14 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U15 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U16 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U17 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U18 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U19 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U22 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U23 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U24 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U25 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U26 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U27 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U28 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U29 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U30 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U31 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U32 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U33 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U34 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U35 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U36 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U37 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U38 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U39 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U40 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U41 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U42 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U43 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U44 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U45 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U46 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U47 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U48 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U49 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U50 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U51 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U52 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U53 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U54 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U55 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U56 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U57 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U58 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U59 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U60 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U61 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U62 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U63 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U64 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_61 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_61;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_61 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_60 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_60;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_60 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(33), B => B(33), S => n1, Z => Y(33));
   U10 : MUX2_X1 port map( A => A(34), B => B(34), S => n1, Z => Y(34));
   U11 : MUX2_X1 port map( A => A(35), B => B(35), S => n1, Z => Y(35));
   U12 : MUX2_X1 port map( A => A(36), B => B(36), S => n1, Z => Y(36));
   U13 : MUX2_X1 port map( A => A(37), B => B(37), S => n1, Z => Y(37));
   U14 : MUX2_X1 port map( A => A(38), B => B(38), S => n1, Z => Y(38));
   U15 : MUX2_X1 port map( A => A(39), B => B(39), S => n1, Z => Y(39));
   U16 : MUX2_X1 port map( A => A(40), B => B(40), S => n1, Z => Y(40));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(32), B => B(32), S => n3, Z => Y(32));
   U41 : MUX2_X1 port map( A => A(31), B => B(31), S => n3, Z => Y(31));
   U42 : MUX2_X1 port map( A => A(30), B => B(30), S => n3, Z => Y(30));
   U43 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U44 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U45 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U46 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U47 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U48 : MUX2_X1 port map( A => A(24), B => B(24), S => n4, Z => Y(24));
   U49 : MUX2_X1 port map( A => A(23), B => B(23), S => n4, Z => Y(23));
   U50 : MUX2_X1 port map( A => A(22), B => B(22), S => n4, Z => Y(22));
   U51 : MUX2_X1 port map( A => A(21), B => B(21), S => n4, Z => Y(21));
   U52 : MUX2_X1 port map( A => A(20), B => B(20), S => n4, Z => Y(20));
   U53 : MUX2_X1 port map( A => A(19), B => B(19), S => n4, Z => Y(19));
   U54 : MUX2_X1 port map( A => A(18), B => B(18), S => n4, Z => Y(18));
   U55 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U56 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U57 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U58 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U59 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U60 : MUX2_X1 port map( A => A(12), B => B(12), S => n5, Z => Y(12));
   U61 : MUX2_X1 port map( A => A(11), B => B(11), S => n5, Z => Y(11));
   U62 : MUX2_X1 port map( A => A(10), B => B(10), S => n5, Z => Y(10));
   U63 : MUX2_X1 port map( A => A(9), B => B(9), S => n5, Z => Y(9));
   U64 : MUX2_X1 port map( A => A(8), B => B(8), S => n5, Z => Y(8));
   U65 : MUX2_X1 port map( A => A(7), B => B(7), S => n5, Z => Y(7));
   U66 : MUX2_X1 port map( A => A(6), B => B(6), S => n5, Z => Y(6));
   U67 : MUX2_X1 port map( A => A(5), B => B(5), S => n6, Z => Y(5));
   U68 : MUX2_X1 port map( A => A(4), B => B(4), S => n6, Z => Y(4));
   U69 : MUX2_X1 port map( A => A(3), B => B(3), S => n6, Z => Y(3));
   U70 : MUX2_X1 port map( A => A(2), B => B(2), S => n6, Z => Y(2));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_59 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_59;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_59 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(34), B => B(34), S => n1, Z => Y(34));
   U11 : MUX2_X1 port map( A => A(35), B => B(35), S => n1, Z => Y(35));
   U12 : MUX2_X1 port map( A => A(36), B => B(36), S => n1, Z => Y(36));
   U13 : MUX2_X1 port map( A => A(37), B => B(37), S => n1, Z => Y(37));
   U14 : MUX2_X1 port map( A => A(38), B => B(38), S => n1, Z => Y(38));
   U15 : MUX2_X1 port map( A => A(39), B => B(39), S => n1, Z => Y(39));
   U16 : MUX2_X1 port map( A => A(40), B => B(40), S => n1, Z => Y(40));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(33), B => B(33), S => n3, Z => Y(33));
   U41 : MUX2_X1 port map( A => A(32), B => B(32), S => n3, Z => Y(32));
   U42 : MUX2_X1 port map( A => A(31), B => B(31), S => n3, Z => Y(31));
   U43 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U44 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U45 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U46 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U47 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U48 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U49 : MUX2_X1 port map( A => A(24), B => B(24), S => n4, Z => Y(24));
   U50 : MUX2_X1 port map( A => A(23), B => B(23), S => n4, Z => Y(23));
   U51 : MUX2_X1 port map( A => A(22), B => B(22), S => n4, Z => Y(22));
   U52 : MUX2_X1 port map( A => A(21), B => B(21), S => n4, Z => Y(21));
   U53 : MUX2_X1 port map( A => A(20), B => B(20), S => n4, Z => Y(20));
   U54 : MUX2_X1 port map( A => A(19), B => B(19), S => n4, Z => Y(19));
   U55 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U56 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U57 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U58 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U59 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U60 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U61 : MUX2_X1 port map( A => A(12), B => B(12), S => n5, Z => Y(12));
   U62 : MUX2_X1 port map( A => A(11), B => B(11), S => n5, Z => Y(11));
   U63 : MUX2_X1 port map( A => A(10), B => B(10), S => n5, Z => Y(10));
   U64 : MUX2_X1 port map( A => A(9), B => B(9), S => n5, Z => Y(9));
   U65 : MUX2_X1 port map( A => A(8), B => B(8), S => n5, Z => Y(8));
   U66 : MUX2_X1 port map( A => A(7), B => B(7), S => n5, Z => Y(7));
   U67 : MUX2_X1 port map( A => A(6), B => B(6), S => n6, Z => Y(6));
   U68 : MUX2_X1 port map( A => A(5), B => B(5), S => n6, Z => Y(5));
   U69 : MUX2_X1 port map( A => A(4), B => B(4), S => n6, Z => Y(4));
   U70 : MUX2_X1 port map( A => A(3), B => B(3), S => n6, Z => Y(3));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_58 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_58;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_58 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U5 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U6 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U7 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U8 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U9 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U10 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U11 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U12 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U13 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U14 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U15 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U16 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U17 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U18 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U19 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U36 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U37 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U38 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U39 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U40 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U41 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U42 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U43 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U44 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U45 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U46 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U47 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U48 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U49 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U50 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U51 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U52 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U53 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U54 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U55 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U56 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U57 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U58 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U59 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U60 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U61 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U62 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U63 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U64 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_57 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_57;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_57 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_56 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_56;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_56 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(35), B => B(35), S => n1, Z => Y(35));
   U12 : MUX2_X1 port map( A => A(36), B => B(36), S => n1, Z => Y(36));
   U13 : MUX2_X1 port map( A => A(37), B => B(37), S => n1, Z => Y(37));
   U14 : MUX2_X1 port map( A => A(38), B => B(38), S => n1, Z => Y(38));
   U15 : MUX2_X1 port map( A => A(39), B => B(39), S => n1, Z => Y(39));
   U16 : MUX2_X1 port map( A => A(40), B => B(40), S => n1, Z => Y(40));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(34), B => B(34), S => n3, Z => Y(34));
   U41 : MUX2_X1 port map( A => A(33), B => B(33), S => n3, Z => Y(33));
   U42 : MUX2_X1 port map( A => A(32), B => B(32), S => n3, Z => Y(32));
   U43 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U44 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U45 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U46 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U47 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U48 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U49 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U50 : MUX2_X1 port map( A => A(24), B => B(24), S => n4, Z => Y(24));
   U51 : MUX2_X1 port map( A => A(23), B => B(23), S => n4, Z => Y(23));
   U52 : MUX2_X1 port map( A => A(22), B => B(22), S => n4, Z => Y(22));
   U53 : MUX2_X1 port map( A => A(21), B => B(21), S => n4, Z => Y(21));
   U54 : MUX2_X1 port map( A => A(20), B => B(20), S => n4, Z => Y(20));
   U55 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U56 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U57 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U58 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U59 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U60 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U61 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U62 : MUX2_X1 port map( A => A(12), B => B(12), S => n5, Z => Y(12));
   U63 : MUX2_X1 port map( A => A(11), B => B(11), S => n5, Z => Y(11));
   U64 : MUX2_X1 port map( A => A(10), B => B(10), S => n5, Z => Y(10));
   U65 : MUX2_X1 port map( A => A(9), B => B(9), S => n5, Z => Y(9));
   U66 : MUX2_X1 port map( A => A(8), B => B(8), S => n5, Z => Y(8));
   U67 : MUX2_X1 port map( A => A(7), B => B(7), S => n6, Z => Y(7));
   U68 : MUX2_X1 port map( A => A(6), B => B(6), S => n6, Z => Y(6));
   U69 : MUX2_X1 port map( A => A(5), B => B(5), S => n6, Z => Y(5));
   U70 : MUX2_X1 port map( A => A(4), B => B(4), S => n6, Z => Y(4));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_55 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_55;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_55 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(36), B => B(36), S => n1, Z => Y(36));
   U13 : MUX2_X1 port map( A => A(37), B => B(37), S => n1, Z => Y(37));
   U14 : MUX2_X1 port map( A => A(38), B => B(38), S => n1, Z => Y(38));
   U15 : MUX2_X1 port map( A => A(39), B => B(39), S => n1, Z => Y(39));
   U16 : MUX2_X1 port map( A => A(40), B => B(40), S => n1, Z => Y(40));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(35), B => B(35), S => n3, Z => Y(35));
   U41 : MUX2_X1 port map( A => A(34), B => B(34), S => n3, Z => Y(34));
   U42 : MUX2_X1 port map( A => A(33), B => B(33), S => n3, Z => Y(33));
   U43 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U44 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U45 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U46 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U47 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U48 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U49 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U50 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U51 : MUX2_X1 port map( A => A(24), B => B(24), S => n4, Z => Y(24));
   U52 : MUX2_X1 port map( A => A(23), B => B(23), S => n4, Z => Y(23));
   U53 : MUX2_X1 port map( A => A(22), B => B(22), S => n4, Z => Y(22));
   U54 : MUX2_X1 port map( A => A(21), B => B(21), S => n4, Z => Y(21));
   U55 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U56 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U57 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U58 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U59 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U60 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U61 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U62 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U63 : MUX2_X1 port map( A => A(12), B => B(12), S => n5, Z => Y(12));
   U64 : MUX2_X1 port map( A => A(11), B => B(11), S => n5, Z => Y(11));
   U65 : MUX2_X1 port map( A => A(10), B => B(10), S => n5, Z => Y(10));
   U66 : MUX2_X1 port map( A => A(9), B => B(9), S => n5, Z => Y(9));
   U67 : MUX2_X1 port map( A => A(8), B => B(8), S => n6, Z => Y(8));
   U68 : MUX2_X1 port map( A => A(7), B => B(7), S => n6, Z => Y(7));
   U69 : MUX2_X1 port map( A => A(6), B => B(6), S => n6, Z => Y(6));
   U70 : MUX2_X1 port map( A => A(5), B => B(5), S => n6, Z => Y(5));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_54 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_54;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_54 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U7 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U8 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U9 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U10 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U11 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U12 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U13 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U14 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U15 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U16 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U17 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U18 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U19 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U37 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U38 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U39 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U40 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U41 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U42 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U43 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U44 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U45 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U46 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U47 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U48 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U49 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U50 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U51 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U52 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U53 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U54 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U55 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U56 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U57 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U58 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U59 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U60 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U61 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U62 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U63 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U64 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_53 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_53;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_53 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_52 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_52;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_52 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(37), B => B(37), S => n1, Z => Y(37));
   U14 : MUX2_X1 port map( A => A(38), B => B(38), S => n1, Z => Y(38));
   U15 : MUX2_X1 port map( A => A(39), B => B(39), S => n1, Z => Y(39));
   U16 : MUX2_X1 port map( A => A(40), B => B(40), S => n1, Z => Y(40));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(36), B => B(36), S => n3, Z => Y(36));
   U41 : MUX2_X1 port map( A => A(35), B => B(35), S => n3, Z => Y(35));
   U42 : MUX2_X1 port map( A => A(34), B => B(34), S => n3, Z => Y(34));
   U43 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U44 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U45 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U46 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U47 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U48 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U49 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U50 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U51 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U52 : MUX2_X1 port map( A => A(24), B => B(24), S => n4, Z => Y(24));
   U53 : MUX2_X1 port map( A => A(23), B => B(23), S => n4, Z => Y(23));
   U54 : MUX2_X1 port map( A => A(22), B => B(22), S => n4, Z => Y(22));
   U55 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U56 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U57 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U58 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U59 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U60 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U61 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U62 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U63 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U64 : MUX2_X1 port map( A => A(12), B => B(12), S => n5, Z => Y(12));
   U65 : MUX2_X1 port map( A => A(11), B => B(11), S => n5, Z => Y(11));
   U66 : MUX2_X1 port map( A => A(10), B => B(10), S => n5, Z => Y(10));
   U67 : MUX2_X1 port map( A => A(9), B => B(9), S => n6, Z => Y(9));
   U68 : MUX2_X1 port map( A => A(8), B => B(8), S => n6, Z => Y(8));
   U69 : MUX2_X1 port map( A => A(7), B => B(7), S => n6, Z => Y(7));
   U70 : MUX2_X1 port map( A => A(6), B => B(6), S => n6, Z => Y(6));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_51 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_51;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_51 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(38), B => B(38), S => n1, Z => Y(38));
   U15 : MUX2_X1 port map( A => A(39), B => B(39), S => n1, Z => Y(39));
   U16 : MUX2_X1 port map( A => A(40), B => B(40), S => n1, Z => Y(40));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(37), B => B(37), S => n3, Z => Y(37));
   U41 : MUX2_X1 port map( A => A(36), B => B(36), S => n3, Z => Y(36));
   U42 : MUX2_X1 port map( A => A(35), B => B(35), S => n3, Z => Y(35));
   U43 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U44 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U45 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U46 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U47 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U48 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U49 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U50 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U51 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U52 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U53 : MUX2_X1 port map( A => A(24), B => B(24), S => n4, Z => Y(24));
   U54 : MUX2_X1 port map( A => A(23), B => B(23), S => n4, Z => Y(23));
   U55 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U56 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U57 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U58 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U59 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U60 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U61 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U62 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U63 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U64 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U65 : MUX2_X1 port map( A => A(12), B => B(12), S => n5, Z => Y(12));
   U66 : MUX2_X1 port map( A => A(11), B => B(11), S => n5, Z => Y(11));
   U67 : MUX2_X1 port map( A => A(10), B => B(10), S => n6, Z => Y(10));
   U68 : MUX2_X1 port map( A => A(9), B => B(9), S => n6, Z => Y(9));
   U69 : MUX2_X1 port map( A => A(8), B => B(8), S => n6, Z => Y(8));
   U70 : MUX2_X1 port map( A => A(7), B => B(7), S => n6, Z => Y(7));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_50 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_50;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_50 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U9 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U10 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U11 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U12 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U13 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U14 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U15 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U16 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U17 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U18 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U19 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U35 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U38 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U39 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U40 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U41 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U42 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U43 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U44 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U45 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U46 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U47 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U48 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U49 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U50 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U51 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U52 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U53 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U54 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U55 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U56 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U57 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U58 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U59 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U60 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U61 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U62 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U63 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U64 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_49 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_49;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_49 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_48 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_48;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_48 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(39), B => B(39), S => n1, Z => Y(39));
   U16 : MUX2_X1 port map( A => A(40), B => B(40), S => n1, Z => Y(40));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(38), B => B(38), S => n3, Z => Y(38));
   U41 : MUX2_X1 port map( A => A(37), B => B(37), S => n3, Z => Y(37));
   U42 : MUX2_X1 port map( A => A(36), B => B(36), S => n3, Z => Y(36));
   U43 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U44 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U45 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U46 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U47 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U48 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U49 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U50 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U51 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U52 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U53 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U54 : MUX2_X1 port map( A => A(24), B => B(24), S => n4, Z => Y(24));
   U55 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U56 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U57 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U58 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U59 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U60 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U61 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U62 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U63 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U64 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U65 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U66 : MUX2_X1 port map( A => A(12), B => B(12), S => n5, Z => Y(12));
   U67 : MUX2_X1 port map( A => A(11), B => B(11), S => n6, Z => Y(11));
   U68 : MUX2_X1 port map( A => A(10), B => B(10), S => n6, Z => Y(10));
   U69 : MUX2_X1 port map( A => A(9), B => B(9), S => n6, Z => Y(9));
   U70 : MUX2_X1 port map( A => A(8), B => B(8), S => n6, Z => Y(8));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_47 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_47;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_47 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(40), B => B(40), S => n1, Z => Y(40));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => n3, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(38), B => B(38), S => n3, Z => Y(38));
   U42 : MUX2_X1 port map( A => A(37), B => B(37), S => n3, Z => Y(37));
   U43 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U44 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U45 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U46 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U47 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U48 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U49 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U50 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U51 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U52 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U53 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U54 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U55 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U56 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U57 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U58 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U59 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U60 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U61 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U62 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U63 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U64 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U65 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U66 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U67 : MUX2_X1 port map( A => A(12), B => B(12), S => n6, Z => Y(12));
   U68 : MUX2_X1 port map( A => A(11), B => B(11), S => n6, Z => Y(11));
   U69 : MUX2_X1 port map( A => A(10), B => B(10), S => n6, Z => Y(10));
   U70 : MUX2_X1 port map( A => A(9), B => B(9), S => n6, Z => Y(9));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_46 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_46;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_46 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U11 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U12 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U13 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U14 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U15 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U16 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U17 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U18 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U19 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U35 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U36 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U39 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U40 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U41 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U42 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U43 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U44 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U45 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U46 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U47 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U48 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U49 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U50 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U51 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U52 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U53 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U54 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U55 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U56 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U57 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U58 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U59 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U60 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U61 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U62 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U63 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U64 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_45 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_45;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_45 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_44 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_44;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_44 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(41), B => B(41), S => n1, Z => Y(41));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(40), B => B(40), S => n3, Z => Y(40));
   U41 : MUX2_X1 port map( A => A(39), B => B(39), S => n3, Z => Y(39));
   U42 : MUX2_X1 port map( A => A(38), B => B(38), S => n3, Z => Y(38));
   U43 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U44 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U45 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U46 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U47 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U48 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U49 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U50 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U51 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U52 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U53 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U54 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U55 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U56 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U57 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U58 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U59 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U60 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U61 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U62 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U63 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U64 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U65 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U66 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U67 : MUX2_X1 port map( A => A(13), B => B(13), S => n6, Z => Y(13));
   U68 : MUX2_X1 port map( A => A(12), B => B(12), S => n6, Z => Y(12));
   U69 : MUX2_X1 port map( A => A(11), B => B(11), S => n6, Z => Y(11));
   U70 : MUX2_X1 port map( A => A(10), B => B(10), S => n6, Z => Y(10));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_43 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_43;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_43 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(42), B => B(42), S => n1, Z => Y(42));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(41), B => B(41), S => n3, Z => Y(41));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => n3, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(39), B => B(39), S => n3, Z => Y(39));
   U43 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U44 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U45 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U46 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U47 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U48 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U49 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U50 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U51 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U52 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U53 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U54 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U55 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U56 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U57 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U58 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U59 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U60 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U61 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U62 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U63 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U64 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U65 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U66 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U67 : MUX2_X1 port map( A => A(14), B => B(14), S => n6, Z => Y(14));
   U68 : MUX2_X1 port map( A => A(13), B => B(13), S => n6, Z => Y(13));
   U69 : MUX2_X1 port map( A => A(12), B => B(12), S => n6, Z => Y(12));
   U70 : MUX2_X1 port map( A => A(11), B => B(11), S => n6, Z => Y(11));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_42 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_42;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_42 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U13 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U14 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U15 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U16 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U17 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U18 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U19 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U35 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U36 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U37 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U40 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U41 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U42 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U43 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U44 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U45 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U46 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U47 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U48 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U49 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U50 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U51 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U52 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U53 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U54 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U55 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U56 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U57 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U58 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U59 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U60 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U61 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U62 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U63 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U64 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_41 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_41;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_41 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_40 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_40;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_40 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(43), B => B(43), S => n2, Z => Y(43));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(42), B => B(42), S => n3, Z => Y(42));
   U41 : MUX2_X1 port map( A => A(41), B => B(41), S => n3, Z => Y(41));
   U42 : MUX2_X1 port map( A => A(40), B => B(40), S => n3, Z => Y(40));
   U43 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U44 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U45 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U46 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U47 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U48 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U49 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U50 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U51 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U52 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U53 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U54 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U55 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U56 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U57 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U58 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U59 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U60 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U61 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U62 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U63 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U64 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U65 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U66 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U67 : MUX2_X1 port map( A => A(15), B => B(15), S => n6, Z => Y(15));
   U68 : MUX2_X1 port map( A => A(14), B => B(14), S => n6, Z => Y(14));
   U69 : MUX2_X1 port map( A => A(13), B => B(13), S => n6, Z => Y(13));
   U70 : MUX2_X1 port map( A => A(12), B => B(12), S => n6, Z => Y(12));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_39 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_39;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_39 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(44), B => B(44), S => n2, Z => Y(44));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(43), B => B(43), S => n3, Z => Y(43));
   U41 : MUX2_X1 port map( A => A(42), B => B(42), S => n3, Z => Y(42));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => n3, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U44 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U45 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U46 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U47 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U48 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U49 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U50 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U51 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U52 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U53 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U54 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U55 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U56 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U57 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U58 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U59 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U60 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U61 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U62 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U63 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U64 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U65 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U66 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U67 : MUX2_X1 port map( A => A(16), B => B(16), S => n6, Z => Y(16));
   U68 : MUX2_X1 port map( A => A(15), B => B(15), S => n6, Z => Y(15));
   U69 : MUX2_X1 port map( A => A(14), B => B(14), S => n6, Z => Y(14));
   U70 : MUX2_X1 port map( A => A(13), B => B(13), S => n6, Z => Y(13));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_38 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_38;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_38 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U15 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U16 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U17 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U18 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U19 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U35 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U36 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U37 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U38 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U41 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U42 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U43 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U44 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U45 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U46 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U47 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U48 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U49 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U50 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U51 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U52 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U53 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U54 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U55 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U56 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U57 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U58 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U59 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U60 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U61 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U62 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U63 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U64 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_37 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_37;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_37 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_36 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_36;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_36 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(45), B => B(45), S => n2, Z => Y(45));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(44), B => B(44), S => n3, Z => Y(44));
   U41 : MUX2_X1 port map( A => A(43), B => B(43), S => n3, Z => Y(43));
   U42 : MUX2_X1 port map( A => A(42), B => B(42), S => n3, Z => Y(42));
   U43 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U44 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U45 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U46 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U47 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U48 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U49 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U50 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U51 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U52 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U53 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U54 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U55 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U56 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U57 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U58 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U59 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U60 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U61 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U62 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U63 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U64 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U65 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U66 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U67 : MUX2_X1 port map( A => A(17), B => B(17), S => n6, Z => Y(17));
   U68 : MUX2_X1 port map( A => A(16), B => B(16), S => n6, Z => Y(16));
   U69 : MUX2_X1 port map( A => A(15), B => B(15), S => n6, Z => Y(15));
   U70 : MUX2_X1 port map( A => A(14), B => B(14), S => n6, Z => Y(14));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_35 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_35;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_35 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(45), B => B(45), S => n3, Z => Y(45));
   U41 : MUX2_X1 port map( A => A(44), B => B(44), S => n3, Z => Y(44));
   U42 : MUX2_X1 port map( A => A(43), B => B(43), S => n3, Z => Y(43));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U45 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U46 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U47 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U48 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U49 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U50 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U51 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U52 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U53 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U54 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U55 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U56 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U57 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U58 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U59 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U60 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U61 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U62 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U63 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U64 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U65 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U66 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U67 : MUX2_X1 port map( A => A(18), B => B(18), S => n6, Z => Y(18));
   U68 : MUX2_X1 port map( A => A(17), B => B(17), S => n6, Z => Y(17));
   U69 : MUX2_X1 port map( A => A(16), B => B(16), S => n6, Z => Y(16));
   U70 : MUX2_X1 port map( A => A(15), B => B(15), S => n6, Z => Y(15));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_34 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_34;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_34 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U17 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U18 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U19 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U35 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U36 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U37 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U38 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U39 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U42 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U43 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U44 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U45 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U46 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U47 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U48 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U49 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U50 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U51 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U52 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U53 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U54 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U55 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U56 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U57 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U58 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U59 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U60 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U61 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U62 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U63 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U64 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_33 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_33;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_33 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_32 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_32;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(46), B => B(46), S => n3, Z => Y(46));
   U41 : MUX2_X1 port map( A => A(45), B => B(45), S => n3, Z => Y(45));
   U42 : MUX2_X1 port map( A => A(44), B => B(44), S => n3, Z => Y(44));
   U43 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U44 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U45 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U46 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U47 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U48 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U49 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U50 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U51 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U52 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U53 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U54 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U55 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U56 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U57 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U58 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U59 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U60 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U61 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U62 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U63 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U64 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U65 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U66 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U67 : MUX2_X1 port map( A => A(19), B => B(19), S => n6, Z => Y(19));
   U68 : MUX2_X1 port map( A => A(18), B => B(18), S => n6, Z => Y(18));
   U69 : MUX2_X1 port map( A => A(17), B => B(17), S => n6, Z => Y(17));
   U70 : MUX2_X1 port map( A => A(16), B => B(16), S => n6, Z => Y(16));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_31 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_31;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_31 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(47), B => B(47), S => n3, Z => Y(47));
   U41 : MUX2_X1 port map( A => A(46), B => B(46), S => n3, Z => Y(46));
   U42 : MUX2_X1 port map( A => A(45), B => B(45), S => n3, Z => Y(45));
   U43 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U46 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U47 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U48 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U49 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U50 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U51 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U52 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U53 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U54 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U55 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U56 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U57 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U58 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U59 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U60 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U61 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U62 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U63 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U64 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U65 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U66 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U67 : MUX2_X1 port map( A => A(20), B => B(20), S => n6, Z => Y(20));
   U68 : MUX2_X1 port map( A => A(19), B => B(19), S => n6, Z => Y(19));
   U69 : MUX2_X1 port map( A => A(18), B => B(18), S => n6, Z => Y(18));
   U70 : MUX2_X1 port map( A => A(17), B => B(17), S => n6, Z => Y(17));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_30 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_30;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_30 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U19 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U35 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U36 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U37 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U38 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U39 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U40 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U43 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U44 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U45 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U46 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U47 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U48 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U49 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U50 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U51 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U52 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U53 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U54 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U55 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U56 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U57 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U58 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U59 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U60 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U61 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U62 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U63 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U64 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_29 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_29;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_29 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_28 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_28;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_28 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(48), B => B(48), S => n3, Z => Y(48));
   U41 : MUX2_X1 port map( A => A(47), B => B(47), S => n3, Z => Y(47));
   U42 : MUX2_X1 port map( A => A(46), B => B(46), S => n3, Z => Y(46));
   U43 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U44 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U45 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U46 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U47 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U48 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U49 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U50 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U51 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U52 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U53 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U54 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U55 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U56 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U57 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U58 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U59 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U60 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U61 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U62 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U63 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U64 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U65 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U66 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U67 : MUX2_X1 port map( A => A(21), B => B(21), S => n6, Z => Y(21));
   U68 : MUX2_X1 port map( A => A(20), B => B(20), S => n6, Z => Y(20));
   U69 : MUX2_X1 port map( A => A(19), B => B(19), S => n6, Z => Y(19));
   U70 : MUX2_X1 port map( A => A(18), B => B(18), S => n6, Z => Y(18));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_27 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_27;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_27 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(49), B => B(49), S => n3, Z => Y(49));
   U41 : MUX2_X1 port map( A => A(48), B => B(48), S => n3, Z => Y(48));
   U42 : MUX2_X1 port map( A => A(47), B => B(47), S => n3, Z => Y(47));
   U43 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U44 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U47 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U48 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U49 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U50 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U51 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U52 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U53 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U54 : MUX2_X1 port map( A => A(35), B => B(35), S => n4, Z => Y(35));
   U55 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U56 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U57 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U58 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U59 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U60 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U61 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U62 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U63 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U64 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U65 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U66 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U67 : MUX2_X1 port map( A => A(22), B => B(22), S => n6, Z => Y(22));
   U68 : MUX2_X1 port map( A => A(21), B => B(21), S => n6, Z => Y(21));
   U69 : MUX2_X1 port map( A => A(20), B => B(20), S => n6, Z => Y(20));
   U70 : MUX2_X1 port map( A => A(19), B => B(19), S => n6, Z => Y(19));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_26 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_26;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_26 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U21 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U35 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U36 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U37 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U38 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U39 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U40 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U41 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U44 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U45 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U46 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U47 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U48 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U49 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U50 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U51 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U52 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U53 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U54 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U55 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U56 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U57 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U58 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U59 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U60 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U61 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U62 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U63 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U64 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_25 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_25;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_25 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_24 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_24;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_24 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(50), B => B(50), S => n3, Z => Y(50));
   U41 : MUX2_X1 port map( A => A(49), B => B(49), S => n3, Z => Y(49));
   U42 : MUX2_X1 port map( A => A(48), B => B(48), S => n3, Z => Y(48));
   U43 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U44 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U45 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U46 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U47 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U48 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U49 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U50 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U51 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U52 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U53 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U54 : MUX2_X1 port map( A => A(36), B => B(36), S => n4, Z => Y(36));
   U55 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U56 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U57 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U58 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U59 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U60 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U61 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U62 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U63 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U64 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U65 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U66 : MUX2_X1 port map( A => A(24), B => B(24), S => n5, Z => Y(24));
   U67 : MUX2_X1 port map( A => A(23), B => B(23), S => n6, Z => Y(23));
   U68 : MUX2_X1 port map( A => A(22), B => B(22), S => n6, Z => Y(22));
   U69 : MUX2_X1 port map( A => A(21), B => B(21), S => n6, Z => Y(21));
   U70 : MUX2_X1 port map( A => A(20), B => B(20), S => n6, Z => Y(20));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_23 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_23;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_23 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(51), B => B(51), S => n3, Z => Y(51));
   U41 : MUX2_X1 port map( A => A(50), B => B(50), S => n3, Z => Y(50));
   U42 : MUX2_X1 port map( A => A(49), B => B(49), S => n3, Z => Y(49));
   U43 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U44 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U45 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U48 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U49 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U50 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U51 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U52 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U53 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U54 : MUX2_X1 port map( A => A(37), B => B(37), S => n4, Z => Y(37));
   U55 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U56 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U57 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U58 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U59 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U60 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U61 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U62 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U63 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U64 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U65 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U66 : MUX2_X1 port map( A => A(25), B => B(25), S => n5, Z => Y(25));
   U67 : MUX2_X1 port map( A => A(24), B => B(24), S => n6, Z => Y(24));
   U68 : MUX2_X1 port map( A => A(23), B => B(23), S => n6, Z => Y(23));
   U69 : MUX2_X1 port map( A => A(22), B => B(22), S => n6, Z => Y(22));
   U70 : MUX2_X1 port map( A => A(21), B => B(21), S => n6, Z => Y(21));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_22 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_22;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_22 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U23 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U35 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U36 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U37 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U38 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U39 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U40 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U41 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U42 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U45 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U46 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U47 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U48 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U49 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U50 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U51 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U52 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U53 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U54 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U55 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U56 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U57 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U58 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U59 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U60 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U61 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U62 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U63 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U64 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_21 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_21;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_21 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_20 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_20;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(52), B => B(52), S => n3, Z => Y(52));
   U41 : MUX2_X1 port map( A => A(51), B => B(51), S => n3, Z => Y(51));
   U42 : MUX2_X1 port map( A => A(50), B => B(50), S => n3, Z => Y(50));
   U43 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U44 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U45 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U46 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U47 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U48 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U49 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U50 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U51 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U52 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U53 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U54 : MUX2_X1 port map( A => A(38), B => B(38), S => n4, Z => Y(38));
   U55 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U56 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U57 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U58 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U59 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U60 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U61 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U62 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U63 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U64 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U65 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U66 : MUX2_X1 port map( A => A(26), B => B(26), S => n5, Z => Y(26));
   U67 : MUX2_X1 port map( A => A(25), B => B(25), S => n6, Z => Y(25));
   U68 : MUX2_X1 port map( A => A(24), B => B(24), S => n6, Z => Y(24));
   U69 : MUX2_X1 port map( A => A(23), B => B(23), S => n6, Z => Y(23));
   U70 : MUX2_X1 port map( A => A(22), B => B(22), S => n6, Z => Y(22));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_19 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_19;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(53), B => B(53), S => n3, Z => Y(53));
   U41 : MUX2_X1 port map( A => A(52), B => B(52), S => n3, Z => Y(52));
   U42 : MUX2_X1 port map( A => A(51), B => B(51), S => n3, Z => Y(51));
   U43 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U44 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U45 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U46 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U49 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U50 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U51 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U52 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U53 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U54 : MUX2_X1 port map( A => A(39), B => B(39), S => n4, Z => Y(39));
   U55 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U56 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U57 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U58 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U59 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U60 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U61 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U62 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U63 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U64 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U65 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U66 : MUX2_X1 port map( A => A(27), B => B(27), S => n5, Z => Y(27));
   U67 : MUX2_X1 port map( A => A(26), B => B(26), S => n6, Z => Y(26));
   U68 : MUX2_X1 port map( A => A(25), B => B(25), S => n6, Z => Y(25));
   U69 : MUX2_X1 port map( A => A(24), B => B(24), S => n6, Z => Y(24));
   U70 : MUX2_X1 port map( A => A(23), B => B(23), S => n6, Z => Y(23));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_18 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_18;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U25 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U35 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U36 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U37 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U38 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U39 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U40 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U41 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U42 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U43 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U46 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U47 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U48 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U49 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U50 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U51 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U52 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U53 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U54 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U55 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U56 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U57 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U58 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U59 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U60 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U61 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U62 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U63 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U64 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_17 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_17;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_16 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_16;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(54), B => B(54), S => n3, Z => Y(54));
   U41 : MUX2_X1 port map( A => A(53), B => B(53), S => n3, Z => Y(53));
   U42 : MUX2_X1 port map( A => A(52), B => B(52), S => n3, Z => Y(52));
   U43 : MUX2_X1 port map( A => A(51), B => B(51), S => n4, Z => Y(51));
   U44 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U45 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U46 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U47 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U48 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U49 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U50 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U51 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U52 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U53 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U54 : MUX2_X1 port map( A => A(40), B => B(40), S => n4, Z => Y(40));
   U55 : MUX2_X1 port map( A => A(39), B => B(39), S => n5, Z => Y(39));
   U56 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U57 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U58 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U59 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U60 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U61 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U62 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U63 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U64 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U65 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U66 : MUX2_X1 port map( A => A(28), B => B(28), S => n5, Z => Y(28));
   U67 : MUX2_X1 port map( A => A(27), B => B(27), S => n6, Z => Y(27));
   U68 : MUX2_X1 port map( A => A(26), B => B(26), S => n6, Z => Y(26));
   U69 : MUX2_X1 port map( A => A(25), B => B(25), S => n6, Z => Y(25));
   U70 : MUX2_X1 port map( A => A(24), B => B(24), S => n6, Z => Y(24));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_15 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_15;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U32 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U41 : MUX2_X1 port map( A => A(54), B => B(54), S => n3, Z => Y(54));
   U42 : MUX2_X1 port map( A => A(53), B => B(53), S => n3, Z => Y(53));
   U43 : MUX2_X1 port map( A => A(52), B => B(52), S => n4, Z => Y(52));
   U44 : MUX2_X1 port map( A => A(51), B => B(51), S => n4, Z => Y(51));
   U45 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U46 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U47 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U50 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U51 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U52 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U53 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U54 : MUX2_X1 port map( A => A(41), B => B(41), S => n4, Z => Y(41));
   U55 : MUX2_X1 port map( A => A(40), B => B(40), S => n5, Z => Y(40));
   U56 : MUX2_X1 port map( A => A(39), B => B(39), S => n5, Z => Y(39));
   U57 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U58 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U59 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U60 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U61 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U62 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U63 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U64 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U65 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U66 : MUX2_X1 port map( A => A(29), B => B(29), S => n5, Z => Y(29));
   U67 : MUX2_X1 port map( A => A(28), B => B(28), S => n6, Z => Y(28));
   U68 : MUX2_X1 port map( A => A(27), B => B(27), S => n6, Z => Y(27));
   U69 : MUX2_X1 port map( A => A(26), B => B(26), S => n6, Z => Y(26));
   U70 : MUX2_X1 port map( A => A(25), B => B(25), S => n6, Z => Y(25));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_14 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_14;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U27 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U35 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U36 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U37 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U38 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U39 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U40 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U41 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U42 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U43 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U44 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U47 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U48 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U49 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U50 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U51 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U52 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U53 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U54 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U55 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U56 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U57 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U58 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U59 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U60 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U61 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U62 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U63 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U64 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_13 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_13;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_12 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_12;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U32 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U33 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U41 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U42 : MUX2_X1 port map( A => A(54), B => B(54), S => n3, Z => Y(54));
   U43 : MUX2_X1 port map( A => A(53), B => B(53), S => n4, Z => Y(53));
   U44 : MUX2_X1 port map( A => A(52), B => B(52), S => n4, Z => Y(52));
   U45 : MUX2_X1 port map( A => A(51), B => B(51), S => n4, Z => Y(51));
   U46 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U47 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U48 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U49 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U50 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U51 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U52 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U53 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U54 : MUX2_X1 port map( A => A(42), B => B(42), S => n4, Z => Y(42));
   U55 : MUX2_X1 port map( A => A(41), B => B(41), S => n5, Z => Y(41));
   U56 : MUX2_X1 port map( A => A(40), B => B(40), S => n5, Z => Y(40));
   U57 : MUX2_X1 port map( A => A(39), B => B(39), S => n5, Z => Y(39));
   U58 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U59 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U60 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U61 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U62 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U63 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U64 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U65 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U66 : MUX2_X1 port map( A => A(30), B => B(30), S => n5, Z => Y(30));
   U67 : MUX2_X1 port map( A => A(29), B => B(29), S => n6, Z => Y(29));
   U68 : MUX2_X1 port map( A => A(28), B => B(28), S => n6, Z => Y(28));
   U69 : MUX2_X1 port map( A => A(27), B => B(27), S => n6, Z => Y(27));
   U70 : MUX2_X1 port map( A => A(26), B => B(26), S => n6, Z => Y(26));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_11 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_11;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U32 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U33 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U34 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U41 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U42 : MUX2_X1 port map( A => A(55), B => B(55), S => n3, Z => Y(55));
   U43 : MUX2_X1 port map( A => A(54), B => B(54), S => n4, Z => Y(54));
   U44 : MUX2_X1 port map( A => A(53), B => B(53), S => n4, Z => Y(53));
   U45 : MUX2_X1 port map( A => A(52), B => B(52), S => n4, Z => Y(52));
   U46 : MUX2_X1 port map( A => A(51), B => B(51), S => n4, Z => Y(51));
   U47 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U48 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U51 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U52 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U53 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U54 : MUX2_X1 port map( A => A(43), B => B(43), S => n4, Z => Y(43));
   U55 : MUX2_X1 port map( A => A(42), B => B(42), S => n5, Z => Y(42));
   U56 : MUX2_X1 port map( A => A(41), B => B(41), S => n5, Z => Y(41));
   U57 : MUX2_X1 port map( A => A(40), B => B(40), S => n5, Z => Y(40));
   U58 : MUX2_X1 port map( A => A(39), B => B(39), S => n5, Z => Y(39));
   U59 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U60 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U61 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U62 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U63 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U64 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U65 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U66 : MUX2_X1 port map( A => A(31), B => B(31), S => n5, Z => Y(31));
   U67 : MUX2_X1 port map( A => A(30), B => B(30), S => n6, Z => Y(30));
   U68 : MUX2_X1 port map( A => A(29), B => B(29), S => n6, Z => Y(29));
   U69 : MUX2_X1 port map( A => A(28), B => B(28), S => n6, Z => Y(28));
   U70 : MUX2_X1 port map( A => A(27), B => B(27), S => n6, Z => Y(27));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_10 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_10;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U29 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U35 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U36 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U37 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U38 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U39 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U40 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U41 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U42 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U43 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U44 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U45 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U48 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U49 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U50 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U51 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U52 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U53 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U54 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U55 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U56 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U57 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U58 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U59 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U60 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U61 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U62 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U63 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U64 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_9 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_9;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_8 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_8;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U32 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U33 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U34 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U35 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U41 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U42 : MUX2_X1 port map( A => A(56), B => B(56), S => n3, Z => Y(56));
   U43 : MUX2_X1 port map( A => A(55), B => B(55), S => n4, Z => Y(55));
   U44 : MUX2_X1 port map( A => A(54), B => B(54), S => n4, Z => Y(54));
   U45 : MUX2_X1 port map( A => A(53), B => B(53), S => n4, Z => Y(53));
   U46 : MUX2_X1 port map( A => A(52), B => B(52), S => n4, Z => Y(52));
   U47 : MUX2_X1 port map( A => A(51), B => B(51), S => n4, Z => Y(51));
   U48 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U49 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U50 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U51 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U52 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U53 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U54 : MUX2_X1 port map( A => A(44), B => B(44), S => n4, Z => Y(44));
   U55 : MUX2_X1 port map( A => A(43), B => B(43), S => n5, Z => Y(43));
   U56 : MUX2_X1 port map( A => A(42), B => B(42), S => n5, Z => Y(42));
   U57 : MUX2_X1 port map( A => A(41), B => B(41), S => n5, Z => Y(41));
   U58 : MUX2_X1 port map( A => A(40), B => B(40), S => n5, Z => Y(40));
   U59 : MUX2_X1 port map( A => A(39), B => B(39), S => n5, Z => Y(39));
   U60 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U61 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U62 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U63 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U64 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U65 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U66 : MUX2_X1 port map( A => A(32), B => B(32), S => n5, Z => Y(32));
   U67 : MUX2_X1 port map( A => A(31), B => B(31), S => n6, Z => Y(31));
   U68 : MUX2_X1 port map( A => A(30), B => B(30), S => n6, Z => Y(30));
   U69 : MUX2_X1 port map( A => A(29), B => B(29), S => n6, Z => Y(29));
   U70 : MUX2_X1 port map( A => A(28), B => B(28), S => n6, Z => Y(28));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_7 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_7;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U32 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U33 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U34 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U35 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Y(28));
   U36 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U41 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U42 : MUX2_X1 port map( A => A(57), B => B(57), S => n3, Z => Y(57));
   U43 : MUX2_X1 port map( A => A(56), B => B(56), S => n4, Z => Y(56));
   U44 : MUX2_X1 port map( A => A(55), B => B(55), S => n4, Z => Y(55));
   U45 : MUX2_X1 port map( A => A(54), B => B(54), S => n4, Z => Y(54));
   U46 : MUX2_X1 port map( A => A(53), B => B(53), S => n4, Z => Y(53));
   U47 : MUX2_X1 port map( A => A(52), B => B(52), S => n4, Z => Y(52));
   U48 : MUX2_X1 port map( A => A(51), B => B(51), S => n4, Z => Y(51));
   U49 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U52 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U53 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U54 : MUX2_X1 port map( A => A(45), B => B(45), S => n4, Z => Y(45));
   U55 : MUX2_X1 port map( A => A(44), B => B(44), S => n5, Z => Y(44));
   U56 : MUX2_X1 port map( A => A(43), B => B(43), S => n5, Z => Y(43));
   U57 : MUX2_X1 port map( A => A(42), B => B(42), S => n5, Z => Y(42));
   U58 : MUX2_X1 port map( A => A(41), B => B(41), S => n5, Z => Y(41));
   U59 : MUX2_X1 port map( A => A(40), B => B(40), S => n5, Z => Y(40));
   U60 : MUX2_X1 port map( A => A(39), B => B(39), S => n5, Z => Y(39));
   U61 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U62 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U63 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U64 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U65 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U66 : MUX2_X1 port map( A => A(33), B => B(33), S => n5, Z => Y(33));
   U67 : MUX2_X1 port map( A => A(32), B => B(32), S => n6, Z => Y(32));
   U68 : MUX2_X1 port map( A => A(31), B => B(31), S => n6, Z => Y(31));
   U69 : MUX2_X1 port map( A => A(30), B => B(30), S => n6, Z => Y(30));
   U70 : MUX2_X1 port map( A => A(29), B => B(29), S => n6, Z => Y(29));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_6 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_6;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U31 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U35 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U36 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U37 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U38 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U39 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U40 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U41 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U42 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U43 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U44 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U45 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U46 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U49 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U50 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U51 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U52 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U53 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U54 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U55 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U56 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U57 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U58 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U59 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U60 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U61 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U62 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U63 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U64 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_5 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_5;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_4 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_4;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U32 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U33 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U34 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U35 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Y(28));
   U36 : MUX2_X1 port map( A => A(29), B => B(29), S => n3, Z => Y(29));
   U37 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U41 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U42 : MUX2_X1 port map( A => A(58), B => B(58), S => n3, Z => Y(58));
   U43 : MUX2_X1 port map( A => A(57), B => B(57), S => n4, Z => Y(57));
   U44 : MUX2_X1 port map( A => A(56), B => B(56), S => n4, Z => Y(56));
   U45 : MUX2_X1 port map( A => A(55), B => B(55), S => n4, Z => Y(55));
   U46 : MUX2_X1 port map( A => A(54), B => B(54), S => n4, Z => Y(54));
   U47 : MUX2_X1 port map( A => A(53), B => B(53), S => n4, Z => Y(53));
   U48 : MUX2_X1 port map( A => A(52), B => B(52), S => n4, Z => Y(52));
   U49 : MUX2_X1 port map( A => A(51), B => B(51), S => n4, Z => Y(51));
   U50 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U51 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U52 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U53 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U54 : MUX2_X1 port map( A => A(46), B => B(46), S => n4, Z => Y(46));
   U55 : MUX2_X1 port map( A => A(45), B => B(45), S => n5, Z => Y(45));
   U56 : MUX2_X1 port map( A => A(44), B => B(44), S => n5, Z => Y(44));
   U57 : MUX2_X1 port map( A => A(43), B => B(43), S => n5, Z => Y(43));
   U58 : MUX2_X1 port map( A => A(42), B => B(42), S => n5, Z => Y(42));
   U59 : MUX2_X1 port map( A => A(41), B => B(41), S => n5, Z => Y(41));
   U60 : MUX2_X1 port map( A => A(40), B => B(40), S => n5, Z => Y(40));
   U61 : MUX2_X1 port map( A => A(39), B => B(39), S => n5, Z => Y(39));
   U62 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U63 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U64 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U65 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U66 : MUX2_X1 port map( A => A(34), B => B(34), S => n5, Z => Y(34));
   U67 : MUX2_X1 port map( A => A(33), B => B(33), S => n6, Z => Y(33));
   U68 : MUX2_X1 port map( A => A(32), B => B(32), S => n6, Z => Y(32));
   U69 : MUX2_X1 port map( A => A(31), B => B(31), S => n6, Z => Y(31));
   U70 : MUX2_X1 port map( A => A(30), B => B(30), S => n6, Z => Y(30));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_3 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_3;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(0), B => B(0), S => n1, Z => Y(0));
   U8 : MUX2_X1 port map( A => A(1), B => B(1), S => n1, Z => Y(1));
   U9 : MUX2_X1 port map( A => A(2), B => B(2), S => n1, Z => Y(2));
   U10 : MUX2_X1 port map( A => A(3), B => B(3), S => n1, Z => Y(3));
   U11 : MUX2_X1 port map( A => A(4), B => B(4), S => n1, Z => Y(4));
   U12 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U13 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U16 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U17 : MUX2_X1 port map( A => A(10), B => B(10), S => n1, Z => Y(10));
   U18 : MUX2_X1 port map( A => A(11), B => B(11), S => n1, Z => Y(11));
   U19 : MUX2_X1 port map( A => A(12), B => B(12), S => n2, Z => Y(12));
   U20 : MUX2_X1 port map( A => A(13), B => B(13), S => n2, Z => Y(13));
   U21 : MUX2_X1 port map( A => A(14), B => B(14), S => n2, Z => Y(14));
   U22 : MUX2_X1 port map( A => A(15), B => B(15), S => n2, Z => Y(15));
   U23 : MUX2_X1 port map( A => A(16), B => B(16), S => n2, Z => Y(16));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => n2, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => n2, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(19), B => B(19), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => A(20), B => B(20), S => n2, Z => Y(20));
   U28 : MUX2_X1 port map( A => A(21), B => B(21), S => n2, Z => Y(21));
   U29 : MUX2_X1 port map( A => A(22), B => B(22), S => n2, Z => Y(22));
   U30 : MUX2_X1 port map( A => A(23), B => B(23), S => n2, Z => Y(23));
   U31 : MUX2_X1 port map( A => A(24), B => B(24), S => n3, Z => Y(24));
   U32 : MUX2_X1 port map( A => A(25), B => B(25), S => n3, Z => Y(25));
   U33 : MUX2_X1 port map( A => A(26), B => B(26), S => n3, Z => Y(26));
   U34 : MUX2_X1 port map( A => A(27), B => B(27), S => n3, Z => Y(27));
   U35 : MUX2_X1 port map( A => A(28), B => B(28), S => n3, Z => Y(28));
   U36 : MUX2_X1 port map( A => A(29), B => B(29), S => n3, Z => Y(29));
   U37 : MUX2_X1 port map( A => A(30), B => B(30), S => n3, Z => Y(30));
   U38 : MUX2_X1 port map( A => A(62), B => B(62), S => n3, Z => Y(62));
   U39 : MUX2_X1 port map( A => A(63), B => B(63), S => n3, Z => Y(63));
   U40 : MUX2_X1 port map( A => A(61), B => B(61), S => n3, Z => Y(61));
   U41 : MUX2_X1 port map( A => A(60), B => B(60), S => n3, Z => Y(60));
   U42 : MUX2_X1 port map( A => A(59), B => B(59), S => n3, Z => Y(59));
   U43 : MUX2_X1 port map( A => A(58), B => B(58), S => n4, Z => Y(58));
   U44 : MUX2_X1 port map( A => A(57), B => B(57), S => n4, Z => Y(57));
   U45 : MUX2_X1 port map( A => A(56), B => B(56), S => n4, Z => Y(56));
   U46 : MUX2_X1 port map( A => A(55), B => B(55), S => n4, Z => Y(55));
   U47 : MUX2_X1 port map( A => A(54), B => B(54), S => n4, Z => Y(54));
   U48 : MUX2_X1 port map( A => A(53), B => B(53), S => n4, Z => Y(53));
   U49 : MUX2_X1 port map( A => A(52), B => B(52), S => n4, Z => Y(52));
   U50 : MUX2_X1 port map( A => A(51), B => B(51), S => n4, Z => Y(51));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => n4, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(49), B => B(49), S => n4, Z => Y(49));
   U53 : MUX2_X1 port map( A => A(48), B => B(48), S => n4, Z => Y(48));
   U54 : MUX2_X1 port map( A => A(47), B => B(47), S => n4, Z => Y(47));
   U55 : MUX2_X1 port map( A => A(46), B => B(46), S => n5, Z => Y(46));
   U56 : MUX2_X1 port map( A => A(45), B => B(45), S => n5, Z => Y(45));
   U57 : MUX2_X1 port map( A => A(44), B => B(44), S => n5, Z => Y(44));
   U58 : MUX2_X1 port map( A => A(43), B => B(43), S => n5, Z => Y(43));
   U59 : MUX2_X1 port map( A => A(42), B => B(42), S => n5, Z => Y(42));
   U60 : MUX2_X1 port map( A => A(41), B => B(41), S => n5, Z => Y(41));
   U61 : MUX2_X1 port map( A => A(40), B => B(40), S => n5, Z => Y(40));
   U62 : MUX2_X1 port map( A => A(39), B => B(39), S => n5, Z => Y(39));
   U63 : MUX2_X1 port map( A => A(38), B => B(38), S => n5, Z => Y(38));
   U64 : MUX2_X1 port map( A => A(37), B => B(37), S => n5, Z => Y(37));
   U65 : MUX2_X1 port map( A => A(36), B => B(36), S => n5, Z => Y(36));
   U66 : MUX2_X1 port map( A => A(35), B => B(35), S => n5, Z => Y(35));
   U67 : MUX2_X1 port map( A => A(34), B => B(34), S => n6, Z => Y(34));
   U68 : MUX2_X1 port map( A => A(33), B => B(33), S => n6, Z => Y(33));
   U69 : MUX2_X1 port map( A => A(32), B => B(32), S => n6, Z => Y(32));
   U70 : MUX2_X1 port map( A => A(31), B => B(31), S => n6, Z => Y(31));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_2 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_2;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U33 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));
   U34 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U35 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U36 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U37 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U38 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U39 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U40 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U41 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U42 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U43 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U44 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U45 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U46 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U47 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U50 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U51 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U52 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U53 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U54 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U55 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U56 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U57 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U58 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U59 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U60 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U61 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U62 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U63 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U64 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_1;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U5 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U6 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U7 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U8 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U9 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U10 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U11 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U12 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U13 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U14 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U15 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U16 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U17 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U18 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U19 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U22 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U23 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U24 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U25 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U26 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U27 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U28 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U29 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U30 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U31 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U32 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U33 : MUX2_X1 port map( A => A(32), B => B(32), S => SEL, Z => Y(32));
   U34 : MUX2_X1 port map( A => A(33), B => B(33), S => SEL, Z => Y(33));
   U35 : MUX2_X1 port map( A => A(34), B => B(34), S => SEL, Z => Y(34));
   U36 : MUX2_X1 port map( A => A(35), B => B(35), S => SEL, Z => Y(35));
   U37 : MUX2_X1 port map( A => A(36), B => B(36), S => SEL, Z => Y(36));
   U38 : MUX2_X1 port map( A => A(37), B => B(37), S => SEL, Z => Y(37));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => SEL, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(39), B => B(39), S => SEL, Z => Y(39));
   U41 : MUX2_X1 port map( A => A(40), B => B(40), S => SEL, Z => Y(40));
   U42 : MUX2_X1 port map( A => A(41), B => B(41), S => SEL, Z => Y(41));
   U43 : MUX2_X1 port map( A => A(42), B => B(42), S => SEL, Z => Y(42));
   U44 : MUX2_X1 port map( A => A(43), B => B(43), S => SEL, Z => Y(43));
   U45 : MUX2_X1 port map( A => A(44), B => B(44), S => SEL, Z => Y(44));
   U46 : MUX2_X1 port map( A => A(45), B => B(45), S => SEL, Z => Y(45));
   U47 : MUX2_X1 port map( A => A(46), B => B(46), S => SEL, Z => Y(46));
   U48 : MUX2_X1 port map( A => A(47), B => B(47), S => SEL, Z => Y(47));
   U49 : MUX2_X1 port map( A => A(48), B => B(48), S => SEL, Z => Y(48));
   U50 : MUX2_X1 port map( A => A(49), B => B(49), S => SEL, Z => Y(49));
   U51 : MUX2_X1 port map( A => A(50), B => B(50), S => SEL, Z => Y(50));
   U52 : MUX2_X1 port map( A => A(51), B => B(51), S => SEL, Z => Y(51));
   U53 : MUX2_X1 port map( A => A(52), B => B(52), S => SEL, Z => Y(52));
   U54 : MUX2_X1 port map( A => A(53), B => B(53), S => SEL, Z => Y(53));
   U55 : MUX2_X1 port map( A => A(54), B => B(54), S => SEL, Z => Y(54));
   U56 : MUX2_X1 port map( A => A(55), B => B(55), S => SEL, Z => Y(55));
   U57 : MUX2_X1 port map( A => A(56), B => B(56), S => SEL, Z => Y(56));
   U58 : MUX2_X1 port map( A => A(57), B => B(57), S => SEL, Z => Y(57));
   U59 : MUX2_X1 port map( A => A(58), B => B(58), S => SEL, Z => Y(58));
   U60 : MUX2_X1 port map( A => A(59), B => B(59), S => SEL, Z => Y(59));
   U61 : MUX2_X1 port map( A => A(60), B => B(60), S => SEL, Z => Y(60));
   U62 : MUX2_X1 port map( A => A(61), B => B(61), S => SEL, Z => Y(61));
   U63 : MUX2_X1 port map( A => A(62), B => B(62), S => SEL, Z => Y(62));
   U64 : MUX2_X1 port map( A => A(63), B => B(63), S => SEL, Z => Y(63));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_14 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_14;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_14 is

   component RCA_GENERIC_NBIT64_14_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1077 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_14_DW01_add_0 port map( A(64) => n2
                           , A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1077);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_13 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_13;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_13 is

   component RCA_GENERIC_NBIT64_13_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1078 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_13_DW01_add_0 port map( A(64) => n2
                           , A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1078);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_12 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_12;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_12 is

   component RCA_GENERIC_NBIT64_12_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1079 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_12_DW01_add_0 port map( A(64) => n2
                           , A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1079);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_11 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_11;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_11 is

   component RCA_GENERIC_NBIT64_11_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1080 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_11_DW01_add_0 port map( A(64) => n2
                           , A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1080);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_10 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_10;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_10 is

   component RCA_GENERIC_NBIT64_10_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1081 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_10_DW01_add_0 port map( A(64) => n2
                           , A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1081);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_9 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_9;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_9 is

   component RCA_GENERIC_NBIT64_9_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1082 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_9_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1082);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_8 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_8;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_8 is

   component RCA_GENERIC_NBIT64_8_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1083 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_8_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1083);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_7 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_7;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_7 is

   component RCA_GENERIC_NBIT64_7_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1084 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_7_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1084);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_6 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_6;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_6 is

   component RCA_GENERIC_NBIT64_6_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1085 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_6_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1085);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_5 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_5;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_5 is

   component RCA_GENERIC_NBIT64_5_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1086 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_5_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1086);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_4 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_4;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_4 is

   component RCA_GENERIC_NBIT64_4_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1087 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_4_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1087);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_3 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_3;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_3 is

   component RCA_GENERIC_NBIT64_3_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1088 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_3_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1088);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_2 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_2;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_2 is

   component RCA_GENERIC_NBIT64_2_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1089 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_2_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1089);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_1;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_1 is

   component RCA_GENERIC_NBIT64_1_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1090 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_1_DW01_add_0 port map( A(64) => n2,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n2, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1090);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_15 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_15;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_15 is

   component MUX21_GENERIC_NBIT64_57
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_58
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_59
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_60
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_60 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_59 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_58 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_57 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_14 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_14;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_14 is

   component MUX21_GENERIC_NBIT64_53
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_54
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_55
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_56
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_56 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_55 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_54 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_53 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_13 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_13;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_13 is

   component MUX21_GENERIC_NBIT64_49
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_50
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_51
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_52
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_52 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_51 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_50 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_49 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_12 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_12;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_12 is

   component MUX21_GENERIC_NBIT64_45
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_46
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_47
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_48
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_48 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_47 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_46 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_45 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_11 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_11;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_11 is

   component MUX21_GENERIC_NBIT64_41
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_42
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_43
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_44
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_44 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_43 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_42 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_41 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_10 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_10;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_10 is

   component MUX21_GENERIC_NBIT64_37
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_38
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_39
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_40
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_40 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_39 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_38 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_37 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_9 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_9;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_9 is

   component MUX21_GENERIC_NBIT64_33
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_34
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_35
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_36
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_36 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_35 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_34 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_33 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_8 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_8;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_8 is

   component MUX21_GENERIC_NBIT64_29
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_30
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_31
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_32
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_32 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_31 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_30 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_29 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_7 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_7;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_7 is

   component MUX21_GENERIC_NBIT64_25
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_26
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_27
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_28
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_28 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_27 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_26 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_25 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_6 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_6;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_6 is

   component MUX21_GENERIC_NBIT64_21
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_22
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_23
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_24
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_24 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_23 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_22 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_21 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_5 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_5;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_5 is

   component MUX21_GENERIC_NBIT64_17
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_18
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_19
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_20
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_20 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_19 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_18 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_17 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_4 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_4;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_4 is

   component MUX21_GENERIC_NBIT64_13
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_14
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_15
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_16
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_16 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_15 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_14 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_13 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_3 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_3;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_3 is

   component MUX21_GENERIC_NBIT64_9
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_10
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_11
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_12
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_12 port map( A(63) => IN2(63), A(62) => IN2(62)
                           , A(61) => IN2(61), A(60) => IN2(60), A(59) => 
                           IN2(59), A(58) => IN2(58), A(57) => IN2(57), A(56) 
                           => IN2(56), A(55) => IN2(55), A(54) => IN2(54), 
                           A(53) => IN2(53), A(52) => IN2(52), A(51) => IN2(51)
                           , A(50) => IN2(50), A(49) => IN2(49), A(48) => 
                           IN2(48), A(47) => IN2(47), A(46) => IN2(46), A(45) 
                           => IN2(45), A(44) => IN2(44), A(43) => IN2(43), 
                           A(42) => IN2(42), A(41) => IN2(41), A(40) => IN2(40)
                           , A(39) => IN2(39), A(38) => IN2(38), A(37) => 
                           IN2(37), A(36) => IN2(36), A(35) => IN2(35), A(34) 
                           => IN2(34), A(33) => IN2(33), A(32) => IN2(32), 
                           A(31) => IN2(31), A(30) => IN2(30), A(29) => IN2(29)
                           , A(28) => IN2(28), A(27) => IN2(27), A(26) => 
                           IN2(26), A(25) => IN2(25), A(24) => IN2(24), A(23) 
                           => IN2(23), A(22) => IN2(22), A(21) => IN2(21), 
                           A(20) => IN2(20), A(19) => IN2(19), A(18) => IN2(18)
                           , A(17) => IN2(17), A(16) => IN2(16), A(15) => 
                           IN2(15), A(14) => IN2(14), A(13) => IN2(13), A(12) 
                           => IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9)
                           => IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_11 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_10 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_9 port map( A(63) => IN0(63), A(62) => IN0(62), 
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_2 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_2;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_2 is

   component MUX21_GENERIC_NBIT64_5
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_6
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_7
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_8
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_8 port map( A(63) => IN2(63), A(62) => IN2(62),
                           A(61) => IN2(61), A(60) => IN2(60), A(59) => IN2(59)
                           , A(58) => IN2(58), A(57) => IN2(57), A(56) => 
                           IN2(56), A(55) => IN2(55), A(54) => IN2(54), A(53) 
                           => IN2(53), A(52) => IN2(52), A(51) => IN2(51), 
                           A(50) => IN2(50), A(49) => IN2(49), A(48) => IN2(48)
                           , A(47) => IN2(47), A(46) => IN2(46), A(45) => 
                           IN2(45), A(44) => IN2(44), A(43) => IN2(43), A(42) 
                           => IN2(42), A(41) => IN2(41), A(40) => IN2(40), 
                           A(39) => IN2(39), A(38) => IN2(38), A(37) => IN2(37)
                           , A(36) => IN2(36), A(35) => IN2(35), A(34) => 
                           IN2(34), A(33) => IN2(33), A(32) => IN2(32), A(31) 
                           => IN2(31), A(30) => IN2(30), A(29) => IN2(29), 
                           A(28) => IN2(28), A(27) => IN2(27), A(26) => IN2(26)
                           , A(25) => IN2(25), A(24) => IN2(24), A(23) => 
                           IN2(23), A(22) => IN2(22), A(21) => IN2(21), A(20) 
                           => IN2(20), A(19) => IN2(19), A(18) => IN2(18), 
                           A(17) => IN2(17), A(16) => IN2(16), A(15) => IN2(15)
                           , A(14) => IN2(14), A(13) => IN2(13), A(12) => 
                           IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9) =>
                           IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_7 port map( A(63) => IN4(63), A(62) => IN4(62),
                           A(61) => IN4(61), A(60) => IN4(60), A(59) => IN4(59)
                           , A(58) => IN4(58), A(57) => IN4(57), A(56) => 
                           IN4(56), A(55) => IN4(55), A(54) => IN4(54), A(53) 
                           => IN4(53), A(52) => IN4(52), A(51) => IN4(51), 
                           A(50) => IN4(50), A(49) => IN4(49), A(48) => IN4(48)
                           , A(47) => IN4(47), A(46) => IN4(46), A(45) => 
                           IN4(45), A(44) => IN4(44), A(43) => IN4(43), A(42) 
                           => IN4(42), A(41) => IN4(41), A(40) => IN4(40), 
                           A(39) => IN4(39), A(38) => IN4(38), A(37) => IN4(37)
                           , A(36) => IN4(36), A(35) => IN4(35), A(34) => 
                           IN4(34), A(33) => IN4(33), A(32) => IN4(32), A(31) 
                           => IN4(31), A(30) => IN4(30), A(29) => IN4(29), 
                           A(28) => IN4(28), A(27) => IN4(27), A(26) => IN4(26)
                           , A(25) => IN4(25), A(24) => IN4(24), A(23) => 
                           IN4(23), A(22) => IN4(22), A(21) => IN4(21), A(20) 
                           => IN4(20), A(19) => IN4(19), A(18) => IN4(18), 
                           A(17) => IN4(17), A(16) => IN4(16), A(15) => IN4(15)
                           , A(14) => IN4(14), A(13) => IN4(13), A(12) => 
                           IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9) =>
                           IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_6 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_5 port map( A(63) => IN0(63), A(62) => IN0(62), 
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_1 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_1;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_1 is

   component MUX21_GENERIC_NBIT64_1
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_2
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_3
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_4
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_4 port map( A(63) => IN2(63), A(62) => IN2(62),
                           A(61) => IN2(61), A(60) => IN2(60), A(59) => IN2(59)
                           , A(58) => IN2(58), A(57) => IN2(57), A(56) => 
                           IN2(56), A(55) => IN2(55), A(54) => IN2(54), A(53) 
                           => IN2(53), A(52) => IN2(52), A(51) => IN2(51), 
                           A(50) => IN2(50), A(49) => IN2(49), A(48) => IN2(48)
                           , A(47) => IN2(47), A(46) => IN2(46), A(45) => 
                           IN2(45), A(44) => IN2(44), A(43) => IN2(43), A(42) 
                           => IN2(42), A(41) => IN2(41), A(40) => IN2(40), 
                           A(39) => IN2(39), A(38) => IN2(38), A(37) => IN2(37)
                           , A(36) => IN2(36), A(35) => IN2(35), A(34) => 
                           IN2(34), A(33) => IN2(33), A(32) => IN2(32), A(31) 
                           => IN2(31), A(30) => IN2(30), A(29) => IN2(29), 
                           A(28) => IN2(28), A(27) => IN2(27), A(26) => IN2(26)
                           , A(25) => IN2(25), A(24) => IN2(24), A(23) => 
                           IN2(23), A(22) => IN2(22), A(21) => IN2(21), A(20) 
                           => IN2(20), A(19) => IN2(19), A(18) => IN2(18), 
                           A(17) => IN2(17), A(16) => IN2(16), A(15) => IN2(15)
                           , A(14) => IN2(14), A(13) => IN2(13), A(12) => 
                           IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9) =>
                           IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_3 port map( A(63) => IN4(63), A(62) => IN4(62),
                           A(61) => IN4(61), A(60) => IN4(60), A(59) => IN4(59)
                           , A(58) => IN4(58), A(57) => IN4(57), A(56) => 
                           IN4(56), A(55) => IN4(55), A(54) => IN4(54), A(53) 
                           => IN4(53), A(52) => IN4(52), A(51) => IN4(51), 
                           A(50) => IN4(50), A(49) => IN4(49), A(48) => IN4(48)
                           , A(47) => IN4(47), A(46) => IN4(46), A(45) => 
                           IN4(45), A(44) => IN4(44), A(43) => IN4(43), A(42) 
                           => IN4(42), A(41) => IN4(41), A(40) => IN4(40), 
                           A(39) => IN4(39), A(38) => IN4(38), A(37) => IN4(37)
                           , A(36) => IN4(36), A(35) => IN4(35), A(34) => 
                           IN4(34), A(33) => IN4(33), A(32) => IN4(32), A(31) 
                           => IN4(31), A(30) => IN4(30), A(29) => IN4(29), 
                           A(28) => IN4(28), A(27) => IN4(27), A(26) => IN4(26)
                           , A(25) => IN4(25), A(24) => IN4(24), A(23) => 
                           IN4(23), A(22) => IN4(22), A(21) => IN4(21), A(20) 
                           => IN4(20), A(19) => IN4(19), A(18) => IN4(18), 
                           A(17) => IN4(17), A(16) => IN4(16), A(15) => IN4(15)
                           , A(14) => IN4(14), A(13) => IN4(13), A(12) => 
                           IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9) =>
                           IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_2 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_1 port map( A(63) => IN0(63), A(62) => IN0(62), 
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_19 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_19;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_18 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_18;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_17 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_17;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_16 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_16;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_15 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_15;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_14 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_14;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_13 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_13;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_12 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_12;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_11 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_11;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_10 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_10;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_9 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_9;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_8 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_8;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_7 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_7;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_6 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_6;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_5 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_5;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX21_GENERIC_NBIT64_0 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_NBIT64_0;

architecture SYN_BEH of MUX21_GENERIC_NBIT64_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X1 port map( A => SEL, Z => n3);
   U4 : CLKBUF_X1 port map( A => SEL, Z => n4);
   U5 : CLKBUF_X1 port map( A => SEL, Z => n5);
   U6 : CLKBUF_X1 port map( A => SEL, Z => n6);
   U7 : MUX2_X1 port map( A => A(9), B => B(9), S => n1, Z => Y(9));
   U8 : MUX2_X1 port map( A => A(8), B => B(8), S => n1, Z => Y(8));
   U9 : MUX2_X1 port map( A => A(7), B => B(7), S => n1, Z => Y(7));
   U10 : MUX2_X1 port map( A => A(6), B => B(6), S => n1, Z => Y(6));
   U11 : MUX2_X1 port map( A => A(63), B => B(63), S => n1, Z => Y(63));
   U12 : MUX2_X1 port map( A => A(62), B => B(62), S => n1, Z => Y(62));
   U13 : MUX2_X1 port map( A => A(61), B => B(61), S => n1, Z => Y(61));
   U14 : MUX2_X1 port map( A => A(60), B => B(60), S => n1, Z => Y(60));
   U15 : MUX2_X1 port map( A => A(5), B => B(5), S => n1, Z => Y(5));
   U16 : MUX2_X1 port map( A => A(59), B => B(59), S => n1, Z => Y(59));
   U17 : MUX2_X1 port map( A => A(58), B => B(58), S => n1, Z => Y(58));
   U18 : MUX2_X1 port map( A => A(57), B => B(57), S => n1, Z => Y(57));
   U19 : MUX2_X1 port map( A => A(56), B => B(56), S => n2, Z => Y(56));
   U20 : MUX2_X1 port map( A => A(55), B => B(55), S => n2, Z => Y(55));
   U21 : MUX2_X1 port map( A => A(54), B => B(54), S => n2, Z => Y(54));
   U22 : MUX2_X1 port map( A => A(53), B => B(53), S => n2, Z => Y(53));
   U23 : MUX2_X1 port map( A => A(52), B => B(52), S => n2, Z => Y(52));
   U24 : MUX2_X1 port map( A => A(51), B => B(51), S => n2, Z => Y(51));
   U25 : MUX2_X1 port map( A => A(50), B => B(50), S => n2, Z => Y(50));
   U26 : MUX2_X1 port map( A => A(4), B => B(4), S => n2, Z => Y(4));
   U27 : MUX2_X1 port map( A => A(49), B => B(49), S => n2, Z => Y(49));
   U28 : MUX2_X1 port map( A => A(48), B => B(48), S => n2, Z => Y(48));
   U29 : MUX2_X1 port map( A => A(47), B => B(47), S => n2, Z => Y(47));
   U30 : MUX2_X1 port map( A => A(46), B => B(46), S => n2, Z => Y(46));
   U31 : MUX2_X1 port map( A => A(45), B => B(45), S => n3, Z => Y(45));
   U32 : MUX2_X1 port map( A => A(44), B => B(44), S => n3, Z => Y(44));
   U33 : MUX2_X1 port map( A => A(43), B => B(43), S => n3, Z => Y(43));
   U34 : MUX2_X1 port map( A => A(42), B => B(42), S => n3, Z => Y(42));
   U35 : MUX2_X1 port map( A => A(41), B => B(41), S => n3, Z => Y(41));
   U36 : MUX2_X1 port map( A => A(40), B => B(40), S => n3, Z => Y(40));
   U37 : MUX2_X1 port map( A => A(3), B => B(3), S => n3, Z => Y(3));
   U38 : MUX2_X1 port map( A => A(39), B => B(39), S => n3, Z => Y(39));
   U39 : MUX2_X1 port map( A => A(38), B => B(38), S => n3, Z => Y(38));
   U40 : MUX2_X1 port map( A => A(37), B => B(37), S => n3, Z => Y(37));
   U41 : MUX2_X1 port map( A => A(36), B => B(36), S => n3, Z => Y(36));
   U42 : MUX2_X1 port map( A => A(35), B => B(35), S => n3, Z => Y(35));
   U43 : MUX2_X1 port map( A => A(34), B => B(34), S => n4, Z => Y(34));
   U44 : MUX2_X1 port map( A => A(33), B => B(33), S => n4, Z => Y(33));
   U45 : MUX2_X1 port map( A => A(32), B => B(32), S => n4, Z => Y(32));
   U46 : MUX2_X1 port map( A => A(31), B => B(31), S => n4, Z => Y(31));
   U47 : MUX2_X1 port map( A => A(30), B => B(30), S => n4, Z => Y(30));
   U48 : MUX2_X1 port map( A => A(2), B => B(2), S => n4, Z => Y(2));
   U49 : MUX2_X1 port map( A => A(29), B => B(29), S => n4, Z => Y(29));
   U50 : MUX2_X1 port map( A => A(28), B => B(28), S => n4, Z => Y(28));
   U51 : MUX2_X1 port map( A => A(27), B => B(27), S => n4, Z => Y(27));
   U52 : MUX2_X1 port map( A => A(26), B => B(26), S => n4, Z => Y(26));
   U53 : MUX2_X1 port map( A => A(25), B => B(25), S => n4, Z => Y(25));
   U54 : MUX2_X1 port map( A => A(24), B => B(24), S => n4, Z => Y(24));
   U55 : MUX2_X1 port map( A => A(23), B => B(23), S => n5, Z => Y(23));
   U56 : MUX2_X1 port map( A => A(22), B => B(22), S => n5, Z => Y(22));
   U57 : MUX2_X1 port map( A => A(21), B => B(21), S => n5, Z => Y(21));
   U58 : MUX2_X1 port map( A => A(20), B => B(20), S => n5, Z => Y(20));
   U59 : MUX2_X1 port map( A => A(1), B => B(1), S => n5, Z => Y(1));
   U60 : MUX2_X1 port map( A => A(19), B => B(19), S => n5, Z => Y(19));
   U61 : MUX2_X1 port map( A => A(18), B => B(18), S => n5, Z => Y(18));
   U62 : MUX2_X1 port map( A => A(17), B => B(17), S => n5, Z => Y(17));
   U63 : MUX2_X1 port map( A => A(16), B => B(16), S => n5, Z => Y(16));
   U64 : MUX2_X1 port map( A => A(15), B => B(15), S => n5, Z => Y(15));
   U65 : MUX2_X1 port map( A => A(14), B => B(14), S => n5, Z => Y(14));
   U66 : MUX2_X1 port map( A => A(13), B => B(13), S => n5, Z => Y(13));
   U67 : MUX2_X1 port map( A => A(12), B => B(12), S => n6, Z => Y(12));
   U68 : MUX2_X1 port map( A => A(11), B => B(11), S => n6, Z => Y(11));
   U69 : MUX2_X1 port map( A => A(10), B => B(10), S => n6, Z => Y(10));
   U70 : MUX2_X1 port map( A => A(0), B => B(0), S => n6, Z => Y(0));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_GENERIC_NBIT64_0 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT64_0;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT64_0 is

   component RCA_GENERIC_NBIT64_0_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1091 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_23_2 : RCA_GENERIC_NBIT64_0_DW01_add_0 port map( A(64) => n1,
                           A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(64) => n1, B(63)
                           => B(63), B(62) => B(62), B(61) => B(61), B(60) => 
                           B(60), B(59) => B(59), B(58) => B(58), B(57) => 
                           B(57), B(56) => B(56), B(55) => B(55), B(54) => 
                           B(54), B(53) => B(53), B(52) => B(52), B(51) => 
                           B(51), B(50) => B(50), B(49) => B(49), B(48) => 
                           B(48), B(47) => B(47), B(46) => B(46), B(45) => 
                           B(45), B(44) => B(44), B(43) => B(43), B(42) => 
                           B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, 
                           SUM(63) => S(63), SUM(62) => S(62), SUM(61) => S(61)
                           , SUM(60) => S(60), SUM(59) => S(59), SUM(58) => 
                           S(58), SUM(57) => S(57), SUM(56) => S(56), SUM(55) 
                           => S(55), SUM(54) => S(54), SUM(53) => S(53), 
                           SUM(52) => S(52), SUM(51) => S(51), SUM(50) => S(50)
                           , SUM(49) => S(49), SUM(48) => S(48), SUM(47) => 
                           S(47), SUM(46) => S(46), SUM(45) => S(45), SUM(44) 
                           => S(44), SUM(43) => S(43), SUM(42) => S(42), 
                           SUM(41) => S(41), SUM(40) => S(40), SUM(39) => S(39)
                           , SUM(38) => S(38), SUM(37) => S(37), SUM(36) => 
                           S(36), SUM(35) => S(35), SUM(34) => S(34), SUM(33) 
                           => S(33), SUM(32) => S(32), SUM(31) => S(31), 
                           SUM(30) => S(30), SUM(29) => S(29), SUM(28) => S(28)
                           , SUM(27) => S(27), SUM(26) => S(26), SUM(25) => 
                           S(25), SUM(24) => S(24), SUM(23) => S(23), SUM(22) 
                           => S(22), SUM(21) => S(21), SUM(20) => S(20), 
                           SUM(19) => S(19), SUM(18) => S(18), SUM(17) => S(17)
                           , SUM(16) => S(16), SUM(15) => S(15), SUM(14) => 
                           S(14), SUM(13) => S(13), SUM(12) => S(12), SUM(11) 
                           => S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) 
                           => S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => 
                           S(5), SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2)
                           , SUM(1) => S(1), SUM(0) => S(0), CO => n_1091);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity MUX51_GENERIC_NBIT64_0 is

   port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : in 
         std_logic_vector (2 downto 0);  O : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_NBIT64_0;

architecture SYN_mux51_struct of MUX51_GENERIC_NBIT64_0 is

   component MUX21_GENERIC_NBIT64_61
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_62
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_63
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT64_0
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal temp00_63_port, temp00_62_port, temp00_61_port, temp00_60_port, 
      temp00_59_port, temp00_58_port, temp00_57_port, temp00_56_port, 
      temp00_55_port, temp00_54_port, temp00_53_port, temp00_52_port, 
      temp00_51_port, temp00_50_port, temp00_49_port, temp00_48_port, 
      temp00_47_port, temp00_46_port, temp00_45_port, temp00_44_port, 
      temp00_43_port, temp00_42_port, temp00_41_port, temp00_40_port, 
      temp00_39_port, temp00_38_port, temp00_37_port, temp00_36_port, 
      temp00_35_port, temp00_34_port, temp00_33_port, temp00_32_port, 
      temp00_31_port, temp00_30_port, temp00_29_port, temp00_28_port, 
      temp00_27_port, temp00_26_port, temp00_25_port, temp00_24_port, 
      temp00_23_port, temp00_22_port, temp00_21_port, temp00_20_port, 
      temp00_19_port, temp00_18_port, temp00_17_port, temp00_16_port, 
      temp00_15_port, temp00_14_port, temp00_13_port, temp00_12_port, 
      temp00_11_port, temp00_10_port, temp00_9_port, temp00_8_port, 
      temp00_7_port, temp00_6_port, temp00_5_port, temp00_4_port, temp00_3_port
      , temp00_2_port, temp00_1_port, temp00_0_port, temp01_63_port, 
      temp01_62_port, temp01_61_port, temp01_60_port, temp01_59_port, 
      temp01_58_port, temp01_57_port, temp01_56_port, temp01_55_port, 
      temp01_54_port, temp01_53_port, temp01_52_port, temp01_51_port, 
      temp01_50_port, temp01_49_port, temp01_48_port, temp01_47_port, 
      temp01_46_port, temp01_45_port, temp01_44_port, temp01_43_port, 
      temp01_42_port, temp01_41_port, temp01_40_port, temp01_39_port, 
      temp01_38_port, temp01_37_port, temp01_36_port, temp01_35_port, 
      temp01_34_port, temp01_33_port, temp01_32_port, temp01_31_port, 
      temp01_30_port, temp01_29_port, temp01_28_port, temp01_27_port, 
      temp01_26_port, temp01_25_port, temp01_24_port, temp01_23_port, 
      temp01_22_port, temp01_21_port, temp01_20_port, temp01_19_port, 
      temp01_18_port, temp01_17_port, temp01_16_port, temp01_15_port, 
      temp01_14_port, temp01_13_port, temp01_12_port, temp01_11_port, 
      temp01_10_port, temp01_9_port, temp01_8_port, temp01_7_port, 
      temp01_6_port, temp01_5_port, temp01_4_port, temp01_3_port, temp01_2_port
      , temp01_1_port, temp01_0_port, temp1_63_port, temp1_62_port, 
      temp1_61_port, temp1_60_port, temp1_59_port, temp1_58_port, temp1_57_port
      , temp1_56_port, temp1_55_port, temp1_54_port, temp1_53_port, 
      temp1_52_port, temp1_51_port, temp1_50_port, temp1_49_port, temp1_48_port
      , temp1_47_port, temp1_46_port, temp1_45_port, temp1_44_port, 
      temp1_43_port, temp1_42_port, temp1_41_port, temp1_40_port, temp1_39_port
      , temp1_38_port, temp1_37_port, temp1_36_port, temp1_35_port, 
      temp1_34_port, temp1_33_port, temp1_32_port, temp1_31_port, temp1_30_port
      , temp1_29_port, temp1_28_port, temp1_27_port, temp1_26_port, 
      temp1_25_port, temp1_24_port, temp1_23_port, temp1_22_port, temp1_21_port
      , temp1_20_port, temp1_19_port, temp1_18_port, temp1_17_port, 
      temp1_16_port, temp1_15_port, temp1_14_port, temp1_13_port, temp1_12_port
      , temp1_11_port, temp1_10_port, temp1_9_port, temp1_8_port, temp1_7_port,
      temp1_6_port, temp1_5_port, temp1_4_port, temp1_3_port, temp1_2_port, 
      temp1_1_port, temp1_0_port : std_logic;

begin
   
   mux00 : MUX21_GENERIC_NBIT64_0 port map( A(63) => IN2(63), A(62) => IN2(62),
                           A(61) => IN2(61), A(60) => IN2(60), A(59) => IN2(59)
                           , A(58) => IN2(58), A(57) => IN2(57), A(56) => 
                           IN2(56), A(55) => IN2(55), A(54) => IN2(54), A(53) 
                           => IN2(53), A(52) => IN2(52), A(51) => IN2(51), 
                           A(50) => IN2(50), A(49) => IN2(49), A(48) => IN2(48)
                           , A(47) => IN2(47), A(46) => IN2(46), A(45) => 
                           IN2(45), A(44) => IN2(44), A(43) => IN2(43), A(42) 
                           => IN2(42), A(41) => IN2(41), A(40) => IN2(40), 
                           A(39) => IN2(39), A(38) => IN2(38), A(37) => IN2(37)
                           , A(36) => IN2(36), A(35) => IN2(35), A(34) => 
                           IN2(34), A(33) => IN2(33), A(32) => IN2(32), A(31) 
                           => IN2(31), A(30) => IN2(30), A(29) => IN2(29), 
                           A(28) => IN2(28), A(27) => IN2(27), A(26) => IN2(26)
                           , A(25) => IN2(25), A(24) => IN2(24), A(23) => 
                           IN2(23), A(22) => IN2(22), A(21) => IN2(21), A(20) 
                           => IN2(20), A(19) => IN2(19), A(18) => IN2(18), 
                           A(17) => IN2(17), A(16) => IN2(16), A(15) => IN2(15)
                           , A(14) => IN2(14), A(13) => IN2(13), A(12) => 
                           IN2(12), A(11) => IN2(11), A(10) => IN2(10), A(9) =>
                           IN2(9), A(8) => IN2(8), A(7) => IN2(7), A(6) => 
                           IN2(6), A(5) => IN2(5), A(4) => IN2(4), A(3) => 
                           IN2(3), A(2) => IN2(2), A(1) => IN2(1), A(0) => 
                           IN2(0), B(63) => IN1(63), B(62) => IN1(62), B(61) =>
                           IN1(61), B(60) => IN1(60), B(59) => IN1(59), B(58) 
                           => IN1(58), B(57) => IN1(57), B(56) => IN1(56), 
                           B(55) => IN1(55), B(54) => IN1(54), B(53) => IN1(53)
                           , B(52) => IN1(52), B(51) => IN1(51), B(50) => 
                           IN1(50), B(49) => IN1(49), B(48) => IN1(48), B(47) 
                           => IN1(47), B(46) => IN1(46), B(45) => IN1(45), 
                           B(44) => IN1(44), B(43) => IN1(43), B(42) => IN1(42)
                           , B(41) => IN1(41), B(40) => IN1(40), B(39) => 
                           IN1(39), B(38) => IN1(38), B(37) => IN1(37), B(36) 
                           => IN1(36), B(35) => IN1(35), B(34) => IN1(34), 
                           B(33) => IN1(33), B(32) => IN1(32), B(31) => IN1(31)
                           , B(30) => IN1(30), B(29) => IN1(29), B(28) => 
                           IN1(28), B(27) => IN1(27), B(26) => IN1(26), B(25) 
                           => IN1(25), B(24) => IN1(24), B(23) => IN1(23), 
                           B(22) => IN1(22), B(21) => IN1(21), B(20) => IN1(20)
                           , B(19) => IN1(19), B(18) => IN1(18), B(17) => 
                           IN1(17), B(16) => IN1(16), B(15) => IN1(15), B(14) 
                           => IN1(14), B(13) => IN1(13), B(12) => IN1(12), 
                           B(11) => IN1(11), B(10) => IN1(10), B(9) => IN1(9), 
                           B(8) => IN1(8), B(7) => IN1(7), B(6) => IN1(6), B(5)
                           => IN1(5), B(4) => IN1(4), B(3) => IN1(3), B(2) => 
                           IN1(2), B(1) => IN1(1), B(0) => IN1(0), SEL => S(0),
                           Y(63) => temp00_63_port, Y(62) => temp00_62_port, 
                           Y(61) => temp00_61_port, Y(60) => temp00_60_port, 
                           Y(59) => temp00_59_port, Y(58) => temp00_58_port, 
                           Y(57) => temp00_57_port, Y(56) => temp00_56_port, 
                           Y(55) => temp00_55_port, Y(54) => temp00_54_port, 
                           Y(53) => temp00_53_port, Y(52) => temp00_52_port, 
                           Y(51) => temp00_51_port, Y(50) => temp00_50_port, 
                           Y(49) => temp00_49_port, Y(48) => temp00_48_port, 
                           Y(47) => temp00_47_port, Y(46) => temp00_46_port, 
                           Y(45) => temp00_45_port, Y(44) => temp00_44_port, 
                           Y(43) => temp00_43_port, Y(42) => temp00_42_port, 
                           Y(41) => temp00_41_port, Y(40) => temp00_40_port, 
                           Y(39) => temp00_39_port, Y(38) => temp00_38_port, 
                           Y(37) => temp00_37_port, Y(36) => temp00_36_port, 
                           Y(35) => temp00_35_port, Y(34) => temp00_34_port, 
                           Y(33) => temp00_33_port, Y(32) => temp00_32_port, 
                           Y(31) => temp00_31_port, Y(30) => temp00_30_port, 
                           Y(29) => temp00_29_port, Y(28) => temp00_28_port, 
                           Y(27) => temp00_27_port, Y(26) => temp00_26_port, 
                           Y(25) => temp00_25_port, Y(24) => temp00_24_port, 
                           Y(23) => temp00_23_port, Y(22) => temp00_22_port, 
                           Y(21) => temp00_21_port, Y(20) => temp00_20_port, 
                           Y(19) => temp00_19_port, Y(18) => temp00_18_port, 
                           Y(17) => temp00_17_port, Y(16) => temp00_16_port, 
                           Y(15) => temp00_15_port, Y(14) => temp00_14_port, 
                           Y(13) => temp00_13_port, Y(12) => temp00_12_port, 
                           Y(11) => temp00_11_port, Y(10) => temp00_10_port, 
                           Y(9) => temp00_9_port, Y(8) => temp00_8_port, Y(7) 
                           => temp00_7_port, Y(6) => temp00_6_port, Y(5) => 
                           temp00_5_port, Y(4) => temp00_4_port, Y(3) => 
                           temp00_3_port, Y(2) => temp00_2_port, Y(1) => 
                           temp00_1_port, Y(0) => temp00_0_port);
   mux01 : MUX21_GENERIC_NBIT64_63 port map( A(63) => IN4(63), A(62) => IN4(62)
                           , A(61) => IN4(61), A(60) => IN4(60), A(59) => 
                           IN4(59), A(58) => IN4(58), A(57) => IN4(57), A(56) 
                           => IN4(56), A(55) => IN4(55), A(54) => IN4(54), 
                           A(53) => IN4(53), A(52) => IN4(52), A(51) => IN4(51)
                           , A(50) => IN4(50), A(49) => IN4(49), A(48) => 
                           IN4(48), A(47) => IN4(47), A(46) => IN4(46), A(45) 
                           => IN4(45), A(44) => IN4(44), A(43) => IN4(43), 
                           A(42) => IN4(42), A(41) => IN4(41), A(40) => IN4(40)
                           , A(39) => IN4(39), A(38) => IN4(38), A(37) => 
                           IN4(37), A(36) => IN4(36), A(35) => IN4(35), A(34) 
                           => IN4(34), A(33) => IN4(33), A(32) => IN4(32), 
                           A(31) => IN4(31), A(30) => IN4(30), A(29) => IN4(29)
                           , A(28) => IN4(28), A(27) => IN4(27), A(26) => 
                           IN4(26), A(25) => IN4(25), A(24) => IN4(24), A(23) 
                           => IN4(23), A(22) => IN4(22), A(21) => IN4(21), 
                           A(20) => IN4(20), A(19) => IN4(19), A(18) => IN4(18)
                           , A(17) => IN4(17), A(16) => IN4(16), A(15) => 
                           IN4(15), A(14) => IN4(14), A(13) => IN4(13), A(12) 
                           => IN4(12), A(11) => IN4(11), A(10) => IN4(10), A(9)
                           => IN4(9), A(8) => IN4(8), A(7) => IN4(7), A(6) => 
                           IN4(6), A(5) => IN4(5), A(4) => IN4(4), A(3) => 
                           IN4(3), A(2) => IN4(2), A(1) => IN4(1), A(0) => 
                           IN4(0), B(63) => IN3(63), B(62) => IN3(62), B(61) =>
                           IN3(61), B(60) => IN3(60), B(59) => IN3(59), B(58) 
                           => IN3(58), B(57) => IN3(57), B(56) => IN3(56), 
                           B(55) => IN3(55), B(54) => IN3(54), B(53) => IN3(53)
                           , B(52) => IN3(52), B(51) => IN3(51), B(50) => 
                           IN3(50), B(49) => IN3(49), B(48) => IN3(48), B(47) 
                           => IN3(47), B(46) => IN3(46), B(45) => IN3(45), 
                           B(44) => IN3(44), B(43) => IN3(43), B(42) => IN3(42)
                           , B(41) => IN3(41), B(40) => IN3(40), B(39) => 
                           IN3(39), B(38) => IN3(38), B(37) => IN3(37), B(36) 
                           => IN3(36), B(35) => IN3(35), B(34) => IN3(34), 
                           B(33) => IN3(33), B(32) => IN3(32), B(31) => IN3(31)
                           , B(30) => IN3(30), B(29) => IN3(29), B(28) => 
                           IN3(28), B(27) => IN3(27), B(26) => IN3(26), B(25) 
                           => IN3(25), B(24) => IN3(24), B(23) => IN3(23), 
                           B(22) => IN3(22), B(21) => IN3(21), B(20) => IN3(20)
                           , B(19) => IN3(19), B(18) => IN3(18), B(17) => 
                           IN3(17), B(16) => IN3(16), B(15) => IN3(15), B(14) 
                           => IN3(14), B(13) => IN3(13), B(12) => IN3(12), 
                           B(11) => IN3(11), B(10) => IN3(10), B(9) => IN3(9), 
                           B(8) => IN3(8), B(7) => IN3(7), B(6) => IN3(6), B(5)
                           => IN3(5), B(4) => IN3(4), B(3) => IN3(3), B(2) => 
                           IN3(2), B(1) => IN3(1), B(0) => IN3(0), SEL => S(0),
                           Y(63) => temp01_63_port, Y(62) => temp01_62_port, 
                           Y(61) => temp01_61_port, Y(60) => temp01_60_port, 
                           Y(59) => temp01_59_port, Y(58) => temp01_58_port, 
                           Y(57) => temp01_57_port, Y(56) => temp01_56_port, 
                           Y(55) => temp01_55_port, Y(54) => temp01_54_port, 
                           Y(53) => temp01_53_port, Y(52) => temp01_52_port, 
                           Y(51) => temp01_51_port, Y(50) => temp01_50_port, 
                           Y(49) => temp01_49_port, Y(48) => temp01_48_port, 
                           Y(47) => temp01_47_port, Y(46) => temp01_46_port, 
                           Y(45) => temp01_45_port, Y(44) => temp01_44_port, 
                           Y(43) => temp01_43_port, Y(42) => temp01_42_port, 
                           Y(41) => temp01_41_port, Y(40) => temp01_40_port, 
                           Y(39) => temp01_39_port, Y(38) => temp01_38_port, 
                           Y(37) => temp01_37_port, Y(36) => temp01_36_port, 
                           Y(35) => temp01_35_port, Y(34) => temp01_34_port, 
                           Y(33) => temp01_33_port, Y(32) => temp01_32_port, 
                           Y(31) => temp01_31_port, Y(30) => temp01_30_port, 
                           Y(29) => temp01_29_port, Y(28) => temp01_28_port, 
                           Y(27) => temp01_27_port, Y(26) => temp01_26_port, 
                           Y(25) => temp01_25_port, Y(24) => temp01_24_port, 
                           Y(23) => temp01_23_port, Y(22) => temp01_22_port, 
                           Y(21) => temp01_21_port, Y(20) => temp01_20_port, 
                           Y(19) => temp01_19_port, Y(18) => temp01_18_port, 
                           Y(17) => temp01_17_port, Y(16) => temp01_16_port, 
                           Y(15) => temp01_15_port, Y(14) => temp01_14_port, 
                           Y(13) => temp01_13_port, Y(12) => temp01_12_port, 
                           Y(11) => temp01_11_port, Y(10) => temp01_10_port, 
                           Y(9) => temp01_9_port, Y(8) => temp01_8_port, Y(7) 
                           => temp01_7_port, Y(6) => temp01_6_port, Y(5) => 
                           temp01_5_port, Y(4) => temp01_4_port, Y(3) => 
                           temp01_3_port, Y(2) => temp01_2_port, Y(1) => 
                           temp01_1_port, Y(0) => temp01_0_port);
   mux1 : MUX21_GENERIC_NBIT64_62 port map( A(63) => temp01_63_port, A(62) => 
                           temp01_62_port, A(61) => temp01_61_port, A(60) => 
                           temp01_60_port, A(59) => temp01_59_port, A(58) => 
                           temp01_58_port, A(57) => temp01_57_port, A(56) => 
                           temp01_56_port, A(55) => temp01_55_port, A(54) => 
                           temp01_54_port, A(53) => temp01_53_port, A(52) => 
                           temp01_52_port, A(51) => temp01_51_port, A(50) => 
                           temp01_50_port, A(49) => temp01_49_port, A(48) => 
                           temp01_48_port, A(47) => temp01_47_port, A(46) => 
                           temp01_46_port, A(45) => temp01_45_port, A(44) => 
                           temp01_44_port, A(43) => temp01_43_port, A(42) => 
                           temp01_42_port, A(41) => temp01_41_port, A(40) => 
                           temp01_40_port, A(39) => temp01_39_port, A(38) => 
                           temp01_38_port, A(37) => temp01_37_port, A(36) => 
                           temp01_36_port, A(35) => temp01_35_port, A(34) => 
                           temp01_34_port, A(33) => temp01_33_port, A(32) => 
                           temp01_32_port, A(31) => temp01_31_port, A(30) => 
                           temp01_30_port, A(29) => temp01_29_port, A(28) => 
                           temp01_28_port, A(27) => temp01_27_port, A(26) => 
                           temp01_26_port, A(25) => temp01_25_port, A(24) => 
                           temp01_24_port, A(23) => temp01_23_port, A(22) => 
                           temp01_22_port, A(21) => temp01_21_port, A(20) => 
                           temp01_20_port, A(19) => temp01_19_port, A(18) => 
                           temp01_18_port, A(17) => temp01_17_port, A(16) => 
                           temp01_16_port, A(15) => temp01_15_port, A(14) => 
                           temp01_14_port, A(13) => temp01_13_port, A(12) => 
                           temp01_12_port, A(11) => temp01_11_port, A(10) => 
                           temp01_10_port, A(9) => temp01_9_port, A(8) => 
                           temp01_8_port, A(7) => temp01_7_port, A(6) => 
                           temp01_6_port, A(5) => temp01_5_port, A(4) => 
                           temp01_4_port, A(3) => temp01_3_port, A(2) => 
                           temp01_2_port, A(1) => temp01_1_port, A(0) => 
                           temp01_0_port, B(63) => temp00_63_port, B(62) => 
                           temp00_62_port, B(61) => temp00_61_port, B(60) => 
                           temp00_60_port, B(59) => temp00_59_port, B(58) => 
                           temp00_58_port, B(57) => temp00_57_port, B(56) => 
                           temp00_56_port, B(55) => temp00_55_port, B(54) => 
                           temp00_54_port, B(53) => temp00_53_port, B(52) => 
                           temp00_52_port, B(51) => temp00_51_port, B(50) => 
                           temp00_50_port, B(49) => temp00_49_port, B(48) => 
                           temp00_48_port, B(47) => temp00_47_port, B(46) => 
                           temp00_46_port, B(45) => temp00_45_port, B(44) => 
                           temp00_44_port, B(43) => temp00_43_port, B(42) => 
                           temp00_42_port, B(41) => temp00_41_port, B(40) => 
                           temp00_40_port, B(39) => temp00_39_port, B(38) => 
                           temp00_38_port, B(37) => temp00_37_port, B(36) => 
                           temp00_36_port, B(35) => temp00_35_port, B(34) => 
                           temp00_34_port, B(33) => temp00_33_port, B(32) => 
                           temp00_32_port, B(31) => temp00_31_port, B(30) => 
                           temp00_30_port, B(29) => temp00_29_port, B(28) => 
                           temp00_28_port, B(27) => temp00_27_port, B(26) => 
                           temp00_26_port, B(25) => temp00_25_port, B(24) => 
                           temp00_24_port, B(23) => temp00_23_port, B(22) => 
                           temp00_22_port, B(21) => temp00_21_port, B(20) => 
                           temp00_20_port, B(19) => temp00_19_port, B(18) => 
                           temp00_18_port, B(17) => temp00_17_port, B(16) => 
                           temp00_16_port, B(15) => temp00_15_port, B(14) => 
                           temp00_14_port, B(13) => temp00_13_port, B(12) => 
                           temp00_12_port, B(11) => temp00_11_port, B(10) => 
                           temp00_10_port, B(9) => temp00_9_port, B(8) => 
                           temp00_8_port, B(7) => temp00_7_port, B(6) => 
                           temp00_6_port, B(5) => temp00_5_port, B(4) => 
                           temp00_4_port, B(3) => temp00_3_port, B(2) => 
                           temp00_2_port, B(1) => temp00_1_port, B(0) => 
                           temp00_0_port, SEL => S(1), Y(63) => temp1_63_port, 
                           Y(62) => temp1_62_port, Y(61) => temp1_61_port, 
                           Y(60) => temp1_60_port, Y(59) => temp1_59_port, 
                           Y(58) => temp1_58_port, Y(57) => temp1_57_port, 
                           Y(56) => temp1_56_port, Y(55) => temp1_55_port, 
                           Y(54) => temp1_54_port, Y(53) => temp1_53_port, 
                           Y(52) => temp1_52_port, Y(51) => temp1_51_port, 
                           Y(50) => temp1_50_port, Y(49) => temp1_49_port, 
                           Y(48) => temp1_48_port, Y(47) => temp1_47_port, 
                           Y(46) => temp1_46_port, Y(45) => temp1_45_port, 
                           Y(44) => temp1_44_port, Y(43) => temp1_43_port, 
                           Y(42) => temp1_42_port, Y(41) => temp1_41_port, 
                           Y(40) => temp1_40_port, Y(39) => temp1_39_port, 
                           Y(38) => temp1_38_port, Y(37) => temp1_37_port, 
                           Y(36) => temp1_36_port, Y(35) => temp1_35_port, 
                           Y(34) => temp1_34_port, Y(33) => temp1_33_port, 
                           Y(32) => temp1_32_port, Y(31) => temp1_31_port, 
                           Y(30) => temp1_30_port, Y(29) => temp1_29_port, 
                           Y(28) => temp1_28_port, Y(27) => temp1_27_port, 
                           Y(26) => temp1_26_port, Y(25) => temp1_25_port, 
                           Y(24) => temp1_24_port, Y(23) => temp1_23_port, 
                           Y(22) => temp1_22_port, Y(21) => temp1_21_port, 
                           Y(20) => temp1_20_port, Y(19) => temp1_19_port, 
                           Y(18) => temp1_18_port, Y(17) => temp1_17_port, 
                           Y(16) => temp1_16_port, Y(15) => temp1_15_port, 
                           Y(14) => temp1_14_port, Y(13) => temp1_13_port, 
                           Y(12) => temp1_12_port, Y(11) => temp1_11_port, 
                           Y(10) => temp1_10_port, Y(9) => temp1_9_port, Y(8) 
                           => temp1_8_port, Y(7) => temp1_7_port, Y(6) => 
                           temp1_6_port, Y(5) => temp1_5_port, Y(4) => 
                           temp1_4_port, Y(3) => temp1_3_port, Y(2) => 
                           temp1_2_port, Y(1) => temp1_1_port, Y(0) => 
                           temp1_0_port);
   mux2 : MUX21_GENERIC_NBIT64_61 port map( A(63) => IN0(63), A(62) => IN0(62),
                           A(61) => IN0(61), A(60) => IN0(60), A(59) => IN0(59)
                           , A(58) => IN0(58), A(57) => IN0(57), A(56) => 
                           IN0(56), A(55) => IN0(55), A(54) => IN0(54), A(53) 
                           => IN0(53), A(52) => IN0(52), A(51) => IN0(51), 
                           A(50) => IN0(50), A(49) => IN0(49), A(48) => IN0(48)
                           , A(47) => IN0(47), A(46) => IN0(46), A(45) => 
                           IN0(45), A(44) => IN0(44), A(43) => IN0(43), A(42) 
                           => IN0(42), A(41) => IN0(41), A(40) => IN0(40), 
                           A(39) => IN0(39), A(38) => IN0(38), A(37) => IN0(37)
                           , A(36) => IN0(36), A(35) => IN0(35), A(34) => 
                           IN0(34), A(33) => IN0(33), A(32) => IN0(32), A(31) 
                           => IN0(31), A(30) => IN0(30), A(29) => IN0(29), 
                           A(28) => IN0(28), A(27) => IN0(27), A(26) => IN0(26)
                           , A(25) => IN0(25), A(24) => IN0(24), A(23) => 
                           IN0(23), A(22) => IN0(22), A(21) => IN0(21), A(20) 
                           => IN0(20), A(19) => IN0(19), A(18) => IN0(18), 
                           A(17) => IN0(17), A(16) => IN0(16), A(15) => IN0(15)
                           , A(14) => IN0(14), A(13) => IN0(13), A(12) => 
                           IN0(12), A(11) => IN0(11), A(10) => IN0(10), A(9) =>
                           IN0(9), A(8) => IN0(8), A(7) => IN0(7), A(6) => 
                           IN0(6), A(5) => IN0(5), A(4) => IN0(4), A(3) => 
                           IN0(3), A(2) => IN0(2), A(1) => IN0(1), A(0) => 
                           IN0(0), B(63) => temp1_63_port, B(62) => 
                           temp1_62_port, B(61) => temp1_61_port, B(60) => 
                           temp1_60_port, B(59) => temp1_59_port, B(58) => 
                           temp1_58_port, B(57) => temp1_57_port, B(56) => 
                           temp1_56_port, B(55) => temp1_55_port, B(54) => 
                           temp1_54_port, B(53) => temp1_53_port, B(52) => 
                           temp1_52_port, B(51) => temp1_51_port, B(50) => 
                           temp1_50_port, B(49) => temp1_49_port, B(48) => 
                           temp1_48_port, B(47) => temp1_47_port, B(46) => 
                           temp1_46_port, B(45) => temp1_45_port, B(44) => 
                           temp1_44_port, B(43) => temp1_43_port, B(42) => 
                           temp1_42_port, B(41) => temp1_41_port, B(40) => 
                           temp1_40_port, B(39) => temp1_39_port, B(38) => 
                           temp1_38_port, B(37) => temp1_37_port, B(36) => 
                           temp1_36_port, B(35) => temp1_35_port, B(34) => 
                           temp1_34_port, B(33) => temp1_33_port, B(32) => 
                           temp1_32_port, B(31) => temp1_31_port, B(30) => 
                           temp1_30_port, B(29) => temp1_29_port, B(28) => 
                           temp1_28_port, B(27) => temp1_27_port, B(26) => 
                           temp1_26_port, B(25) => temp1_25_port, B(24) => 
                           temp1_24_port, B(23) => temp1_23_port, B(22) => 
                           temp1_22_port, B(21) => temp1_21_port, B(20) => 
                           temp1_20_port, B(19) => temp1_19_port, B(18) => 
                           temp1_18_port, B(17) => temp1_17_port, B(16) => 
                           temp1_16_port, B(15) => temp1_15_port, B(14) => 
                           temp1_14_port, B(13) => temp1_13_port, B(12) => 
                           temp1_12_port, B(11) => temp1_11_port, B(10) => 
                           temp1_10_port, B(9) => temp1_9_port, B(8) => 
                           temp1_8_port, B(7) => temp1_7_port, B(6) => 
                           temp1_6_port, B(5) => temp1_5_port, B(4) => 
                           temp1_4_port, B(3) => temp1_3_port, B(2) => 
                           temp1_2_port, B(1) => temp1_1_port, B(0) => 
                           temp1_0_port, SEL => S(2), Y(63) => O(63), Y(62) => 
                           O(62), Y(61) => O(61), Y(60) => O(60), Y(59) => 
                           O(59), Y(58) => O(58), Y(57) => O(57), Y(56) => 
                           O(56), Y(55) => O(55), Y(54) => O(54), Y(53) => 
                           O(53), Y(52) => O(52), Y(51) => O(51), Y(50) => 
                           O(50), Y(49) => O(49), Y(48) => O(48), Y(47) => 
                           O(47), Y(46) => O(46), Y(45) => O(45), Y(44) => 
                           O(44), Y(43) => O(43), Y(42) => O(42), Y(41) => 
                           O(41), Y(40) => O(40), Y(39) => O(39), Y(38) => 
                           O(38), Y(37) => O(37), Y(36) => O(36), Y(35) => 
                           O(35), Y(34) => O(34), Y(33) => O(33), Y(32) => 
                           O(32), Y(31) => O(31), Y(30) => O(30), Y(29) => 
                           O(29), Y(28) => O(28), Y(27) => O(27), Y(26) => 
                           O(26), Y(25) => O(25), Y(24) => O(24), Y(23) => 
                           O(23), Y(22) => O(22), Y(21) => O(21), Y(20) => 
                           O(20), Y(19) => O(19), Y(18) => O(18), Y(17) => 
                           O(17), Y(16) => O(16), Y(15) => O(15), Y(14) => 
                           O(14), Y(13) => O(13), Y(12) => O(12), Y(11) => 
                           O(11), Y(10) => O(10), Y(9) => O(9), Y(8) => O(8), 
                           Y(7) => O(7), Y(6) => O(6), Y(5) => O(5), Y(4) => 
                           O(4), Y(3) => O(3), Y(2) => O(2), Y(1) => O(1), Y(0)
                           => O(0));

end SYN_mux51_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTH_ENCODER_3BIT_4 is

   port( B : in std_logic_vector (2 downto 0);  ENCODED : out std_logic_vector 
         (2 downto 0));

end BOOTH_ENCODER_3BIT_4;

architecture SYN_dataflow of BOOTH_ENCODER_3BIT_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U3 : INV_X4 port map( A => n1, ZN => ENCODED(1));
   U4 : NAND2_X4 port map( A1 => n2, A2 => n1, ZN => ENCODED(2));
   U5 : XOR2_X1 port map( A => n3, B => B(2), Z => n2);
   U6 : AOI21_X1 port map( B1 => n1, B2 => n3, A => B(2), ZN => ENCODED(0));
   U7 : XOR2_X1 port map( A => n3, B => B(1), Z => n1);
   U8 : INV_X1 port map( A => B(0), ZN => n3);

end SYN_dataflow;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHMUL_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  P : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL_NBIT32;

architecture SYN_BOOTHMUL_STRUCT of BOOTHMUL_NBIT32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BOOTHMUL_NBIT32_DW01_inc_0
      port( A : in std_logic_vector (63 downto 0);  SUM : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_1
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_1
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_5
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_2
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_2
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_6
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_3
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_3
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_7
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_4
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_4
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_8
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_5
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_5
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_9
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_6
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_6
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_10
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_7
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_7
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_11
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_8
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_8
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_12
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_9
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_9
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_13
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_10
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_10
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_14
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_11
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_11
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_15
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_12
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_12
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_16
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_13
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_13
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_17
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_14
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_14
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_18
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT64_0
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT64_15
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_19
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component MUX51_GENERIC_NBIT64_0
      port( IN0, IN1, IN2, IN3, IN4 : in std_logic_vector (63 downto 0);  S : 
            in std_logic_vector (2 downto 0);  O : out std_logic_vector (63 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_3BIT_4
      port( B : in std_logic_vector (2 downto 0);  ENCODED : out 
            std_logic_vector (2 downto 0));
   end component;
   
   signal X_Logic0_port, negative_a_63_port, negative_a_62_port, 
      negative_a_61_port, negative_a_60_port, negative_a_59_port, 
      negative_a_58_port, negative_a_57_port, negative_a_56_port, 
      negative_a_55_port, negative_a_54_port, negative_a_53_port, 
      negative_a_52_port, negative_a_51_port, negative_a_50_port, 
      negative_a_49_port, negative_a_48_port, negative_a_47_port, 
      negative_a_46_port, negative_a_45_port, negative_a_44_port, 
      negative_a_43_port, negative_a_42_port, negative_a_41_port, 
      negative_a_40_port, negative_a_39_port, negative_a_38_port, 
      negative_a_37_port, negative_a_36_port, negative_a_35_port, 
      negative_a_34_port, negative_a_33_port, negative_a_32_port, 
      negative_a_31_port, negative_a_30_port, negative_a_29_port, 
      negative_a_28_port, negative_a_27_port, negative_a_26_port, 
      negative_a_25_port, negative_a_24_port, negative_a_23_port, 
      negative_a_22_port, negative_a_21_port, negative_a_20_port, 
      negative_a_19_port, negative_a_18_port, negative_a_17_port, 
      negative_a_16_port, negative_a_15_port, negative_a_14_port, 
      negative_a_13_port, negative_a_12_port, negative_a_11_port, 
      negative_a_10_port, negative_a_9_port, negative_a_8_port, 
      negative_a_7_port, negative_a_6_port, negative_a_5_port, 
      negative_a_4_port, negative_a_3_port, negative_a_2_port, 
      negative_a_1_port, negative_a_0_port, muxs_encoded_signals_0_2_port, 
      muxs_encoded_signals_0_1_port, muxs_encoded_signals_0_0_port, 
      muxs_encoded_signals_1_2_port, muxs_encoded_signals_1_1_port, 
      muxs_encoded_signals_1_0_port, muxs_encoded_signals_2_2_port, 
      muxs_encoded_signals_2_1_port, muxs_encoded_signals_2_0_port, 
      muxs_encoded_signals_3_2_port, muxs_encoded_signals_3_1_port, 
      muxs_encoded_signals_3_0_port, muxs_encoded_signals_4_2_port, 
      muxs_encoded_signals_4_1_port, muxs_encoded_signals_4_0_port, 
      muxs_encoded_signals_5_2_port, muxs_encoded_signals_5_1_port, 
      muxs_encoded_signals_5_0_port, muxs_encoded_signals_6_2_port, 
      muxs_encoded_signals_6_1_port, muxs_encoded_signals_6_0_port, 
      muxs_encoded_signals_7_2_port, muxs_encoded_signals_7_1_port, 
      muxs_encoded_signals_7_0_port, muxs_encoded_signals_8_2_port, 
      muxs_encoded_signals_8_1_port, muxs_encoded_signals_8_0_port, 
      muxs_encoded_signals_9_2_port, muxs_encoded_signals_9_1_port, 
      muxs_encoded_signals_9_0_port, muxs_encoded_signals_10_2_port, 
      muxs_encoded_signals_10_1_port, muxs_encoded_signals_10_0_port, 
      muxs_encoded_signals_11_2_port, muxs_encoded_signals_11_1_port, 
      muxs_encoded_signals_11_0_port, muxs_encoded_signals_12_2_port, 
      muxs_encoded_signals_12_1_port, muxs_encoded_signals_12_0_port, 
      muxs_encoded_signals_13_2_port, muxs_encoded_signals_13_1_port, 
      muxs_encoded_signals_13_0_port, muxs_encoded_signals_14_2_port, 
      muxs_encoded_signals_14_1_port, muxs_encoded_signals_14_0_port, 
      muxs_encoded_signals_15_2_port, muxs_encoded_signals_15_1_port, 
      muxs_encoded_signals_15_0_port, out_imux_0_63_port, out_imux_0_62_port, 
      out_imux_0_61_port, out_imux_0_60_port, out_imux_0_59_port, 
      out_imux_0_58_port, out_imux_0_57_port, out_imux_0_56_port, 
      out_imux_0_55_port, out_imux_0_54_port, out_imux_0_53_port, 
      out_imux_0_52_port, out_imux_0_51_port, out_imux_0_50_port, 
      out_imux_0_49_port, out_imux_0_48_port, out_imux_0_47_port, 
      out_imux_0_46_port, out_imux_0_45_port, out_imux_0_44_port, 
      out_imux_0_43_port, out_imux_0_42_port, out_imux_0_41_port, 
      out_imux_0_40_port, out_imux_0_39_port, out_imux_0_38_port, 
      out_imux_0_37_port, out_imux_0_36_port, out_imux_0_35_port, 
      out_imux_0_34_port, out_imux_0_33_port, out_imux_0_32_port, 
      out_imux_0_31_port, out_imux_0_30_port, out_imux_0_29_port, 
      out_imux_0_28_port, out_imux_0_27_port, out_imux_0_26_port, 
      out_imux_0_25_port, out_imux_0_24_port, out_imux_0_23_port, 
      out_imux_0_22_port, out_imux_0_21_port, out_imux_0_20_port, 
      out_imux_0_19_port, out_imux_0_18_port, out_imux_0_17_port, 
      out_imux_0_16_port, out_imux_0_15_port, out_imux_0_14_port, 
      out_imux_0_13_port, out_imux_0_12_port, out_imux_0_11_port, 
      out_imux_0_10_port, out_imux_0_9_port, out_imux_0_8_port, 
      out_imux_0_7_port, out_imux_0_6_port, out_imux_0_5_port, 
      out_imux_0_4_port, out_imux_0_3_port, out_imux_0_2_port, 
      out_imux_0_1_port, out_imux_0_0_port, out_imux_1_63_port, 
      out_imux_1_62_port, out_imux_1_61_port, out_imux_1_60_port, 
      out_imux_1_59_port, out_imux_1_58_port, out_imux_1_57_port, 
      out_imux_1_56_port, out_imux_1_55_port, out_imux_1_54_port, 
      out_imux_1_53_port, out_imux_1_52_port, out_imux_1_51_port, 
      out_imux_1_50_port, out_imux_1_49_port, out_imux_1_48_port, 
      out_imux_1_47_port, out_imux_1_46_port, out_imux_1_45_port, 
      out_imux_1_44_port, out_imux_1_43_port, out_imux_1_42_port, 
      out_imux_1_41_port, out_imux_1_40_port, out_imux_1_39_port, 
      out_imux_1_38_port, out_imux_1_37_port, out_imux_1_36_port, 
      out_imux_1_35_port, out_imux_1_34_port, out_imux_1_33_port, 
      out_imux_1_32_port, out_imux_1_31_port, out_imux_1_30_port, 
      out_imux_1_29_port, out_imux_1_28_port, out_imux_1_27_port, 
      out_imux_1_26_port, out_imux_1_25_port, out_imux_1_24_port, 
      out_imux_1_23_port, out_imux_1_22_port, out_imux_1_21_port, 
      out_imux_1_20_port, out_imux_1_19_port, out_imux_1_18_port, 
      out_imux_1_17_port, out_imux_1_16_port, out_imux_1_15_port, 
      out_imux_1_14_port, out_imux_1_13_port, out_imux_1_12_port, 
      out_imux_1_11_port, out_imux_1_10_port, out_imux_1_9_port, 
      out_imux_1_8_port, out_imux_1_7_port, out_imux_1_6_port, 
      out_imux_1_5_port, out_imux_1_4_port, out_imux_1_3_port, 
      out_imux_1_2_port, out_imux_1_1_port, out_imux_1_0_port, 
      out_imux_2_63_port, out_imux_2_62_port, out_imux_2_61_port, 
      out_imux_2_60_port, out_imux_2_59_port, out_imux_2_58_port, 
      out_imux_2_57_port, out_imux_2_56_port, out_imux_2_55_port, 
      out_imux_2_54_port, out_imux_2_53_port, out_imux_2_52_port, 
      out_imux_2_51_port, out_imux_2_50_port, out_imux_2_49_port, 
      out_imux_2_48_port, out_imux_2_47_port, out_imux_2_46_port, 
      out_imux_2_45_port, out_imux_2_44_port, out_imux_2_43_port, 
      out_imux_2_42_port, out_imux_2_41_port, out_imux_2_40_port, 
      out_imux_2_39_port, out_imux_2_38_port, out_imux_2_37_port, 
      out_imux_2_36_port, out_imux_2_35_port, out_imux_2_34_port, 
      out_imux_2_33_port, out_imux_2_32_port, out_imux_2_31_port, 
      out_imux_2_30_port, out_imux_2_29_port, out_imux_2_28_port, 
      out_imux_2_27_port, out_imux_2_26_port, out_imux_2_25_port, 
      out_imux_2_24_port, out_imux_2_23_port, out_imux_2_22_port, 
      out_imux_2_21_port, out_imux_2_20_port, out_imux_2_19_port, 
      out_imux_2_18_port, out_imux_2_17_port, out_imux_2_16_port, 
      out_imux_2_15_port, out_imux_2_14_port, out_imux_2_13_port, 
      out_imux_2_12_port, out_imux_2_11_port, out_imux_2_10_port, 
      out_imux_2_9_port, out_imux_2_8_port, out_imux_2_7_port, 
      out_imux_2_6_port, out_imux_2_5_port, out_imux_2_4_port, 
      out_imux_2_3_port, out_imux_2_2_port, out_imux_2_1_port, 
      out_imux_2_0_port, out_imux_3_63_port, out_imux_3_62_port, 
      out_imux_3_61_port, out_imux_3_60_port, out_imux_3_59_port, 
      out_imux_3_58_port, out_imux_3_57_port, out_imux_3_56_port, 
      out_imux_3_55_port, out_imux_3_54_port, out_imux_3_53_port, 
      out_imux_3_52_port, out_imux_3_51_port, out_imux_3_50_port, 
      out_imux_3_49_port, out_imux_3_48_port, out_imux_3_47_port, 
      out_imux_3_46_port, out_imux_3_45_port, out_imux_3_44_port, 
      out_imux_3_43_port, out_imux_3_42_port, out_imux_3_41_port, 
      out_imux_3_40_port, out_imux_3_39_port, out_imux_3_38_port, 
      out_imux_3_37_port, out_imux_3_36_port, out_imux_3_35_port, 
      out_imux_3_34_port, out_imux_3_33_port, out_imux_3_32_port, 
      out_imux_3_31_port, out_imux_3_30_port, out_imux_3_29_port, 
      out_imux_3_28_port, out_imux_3_27_port, out_imux_3_26_port, 
      out_imux_3_25_port, out_imux_3_24_port, out_imux_3_23_port, 
      out_imux_3_22_port, out_imux_3_21_port, out_imux_3_20_port, 
      out_imux_3_19_port, out_imux_3_18_port, out_imux_3_17_port, 
      out_imux_3_16_port, out_imux_3_15_port, out_imux_3_14_port, 
      out_imux_3_13_port, out_imux_3_12_port, out_imux_3_11_port, 
      out_imux_3_10_port, out_imux_3_9_port, out_imux_3_8_port, 
      out_imux_3_7_port, out_imux_3_6_port, out_imux_3_5_port, 
      out_imux_3_4_port, out_imux_3_3_port, out_imux_3_2_port, 
      out_imux_3_1_port, out_imux_3_0_port, out_imux_4_63_port, 
      out_imux_4_62_port, out_imux_4_61_port, out_imux_4_60_port, 
      out_imux_4_59_port, out_imux_4_58_port, out_imux_4_57_port, 
      out_imux_4_56_port, out_imux_4_55_port, out_imux_4_54_port, 
      out_imux_4_53_port, out_imux_4_52_port, out_imux_4_51_port, 
      out_imux_4_50_port, out_imux_4_49_port, out_imux_4_48_port, 
      out_imux_4_47_port, out_imux_4_46_port, out_imux_4_45_port, 
      out_imux_4_44_port, out_imux_4_43_port, out_imux_4_42_port, 
      out_imux_4_41_port, out_imux_4_40_port, out_imux_4_39_port, 
      out_imux_4_38_port, out_imux_4_37_port, out_imux_4_36_port, 
      out_imux_4_35_port, out_imux_4_34_port, out_imux_4_33_port, 
      out_imux_4_32_port, out_imux_4_31_port, out_imux_4_30_port, 
      out_imux_4_29_port, out_imux_4_28_port, out_imux_4_27_port, 
      out_imux_4_26_port, out_imux_4_25_port, out_imux_4_24_port, 
      out_imux_4_23_port, out_imux_4_22_port, out_imux_4_21_port, 
      out_imux_4_20_port, out_imux_4_19_port, out_imux_4_18_port, 
      out_imux_4_17_port, out_imux_4_16_port, out_imux_4_15_port, 
      out_imux_4_14_port, out_imux_4_13_port, out_imux_4_12_port, 
      out_imux_4_11_port, out_imux_4_10_port, out_imux_4_9_port, 
      out_imux_4_8_port, out_imux_4_7_port, out_imux_4_6_port, 
      out_imux_4_5_port, out_imux_4_4_port, out_imux_4_3_port, 
      out_imux_4_2_port, out_imux_4_1_port, out_imux_4_0_port, 
      out_imux_5_63_port, out_imux_5_62_port, out_imux_5_61_port, 
      out_imux_5_60_port, out_imux_5_59_port, out_imux_5_58_port, 
      out_imux_5_57_port, out_imux_5_56_port, out_imux_5_55_port, 
      out_imux_5_54_port, out_imux_5_53_port, out_imux_5_52_port, 
      out_imux_5_51_port, out_imux_5_50_port, out_imux_5_49_port, 
      out_imux_5_48_port, out_imux_5_47_port, out_imux_5_46_port, 
      out_imux_5_45_port, out_imux_5_44_port, out_imux_5_43_port, 
      out_imux_5_42_port, out_imux_5_41_port, out_imux_5_40_port, 
      out_imux_5_39_port, out_imux_5_38_port, out_imux_5_37_port, 
      out_imux_5_36_port, out_imux_5_35_port, out_imux_5_34_port, 
      out_imux_5_33_port, out_imux_5_32_port, out_imux_5_31_port, 
      out_imux_5_30_port, out_imux_5_29_port, out_imux_5_28_port, 
      out_imux_5_27_port, out_imux_5_26_port, out_imux_5_25_port, 
      out_imux_5_24_port, out_imux_5_23_port, out_imux_5_22_port, 
      out_imux_5_21_port, out_imux_5_20_port, out_imux_5_19_port, 
      out_imux_5_18_port, out_imux_5_17_port, out_imux_5_16_port, 
      out_imux_5_15_port, out_imux_5_14_port, out_imux_5_13_port, 
      out_imux_5_12_port, out_imux_5_11_port, out_imux_5_10_port, 
      out_imux_5_9_port, out_imux_5_8_port, out_imux_5_7_port, 
      out_imux_5_6_port, out_imux_5_5_port, out_imux_5_4_port, 
      out_imux_5_3_port, out_imux_5_2_port, out_imux_5_1_port, 
      out_imux_5_0_port, out_imux_6_63_port, out_imux_6_62_port, 
      out_imux_6_61_port, out_imux_6_60_port, out_imux_6_59_port, 
      out_imux_6_58_port, out_imux_6_57_port, out_imux_6_56_port, 
      out_imux_6_55_port, out_imux_6_54_port, out_imux_6_53_port, 
      out_imux_6_52_port, out_imux_6_51_port, out_imux_6_50_port, 
      out_imux_6_49_port, out_imux_6_48_port, out_imux_6_47_port, 
      out_imux_6_46_port, out_imux_6_45_port, out_imux_6_44_port, 
      out_imux_6_43_port, out_imux_6_42_port, out_imux_6_41_port, 
      out_imux_6_40_port, out_imux_6_39_port, out_imux_6_38_port, 
      out_imux_6_37_port, out_imux_6_36_port, out_imux_6_35_port, 
      out_imux_6_34_port, out_imux_6_33_port, out_imux_6_32_port, 
      out_imux_6_31_port, out_imux_6_30_port, out_imux_6_29_port, 
      out_imux_6_28_port, out_imux_6_27_port, out_imux_6_26_port, 
      out_imux_6_25_port, out_imux_6_24_port, out_imux_6_23_port, 
      out_imux_6_22_port, out_imux_6_21_port, out_imux_6_20_port, 
      out_imux_6_19_port, out_imux_6_18_port, out_imux_6_17_port, 
      out_imux_6_16_port, out_imux_6_15_port, out_imux_6_14_port, 
      out_imux_6_13_port, out_imux_6_12_port, out_imux_6_11_port, 
      out_imux_6_10_port, out_imux_6_9_port, out_imux_6_8_port, 
      out_imux_6_7_port, out_imux_6_6_port, out_imux_6_5_port, 
      out_imux_6_4_port, out_imux_6_3_port, out_imux_6_2_port, 
      out_imux_6_1_port, out_imux_6_0_port, out_imux_7_63_port, 
      out_imux_7_62_port, out_imux_7_61_port, out_imux_7_60_port, 
      out_imux_7_59_port, out_imux_7_58_port, out_imux_7_57_port, 
      out_imux_7_56_port, out_imux_7_55_port, out_imux_7_54_port, 
      out_imux_7_53_port, out_imux_7_52_port, out_imux_7_51_port, 
      out_imux_7_50_port, out_imux_7_49_port, out_imux_7_48_port, 
      out_imux_7_47_port, out_imux_7_46_port, out_imux_7_45_port, 
      out_imux_7_44_port, out_imux_7_43_port, out_imux_7_42_port, 
      out_imux_7_41_port, out_imux_7_40_port, out_imux_7_39_port, 
      out_imux_7_38_port, out_imux_7_37_port, out_imux_7_36_port, 
      out_imux_7_35_port, out_imux_7_34_port, out_imux_7_33_port, 
      out_imux_7_32_port, out_imux_7_31_port, out_imux_7_30_port, 
      out_imux_7_29_port, out_imux_7_28_port, out_imux_7_27_port, 
      out_imux_7_26_port, out_imux_7_25_port, out_imux_7_24_port, 
      out_imux_7_23_port, out_imux_7_22_port, out_imux_7_21_port, 
      out_imux_7_20_port, out_imux_7_19_port, out_imux_7_18_port, 
      out_imux_7_17_port, out_imux_7_16_port, out_imux_7_15_port, 
      out_imux_7_14_port, out_imux_7_13_port, out_imux_7_12_port, 
      out_imux_7_11_port, out_imux_7_10_port, out_imux_7_9_port, 
      out_imux_7_8_port, out_imux_7_7_port, out_imux_7_6_port, 
      out_imux_7_5_port, out_imux_7_4_port, out_imux_7_3_port, 
      out_imux_7_2_port, out_imux_7_1_port, out_imux_7_0_port, 
      predigest_product_1_63_port, predigest_product_1_62_port, 
      predigest_product_1_61_port, predigest_product_1_60_port, 
      predigest_product_1_59_port, predigest_product_1_58_port, 
      predigest_product_1_57_port, predigest_product_1_56_port, 
      predigest_product_1_55_port, predigest_product_1_54_port, 
      predigest_product_1_53_port, predigest_product_1_52_port, 
      predigest_product_1_51_port, predigest_product_1_50_port, 
      predigest_product_1_49_port, predigest_product_1_48_port, 
      predigest_product_1_47_port, predigest_product_1_46_port, 
      predigest_product_1_45_port, predigest_product_1_44_port, 
      predigest_product_1_43_port, predigest_product_1_42_port, 
      predigest_product_1_41_port, predigest_product_1_40_port, 
      predigest_product_1_39_port, predigest_product_1_38_port, 
      predigest_product_1_37_port, predigest_product_1_36_port, 
      predigest_product_1_35_port, predigest_product_1_34_port, 
      predigest_product_1_33_port, predigest_product_1_32_port, 
      predigest_product_1_31_port, predigest_product_1_30_port, 
      predigest_product_1_29_port, predigest_product_1_28_port, 
      predigest_product_1_27_port, predigest_product_1_26_port, 
      predigest_product_1_25_port, predigest_product_1_24_port, 
      predigest_product_1_23_port, predigest_product_1_22_port, 
      predigest_product_1_21_port, predigest_product_1_20_port, 
      predigest_product_1_19_port, predigest_product_1_18_port, 
      predigest_product_1_17_port, predigest_product_1_16_port, 
      predigest_product_1_15_port, predigest_product_1_14_port, 
      predigest_product_1_13_port, predigest_product_1_12_port, 
      predigest_product_1_11_port, predigest_product_1_10_port, 
      predigest_product_1_9_port, predigest_product_1_8_port, 
      predigest_product_1_7_port, predigest_product_1_6_port, 
      predigest_product_1_5_port, predigest_product_1_4_port, 
      predigest_product_1_3_port, predigest_product_1_2_port, 
      predigest_product_1_1_port, predigest_product_1_0_port, 
      predigest_product_2_63_port, predigest_product_2_62_port, 
      predigest_product_2_61_port, predigest_product_2_60_port, 
      predigest_product_2_59_port, predigest_product_2_58_port, 
      predigest_product_2_57_port, predigest_product_2_56_port, 
      predigest_product_2_55_port, predigest_product_2_54_port, 
      predigest_product_2_53_port, predigest_product_2_52_port, 
      predigest_product_2_51_port, predigest_product_2_50_port, 
      predigest_product_2_49_port, predigest_product_2_48_port, 
      predigest_product_2_47_port, predigest_product_2_46_port, 
      predigest_product_2_45_port, predigest_product_2_44_port, 
      predigest_product_2_43_port, predigest_product_2_42_port, 
      predigest_product_2_41_port, predigest_product_2_40_port, 
      predigest_product_2_39_port, predigest_product_2_38_port, 
      predigest_product_2_37_port, predigest_product_2_36_port, 
      predigest_product_2_35_port, predigest_product_2_34_port, 
      predigest_product_2_33_port, predigest_product_2_32_port, 
      predigest_product_2_31_port, predigest_product_2_30_port, 
      predigest_product_2_29_port, predigest_product_2_28_port, 
      predigest_product_2_27_port, predigest_product_2_26_port, 
      predigest_product_2_25_port, predigest_product_2_24_port, 
      predigest_product_2_23_port, predigest_product_2_22_port, 
      predigest_product_2_21_port, predigest_product_2_20_port, 
      predigest_product_2_19_port, predigest_product_2_18_port, 
      predigest_product_2_17_port, predigest_product_2_16_port, 
      predigest_product_2_15_port, predigest_product_2_14_port, 
      predigest_product_2_13_port, predigest_product_2_12_port, 
      predigest_product_2_11_port, predigest_product_2_10_port, 
      predigest_product_2_9_port, predigest_product_2_8_port, 
      predigest_product_2_7_port, predigest_product_2_6_port, 
      predigest_product_2_5_port, predigest_product_2_4_port, 
      predigest_product_2_3_port, predigest_product_2_2_port, 
      predigest_product_2_1_port, predigest_product_2_0_port, 
      predigest_product_3_63_port, predigest_product_3_62_port, 
      predigest_product_3_61_port, predigest_product_3_60_port, 
      predigest_product_3_59_port, predigest_product_3_58_port, 
      predigest_product_3_57_port, predigest_product_3_56_port, 
      predigest_product_3_55_port, predigest_product_3_54_port, 
      predigest_product_3_53_port, predigest_product_3_52_port, 
      predigest_product_3_51_port, predigest_product_3_50_port, 
      predigest_product_3_49_port, predigest_product_3_48_port, 
      predigest_product_3_47_port, predigest_product_3_46_port, 
      predigest_product_3_45_port, predigest_product_3_44_port, 
      predigest_product_3_43_port, predigest_product_3_42_port, 
      predigest_product_3_41_port, predigest_product_3_40_port, 
      predigest_product_3_39_port, predigest_product_3_38_port, 
      predigest_product_3_37_port, predigest_product_3_36_port, 
      predigest_product_3_35_port, predigest_product_3_34_port, 
      predigest_product_3_33_port, predigest_product_3_32_port, 
      predigest_product_3_31_port, predigest_product_3_30_port, 
      predigest_product_3_29_port, predigest_product_3_28_port, 
      predigest_product_3_27_port, predigest_product_3_26_port, 
      predigest_product_3_25_port, predigest_product_3_24_port, 
      predigest_product_3_23_port, predigest_product_3_22_port, 
      predigest_product_3_21_port, predigest_product_3_20_port, 
      predigest_product_3_19_port, predigest_product_3_18_port, 
      predigest_product_3_17_port, predigest_product_3_16_port, 
      predigest_product_3_15_port, predigest_product_3_14_port, 
      predigest_product_3_13_port, predigest_product_3_12_port, 
      predigest_product_3_11_port, predigest_product_3_10_port, 
      predigest_product_3_9_port, predigest_product_3_8_port, 
      predigest_product_3_7_port, predigest_product_3_6_port, 
      predigest_product_3_5_port, predigest_product_3_4_port, 
      predigest_product_3_3_port, predigest_product_3_2_port, 
      predigest_product_3_1_port, predigest_product_3_0_port, 
      predigest_product_4_63_port, predigest_product_4_62_port, 
      predigest_product_4_61_port, predigest_product_4_60_port, 
      predigest_product_4_59_port, predigest_product_4_58_port, 
      predigest_product_4_57_port, predigest_product_4_56_port, 
      predigest_product_4_55_port, predigest_product_4_54_port, 
      predigest_product_4_53_port, predigest_product_4_52_port, 
      predigest_product_4_51_port, predigest_product_4_50_port, 
      predigest_product_4_49_port, predigest_product_4_48_port, 
      predigest_product_4_47_port, predigest_product_4_46_port, 
      predigest_product_4_45_port, predigest_product_4_44_port, 
      predigest_product_4_43_port, predigest_product_4_42_port, 
      predigest_product_4_41_port, predigest_product_4_40_port, 
      predigest_product_4_39_port, predigest_product_4_38_port, 
      predigest_product_4_37_port, predigest_product_4_36_port, 
      predigest_product_4_35_port, predigest_product_4_34_port, 
      predigest_product_4_33_port, predigest_product_4_32_port, 
      predigest_product_4_31_port, predigest_product_4_30_port, 
      predigest_product_4_29_port, predigest_product_4_28_port, 
      predigest_product_4_27_port, predigest_product_4_26_port, 
      predigest_product_4_25_port, predigest_product_4_24_port, 
      predigest_product_4_23_port, predigest_product_4_22_port, 
      predigest_product_4_21_port, predigest_product_4_20_port, 
      predigest_product_4_19_port, predigest_product_4_18_port, 
      predigest_product_4_17_port, predigest_product_4_16_port, 
      predigest_product_4_15_port, predigest_product_4_14_port, 
      predigest_product_4_13_port, predigest_product_4_12_port, 
      predigest_product_4_11_port, predigest_product_4_10_port, 
      predigest_product_4_9_port, predigest_product_4_8_port, 
      predigest_product_4_7_port, predigest_product_4_6_port, 
      predigest_product_4_5_port, predigest_product_4_4_port, 
      predigest_product_4_3_port, predigest_product_4_2_port, 
      predigest_product_4_1_port, predigest_product_4_0_port, 
      predigest_product_5_63_port, predigest_product_5_62_port, 
      predigest_product_5_61_port, predigest_product_5_60_port, 
      predigest_product_5_59_port, predigest_product_5_58_port, 
      predigest_product_5_57_port, predigest_product_5_56_port, 
      predigest_product_5_55_port, predigest_product_5_54_port, 
      predigest_product_5_53_port, predigest_product_5_52_port, 
      predigest_product_5_51_port, predigest_product_5_50_port, 
      predigest_product_5_49_port, predigest_product_5_48_port, 
      predigest_product_5_47_port, predigest_product_5_46_port, 
      predigest_product_5_45_port, predigest_product_5_44_port, 
      predigest_product_5_43_port, predigest_product_5_42_port, 
      predigest_product_5_41_port, predigest_product_5_40_port, 
      predigest_product_5_39_port, predigest_product_5_38_port, 
      predigest_product_5_37_port, predigest_product_5_36_port, 
      predigest_product_5_35_port, predigest_product_5_34_port, 
      predigest_product_5_33_port, predigest_product_5_32_port, 
      predigest_product_5_31_port, predigest_product_5_30_port, 
      predigest_product_5_29_port, predigest_product_5_28_port, 
      predigest_product_5_27_port, predigest_product_5_26_port, 
      predigest_product_5_25_port, predigest_product_5_24_port, 
      predigest_product_5_23_port, predigest_product_5_22_port, 
      predigest_product_5_21_port, predigest_product_5_20_port, 
      predigest_product_5_19_port, predigest_product_5_18_port, 
      predigest_product_5_17_port, predigest_product_5_16_port, 
      predigest_product_5_15_port, predigest_product_5_14_port, 
      predigest_product_5_13_port, predigest_product_5_12_port, 
      predigest_product_5_11_port, predigest_product_5_10_port, 
      predigest_product_5_9_port, predigest_product_5_8_port, 
      predigest_product_5_7_port, predigest_product_5_6_port, 
      predigest_product_5_5_port, predigest_product_5_4_port, 
      predigest_product_5_3_port, predigest_product_5_2_port, 
      predigest_product_5_1_port, predigest_product_5_0_port, 
      predigest_product_6_63_port, predigest_product_6_62_port, 
      predigest_product_6_61_port, predigest_product_6_60_port, 
      predigest_product_6_59_port, predigest_product_6_58_port, 
      predigest_product_6_57_port, predigest_product_6_56_port, 
      predigest_product_6_55_port, predigest_product_6_54_port, 
      predigest_product_6_53_port, predigest_product_6_52_port, 
      predigest_product_6_51_port, predigest_product_6_50_port, 
      predigest_product_6_49_port, predigest_product_6_48_port, 
      predigest_product_6_47_port, predigest_product_6_46_port, 
      predigest_product_6_45_port, predigest_product_6_44_port, 
      predigest_product_6_43_port, predigest_product_6_42_port, 
      predigest_product_6_41_port, predigest_product_6_40_port, 
      predigest_product_6_39_port, predigest_product_6_38_port, 
      predigest_product_6_37_port, predigest_product_6_36_port, 
      predigest_product_6_35_port, predigest_product_6_34_port, 
      predigest_product_6_33_port, predigest_product_6_32_port, 
      predigest_product_6_31_port, predigest_product_6_30_port, 
      predigest_product_6_29_port, predigest_product_6_28_port, 
      predigest_product_6_27_port, predigest_product_6_26_port, 
      predigest_product_6_25_port, predigest_product_6_24_port, 
      predigest_product_6_23_port, predigest_product_6_22_port, 
      predigest_product_6_21_port, predigest_product_6_20_port, 
      predigest_product_6_19_port, predigest_product_6_18_port, 
      predigest_product_6_17_port, predigest_product_6_16_port, 
      predigest_product_6_15_port, predigest_product_6_14_port, 
      predigest_product_6_13_port, predigest_product_6_12_port, 
      predigest_product_6_11_port, predigest_product_6_10_port, 
      predigest_product_6_9_port, predigest_product_6_8_port, 
      predigest_product_6_7_port, predigest_product_6_6_port, 
      predigest_product_6_5_port, predigest_product_6_4_port, 
      predigest_product_6_3_port, predigest_product_6_2_port, 
      predigest_product_6_1_port, predigest_product_6_0_port, 
      predigest_product_7_63_port, predigest_product_7_62_port, 
      predigest_product_7_61_port, predigest_product_7_60_port, 
      predigest_product_7_59_port, predigest_product_7_58_port, 
      predigest_product_7_57_port, predigest_product_7_56_port, 
      predigest_product_7_55_port, predigest_product_7_54_port, 
      predigest_product_7_53_port, predigest_product_7_52_port, 
      predigest_product_7_51_port, predigest_product_7_50_port, 
      predigest_product_7_49_port, predigest_product_7_48_port, 
      predigest_product_7_47_port, predigest_product_7_46_port, 
      predigest_product_7_45_port, predigest_product_7_44_port, 
      predigest_product_7_43_port, predigest_product_7_42_port, 
      predigest_product_7_41_port, predigest_product_7_40_port, 
      predigest_product_7_39_port, predigest_product_7_38_port, 
      predigest_product_7_37_port, predigest_product_7_36_port, 
      predigest_product_7_35_port, predigest_product_7_34_port, 
      predigest_product_7_33_port, predigest_product_7_32_port, 
      predigest_product_7_31_port, predigest_product_7_30_port, 
      predigest_product_7_29_port, predigest_product_7_28_port, 
      predigest_product_7_27_port, predigest_product_7_26_port, 
      predigest_product_7_25_port, predigest_product_7_24_port, 
      predigest_product_7_23_port, predigest_product_7_22_port, 
      predigest_product_7_21_port, predigest_product_7_20_port, 
      predigest_product_7_19_port, predigest_product_7_18_port, 
      predigest_product_7_17_port, predigest_product_7_16_port, 
      predigest_product_7_15_port, predigest_product_7_14_port, 
      predigest_product_7_13_port, predigest_product_7_12_port, 
      predigest_product_7_11_port, predigest_product_7_10_port, 
      predigest_product_7_9_port, predigest_product_7_8_port, 
      predigest_product_7_7_port, predigest_product_7_6_port, 
      predigest_product_7_5_port, predigest_product_7_4_port, 
      predigest_product_7_3_port, predigest_product_7_2_port, 
      predigest_product_7_1_port, predigest_product_7_0_port, 
      out_imux_8_63_port, out_imux_8_62_port, out_imux_8_61_port, 
      out_imux_8_60_port, out_imux_8_59_port, out_imux_8_58_port, 
      out_imux_8_57_port, out_imux_8_56_port, out_imux_8_55_port, 
      out_imux_8_54_port, out_imux_8_53_port, out_imux_8_52_port, 
      out_imux_8_51_port, out_imux_8_50_port, out_imux_8_49_port, 
      out_imux_8_48_port, out_imux_8_47_port, out_imux_8_46_port, 
      out_imux_8_45_port, out_imux_8_44_port, out_imux_8_43_port, 
      out_imux_8_42_port, out_imux_8_41_port, out_imux_8_40_port, 
      out_imux_8_39_port, out_imux_8_38_port, out_imux_8_37_port, 
      out_imux_8_36_port, out_imux_8_35_port, out_imux_8_34_port, 
      out_imux_8_33_port, out_imux_8_32_port, out_imux_8_31_port, 
      out_imux_8_30_port, out_imux_8_29_port, out_imux_8_28_port, 
      out_imux_8_27_port, out_imux_8_26_port, out_imux_8_25_port, 
      out_imux_8_24_port, out_imux_8_23_port, out_imux_8_22_port, 
      out_imux_8_21_port, out_imux_8_20_port, out_imux_8_19_port, 
      out_imux_8_18_port, out_imux_8_17_port, out_imux_8_16_port, 
      out_imux_8_15_port, out_imux_8_14_port, out_imux_8_13_port, 
      out_imux_8_12_port, out_imux_8_11_port, out_imux_8_10_port, 
      out_imux_8_9_port, out_imux_8_8_port, out_imux_8_7_port, 
      out_imux_8_6_port, out_imux_8_5_port, out_imux_8_4_port, 
      out_imux_8_3_port, out_imux_8_2_port, out_imux_8_1_port, 
      out_imux_8_0_port, out_imux_9_63_port, out_imux_9_62_port, 
      out_imux_9_61_port, out_imux_9_60_port, out_imux_9_59_port, 
      out_imux_9_58_port, out_imux_9_57_port, out_imux_9_56_port, 
      out_imux_9_55_port, out_imux_9_54_port, out_imux_9_53_port, 
      out_imux_9_52_port, out_imux_9_51_port, out_imux_9_50_port, 
      out_imux_9_49_port, out_imux_9_48_port, out_imux_9_47_port, 
      out_imux_9_46_port, out_imux_9_45_port, out_imux_9_44_port, 
      out_imux_9_43_port, out_imux_9_42_port, out_imux_9_41_port, 
      out_imux_9_40_port, out_imux_9_39_port, out_imux_9_38_port, 
      out_imux_9_37_port, out_imux_9_36_port, out_imux_9_35_port, 
      out_imux_9_34_port, out_imux_9_33_port, out_imux_9_32_port, 
      out_imux_9_31_port, out_imux_9_30_port, out_imux_9_29_port, 
      out_imux_9_28_port, out_imux_9_27_port, out_imux_9_26_port, 
      out_imux_9_25_port, out_imux_9_24_port, out_imux_9_23_port, 
      out_imux_9_22_port, out_imux_9_21_port, out_imux_9_20_port, 
      out_imux_9_19_port, out_imux_9_18_port, out_imux_9_17_port, 
      out_imux_9_16_port, out_imux_9_15_port, out_imux_9_14_port, 
      out_imux_9_13_port, out_imux_9_12_port, out_imux_9_11_port, 
      out_imux_9_10_port, out_imux_9_9_port, out_imux_9_8_port, 
      out_imux_9_7_port, out_imux_9_6_port, out_imux_9_5_port, 
      out_imux_9_4_port, out_imux_9_3_port, out_imux_9_2_port, 
      out_imux_9_1_port, out_imux_9_0_port, out_imux_10_63_port, 
      out_imux_10_62_port, out_imux_10_61_port, out_imux_10_60_port, 
      out_imux_10_59_port, out_imux_10_58_port, out_imux_10_57_port, 
      out_imux_10_56_port, out_imux_10_55_port, out_imux_10_54_port, 
      out_imux_10_53_port, out_imux_10_52_port, out_imux_10_51_port, 
      out_imux_10_50_port, out_imux_10_49_port, out_imux_10_48_port, 
      out_imux_10_47_port, out_imux_10_46_port, out_imux_10_45_port, 
      out_imux_10_44_port, out_imux_10_43_port, out_imux_10_42_port, 
      out_imux_10_41_port, out_imux_10_40_port, out_imux_10_39_port, 
      out_imux_10_38_port, out_imux_10_37_port, out_imux_10_36_port, 
      out_imux_10_35_port, out_imux_10_34_port, out_imux_10_33_port, 
      out_imux_10_32_port, out_imux_10_31_port, out_imux_10_30_port, 
      out_imux_10_29_port, out_imux_10_28_port, out_imux_10_27_port, 
      out_imux_10_26_port, out_imux_10_25_port, out_imux_10_24_port, 
      out_imux_10_23_port, out_imux_10_22_port, out_imux_10_21_port, 
      out_imux_10_20_port, out_imux_10_19_port, out_imux_10_18_port, 
      out_imux_10_17_port, out_imux_10_16_port, out_imux_10_15_port, 
      out_imux_10_14_port, out_imux_10_13_port, out_imux_10_12_port, 
      out_imux_10_11_port, out_imux_10_10_port, out_imux_10_9_port, 
      out_imux_10_8_port, out_imux_10_7_port, out_imux_10_6_port, 
      out_imux_10_5_port, out_imux_10_4_port, out_imux_10_3_port, 
      out_imux_10_2_port, out_imux_10_1_port, out_imux_10_0_port, 
      out_imux_11_63_port, out_imux_11_62_port, out_imux_11_61_port, 
      out_imux_11_60_port, out_imux_11_59_port, out_imux_11_58_port, 
      out_imux_11_57_port, out_imux_11_56_port, out_imux_11_55_port, 
      out_imux_11_54_port, out_imux_11_53_port, out_imux_11_52_port, 
      out_imux_11_51_port, out_imux_11_50_port, out_imux_11_49_port, 
      out_imux_11_48_port, out_imux_11_47_port, out_imux_11_46_port, 
      out_imux_11_45_port, out_imux_11_44_port, out_imux_11_43_port, 
      out_imux_11_42_port, out_imux_11_41_port, out_imux_11_40_port, 
      out_imux_11_39_port, out_imux_11_38_port, out_imux_11_37_port, 
      out_imux_11_36_port, out_imux_11_35_port, out_imux_11_34_port, 
      out_imux_11_33_port, out_imux_11_32_port, out_imux_11_31_port, 
      out_imux_11_30_port, out_imux_11_29_port, out_imux_11_28_port, 
      out_imux_11_27_port, out_imux_11_26_port, out_imux_11_25_port, 
      out_imux_11_24_port, out_imux_11_23_port, out_imux_11_22_port, 
      out_imux_11_21_port, out_imux_11_20_port, out_imux_11_19_port, 
      out_imux_11_18_port, out_imux_11_17_port, out_imux_11_16_port, 
      out_imux_11_15_port, out_imux_11_14_port, out_imux_11_13_port, 
      out_imux_11_12_port, out_imux_11_11_port, out_imux_11_10_port, 
      out_imux_11_9_port, out_imux_11_8_port, out_imux_11_7_port, 
      out_imux_11_6_port, out_imux_11_5_port, out_imux_11_4_port, 
      out_imux_11_3_port, out_imux_11_2_port, out_imux_11_1_port, 
      out_imux_11_0_port, out_imux_12_63_port, out_imux_12_62_port, 
      out_imux_12_61_port, out_imux_12_60_port, out_imux_12_59_port, 
      out_imux_12_58_port, out_imux_12_57_port, out_imux_12_56_port, 
      out_imux_12_55_port, out_imux_12_54_port, out_imux_12_53_port, 
      out_imux_12_52_port, out_imux_12_51_port, out_imux_12_50_port, 
      out_imux_12_49_port, out_imux_12_48_port, out_imux_12_47_port, 
      out_imux_12_46_port, out_imux_12_45_port, out_imux_12_44_port, 
      out_imux_12_43_port, out_imux_12_42_port, out_imux_12_41_port, 
      out_imux_12_40_port, out_imux_12_39_port, out_imux_12_38_port, 
      out_imux_12_37_port, out_imux_12_36_port, out_imux_12_35_port, 
      out_imux_12_34_port, out_imux_12_33_port, out_imux_12_32_port, 
      out_imux_12_31_port, out_imux_12_30_port, out_imux_12_29_port, 
      out_imux_12_28_port, out_imux_12_27_port, out_imux_12_26_port, 
      out_imux_12_25_port, out_imux_12_24_port, out_imux_12_23_port, 
      out_imux_12_22_port, out_imux_12_21_port, out_imux_12_20_port, 
      out_imux_12_19_port, out_imux_12_18_port, out_imux_12_17_port, 
      out_imux_12_16_port, out_imux_12_15_port, out_imux_12_14_port, 
      out_imux_12_13_port, out_imux_12_12_port, out_imux_12_11_port, 
      out_imux_12_10_port, out_imux_12_9_port, out_imux_12_8_port, 
      out_imux_12_7_port, out_imux_12_6_port, out_imux_12_5_port, 
      out_imux_12_4_port, out_imux_12_3_port, out_imux_12_2_port, 
      out_imux_12_1_port, out_imux_12_0_port, out_imux_13_63_port, 
      out_imux_13_62_port, out_imux_13_61_port, out_imux_13_60_port, 
      out_imux_13_59_port, out_imux_13_58_port, out_imux_13_57_port, 
      out_imux_13_56_port, out_imux_13_55_port, out_imux_13_54_port, 
      out_imux_13_53_port, out_imux_13_52_port, out_imux_13_51_port, 
      out_imux_13_50_port, out_imux_13_49_port, out_imux_13_48_port, 
      out_imux_13_47_port, out_imux_13_46_port, out_imux_13_45_port, 
      out_imux_13_44_port, out_imux_13_43_port, out_imux_13_42_port, 
      out_imux_13_41_port, out_imux_13_40_port, out_imux_13_39_port, 
      out_imux_13_38_port, out_imux_13_37_port, out_imux_13_36_port, 
      out_imux_13_35_port, out_imux_13_34_port, out_imux_13_33_port, 
      out_imux_13_32_port, out_imux_13_31_port, out_imux_13_30_port, 
      out_imux_13_29_port, out_imux_13_28_port, out_imux_13_27_port, 
      out_imux_13_26_port, out_imux_13_25_port, out_imux_13_24_port, 
      out_imux_13_23_port, out_imux_13_22_port, out_imux_13_21_port, 
      out_imux_13_20_port, out_imux_13_19_port, out_imux_13_18_port, 
      out_imux_13_17_port, out_imux_13_16_port, out_imux_13_15_port, 
      out_imux_13_14_port, out_imux_13_13_port, out_imux_13_12_port, 
      out_imux_13_11_port, out_imux_13_10_port, out_imux_13_9_port, 
      out_imux_13_8_port, out_imux_13_7_port, out_imux_13_6_port, 
      out_imux_13_5_port, out_imux_13_4_port, out_imux_13_3_port, 
      out_imux_13_2_port, out_imux_13_1_port, out_imux_13_0_port, 
      out_imux_14_63_port, out_imux_14_62_port, out_imux_14_61_port, 
      out_imux_14_60_port, out_imux_14_59_port, out_imux_14_58_port, 
      out_imux_14_57_port, out_imux_14_56_port, out_imux_14_55_port, 
      out_imux_14_54_port, out_imux_14_53_port, out_imux_14_52_port, 
      out_imux_14_51_port, out_imux_14_50_port, out_imux_14_49_port, 
      out_imux_14_48_port, out_imux_14_47_port, out_imux_14_46_port, 
      out_imux_14_45_port, out_imux_14_44_port, out_imux_14_43_port, 
      out_imux_14_42_port, out_imux_14_41_port, out_imux_14_40_port, 
      out_imux_14_39_port, out_imux_14_38_port, out_imux_14_37_port, 
      out_imux_14_36_port, out_imux_14_35_port, out_imux_14_34_port, 
      out_imux_14_33_port, out_imux_14_32_port, out_imux_14_31_port, 
      out_imux_14_30_port, out_imux_14_29_port, out_imux_14_28_port, 
      out_imux_14_27_port, out_imux_14_26_port, out_imux_14_25_port, 
      out_imux_14_24_port, out_imux_14_23_port, out_imux_14_22_port, 
      out_imux_14_21_port, out_imux_14_20_port, out_imux_14_19_port, 
      out_imux_14_18_port, out_imux_14_17_port, out_imux_14_16_port, 
      out_imux_14_15_port, out_imux_14_14_port, out_imux_14_13_port, 
      out_imux_14_12_port, out_imux_14_11_port, out_imux_14_10_port, 
      out_imux_14_9_port, out_imux_14_8_port, out_imux_14_7_port, 
      out_imux_14_6_port, out_imux_14_5_port, out_imux_14_4_port, 
      out_imux_14_3_port, out_imux_14_2_port, out_imux_14_1_port, 
      out_imux_14_0_port, out_imux_15_63_port, out_imux_15_62_port, 
      out_imux_15_61_port, out_imux_15_60_port, out_imux_15_59_port, 
      out_imux_15_58_port, out_imux_15_57_port, out_imux_15_56_port, 
      out_imux_15_55_port, out_imux_15_54_port, out_imux_15_53_port, 
      out_imux_15_52_port, out_imux_15_51_port, out_imux_15_50_port, 
      out_imux_15_49_port, out_imux_15_48_port, out_imux_15_47_port, 
      out_imux_15_46_port, out_imux_15_45_port, out_imux_15_44_port, 
      out_imux_15_43_port, out_imux_15_42_port, out_imux_15_41_port, 
      out_imux_15_40_port, out_imux_15_39_port, out_imux_15_38_port, 
      out_imux_15_37_port, out_imux_15_36_port, out_imux_15_35_port, 
      out_imux_15_34_port, out_imux_15_33_port, out_imux_15_32_port, 
      out_imux_15_31_port, out_imux_15_30_port, out_imux_15_29_port, 
      out_imux_15_28_port, out_imux_15_27_port, out_imux_15_26_port, 
      out_imux_15_25_port, out_imux_15_24_port, out_imux_15_23_port, 
      out_imux_15_22_port, out_imux_15_21_port, out_imux_15_20_port, 
      out_imux_15_19_port, out_imux_15_18_port, out_imux_15_17_port, 
      out_imux_15_16_port, out_imux_15_15_port, out_imux_15_14_port, 
      out_imux_15_13_port, out_imux_15_12_port, out_imux_15_11_port, 
      out_imux_15_10_port, out_imux_15_9_port, out_imux_15_8_port, 
      out_imux_15_7_port, out_imux_15_6_port, out_imux_15_5_port, 
      out_imux_15_4_port, out_imux_15_3_port, out_imux_15_2_port, 
      out_imux_15_1_port, out_imux_15_0_port, predigest_product_8_63_port, 
      predigest_product_8_62_port, predigest_product_8_61_port, 
      predigest_product_8_60_port, predigest_product_8_59_port, 
      predigest_product_8_58_port, predigest_product_8_57_port, 
      predigest_product_8_56_port, predigest_product_8_55_port, 
      predigest_product_8_54_port, predigest_product_8_53_port, 
      predigest_product_8_52_port, predigest_product_8_51_port, 
      predigest_product_8_50_port, predigest_product_8_49_port, 
      predigest_product_8_48_port, predigest_product_8_47_port, 
      predigest_product_8_46_port, predigest_product_8_45_port, 
      predigest_product_8_44_port, predigest_product_8_43_port, 
      predigest_product_8_42_port, predigest_product_8_41_port, 
      predigest_product_8_40_port, predigest_product_8_39_port, 
      predigest_product_8_38_port, predigest_product_8_37_port, 
      predigest_product_8_36_port, predigest_product_8_35_port, 
      predigest_product_8_34_port, predigest_product_8_33_port, 
      predigest_product_8_32_port, predigest_product_8_31_port, 
      predigest_product_8_30_port, predigest_product_8_29_port, 
      predigest_product_8_28_port, predigest_product_8_27_port, 
      predigest_product_8_26_port, predigest_product_8_25_port, 
      predigest_product_8_24_port, predigest_product_8_23_port, 
      predigest_product_8_22_port, predigest_product_8_21_port, 
      predigest_product_8_20_port, predigest_product_8_19_port, 
      predigest_product_8_18_port, predigest_product_8_17_port, 
      predigest_product_8_16_port, predigest_product_8_15_port, 
      predigest_product_8_14_port, predigest_product_8_13_port, 
      predigest_product_8_12_port, predigest_product_8_11_port, 
      predigest_product_8_10_port, predigest_product_8_9_port, 
      predigest_product_8_8_port, predigest_product_8_7_port, 
      predigest_product_8_6_port, predigest_product_8_5_port, 
      predigest_product_8_4_port, predigest_product_8_3_port, 
      predigest_product_8_2_port, predigest_product_8_1_port, 
      predigest_product_8_0_port, predigest_product_9_63_port, 
      predigest_product_9_62_port, predigest_product_9_61_port, 
      predigest_product_9_60_port, predigest_product_9_59_port, 
      predigest_product_9_58_port, predigest_product_9_57_port, 
      predigest_product_9_56_port, predigest_product_9_55_port, 
      predigest_product_9_54_port, predigest_product_9_53_port, 
      predigest_product_9_52_port, predigest_product_9_51_port, 
      predigest_product_9_50_port, predigest_product_9_49_port, 
      predigest_product_9_48_port, predigest_product_9_47_port, 
      predigest_product_9_46_port, predigest_product_9_45_port, 
      predigest_product_9_44_port, predigest_product_9_43_port, 
      predigest_product_9_42_port, predigest_product_9_41_port, 
      predigest_product_9_40_port, predigest_product_9_39_port, 
      predigest_product_9_38_port, predigest_product_9_37_port, 
      predigest_product_9_36_port, predigest_product_9_35_port, 
      predigest_product_9_34_port, predigest_product_9_33_port, 
      predigest_product_9_32_port, predigest_product_9_31_port, 
      predigest_product_9_30_port, predigest_product_9_29_port, 
      predigest_product_9_28_port, predigest_product_9_27_port, 
      predigest_product_9_26_port, predigest_product_9_25_port, 
      predigest_product_9_24_port, predigest_product_9_23_port, 
      predigest_product_9_22_port, predigest_product_9_21_port, 
      predigest_product_9_20_port, predigest_product_9_19_port, 
      predigest_product_9_18_port, predigest_product_9_17_port, 
      predigest_product_9_16_port, predigest_product_9_15_port, 
      predigest_product_9_14_port, predigest_product_9_13_port, 
      predigest_product_9_12_port, predigest_product_9_11_port, 
      predigest_product_9_10_port, predigest_product_9_9_port, 
      predigest_product_9_8_port, predigest_product_9_7_port, 
      predigest_product_9_6_port, predigest_product_9_5_port, 
      predigest_product_9_4_port, predigest_product_9_3_port, 
      predigest_product_9_2_port, predigest_product_9_1_port, 
      predigest_product_9_0_port, predigest_product_10_63_port, 
      predigest_product_10_62_port, predigest_product_10_61_port, 
      predigest_product_10_60_port, predigest_product_10_59_port, 
      predigest_product_10_58_port, predigest_product_10_57_port, 
      predigest_product_10_56_port, predigest_product_10_55_port, 
      predigest_product_10_54_port, predigest_product_10_53_port, 
      predigest_product_10_52_port, predigest_product_10_51_port, 
      predigest_product_10_50_port, predigest_product_10_49_port, 
      predigest_product_10_48_port, predigest_product_10_47_port, 
      predigest_product_10_46_port, predigest_product_10_45_port, 
      predigest_product_10_44_port, predigest_product_10_43_port, 
      predigest_product_10_42_port, predigest_product_10_41_port, 
      predigest_product_10_40_port, predigest_product_10_39_port, 
      predigest_product_10_38_port, predigest_product_10_37_port, 
      predigest_product_10_36_port, predigest_product_10_35_port, 
      predigest_product_10_34_port, predigest_product_10_33_port, 
      predigest_product_10_32_port, predigest_product_10_31_port, 
      predigest_product_10_30_port, predigest_product_10_29_port, 
      predigest_product_10_28_port, predigest_product_10_27_port, 
      predigest_product_10_26_port, predigest_product_10_25_port, 
      predigest_product_10_24_port, predigest_product_10_23_port, 
      predigest_product_10_22_port, predigest_product_10_21_port, 
      predigest_product_10_20_port, predigest_product_10_19_port, 
      predigest_product_10_18_port, predigest_product_10_17_port, 
      predigest_product_10_16_port, predigest_product_10_15_port, 
      predigest_product_10_14_port, predigest_product_10_13_port, 
      predigest_product_10_12_port, predigest_product_10_11_port, 
      predigest_product_10_10_port, predigest_product_10_9_port, 
      predigest_product_10_8_port, predigest_product_10_7_port, 
      predigest_product_10_6_port, predigest_product_10_5_port, 
      predigest_product_10_4_port, predigest_product_10_3_port, 
      predigest_product_10_2_port, predigest_product_10_1_port, 
      predigest_product_10_0_port, predigest_product_11_63_port, 
      predigest_product_11_62_port, predigest_product_11_61_port, 
      predigest_product_11_60_port, predigest_product_11_59_port, 
      predigest_product_11_58_port, predigest_product_11_57_port, 
      predigest_product_11_56_port, predigest_product_11_55_port, 
      predigest_product_11_54_port, predigest_product_11_53_port, 
      predigest_product_11_52_port, predigest_product_11_51_port, 
      predigest_product_11_50_port, predigest_product_11_49_port, 
      predigest_product_11_48_port, predigest_product_11_47_port, 
      predigest_product_11_46_port, predigest_product_11_45_port, 
      predigest_product_11_44_port, predigest_product_11_43_port, 
      predigest_product_11_42_port, predigest_product_11_41_port, 
      predigest_product_11_40_port, predigest_product_11_39_port, 
      predigest_product_11_38_port, predigest_product_11_37_port, 
      predigest_product_11_36_port, predigest_product_11_35_port, 
      predigest_product_11_34_port, predigest_product_11_33_port, 
      predigest_product_11_32_port, predigest_product_11_31_port, 
      predigest_product_11_30_port, predigest_product_11_29_port, 
      predigest_product_11_28_port, predigest_product_11_27_port, 
      predigest_product_11_26_port, predigest_product_11_25_port, 
      predigest_product_11_24_port, predigest_product_11_23_port, 
      predigest_product_11_22_port, predigest_product_11_21_port, 
      predigest_product_11_20_port, predigest_product_11_19_port, 
      predigest_product_11_18_port, predigest_product_11_17_port, 
      predigest_product_11_16_port, predigest_product_11_15_port, 
      predigest_product_11_14_port, predigest_product_11_13_port, 
      predigest_product_11_12_port, predigest_product_11_11_port, 
      predigest_product_11_10_port, predigest_product_11_9_port, 
      predigest_product_11_8_port, predigest_product_11_7_port, 
      predigest_product_11_6_port, predigest_product_11_5_port, 
      predigest_product_11_4_port, predigest_product_11_3_port, 
      predigest_product_11_2_port, predigest_product_11_1_port, 
      predigest_product_11_0_port, predigest_product_12_63_port, 
      predigest_product_12_62_port, predigest_product_12_61_port, 
      predigest_product_12_60_port, predigest_product_12_59_port, 
      predigest_product_12_58_port, predigest_product_12_57_port, 
      predigest_product_12_56_port, predigest_product_12_55_port, 
      predigest_product_12_54_port, predigest_product_12_53_port, 
      predigest_product_12_52_port, predigest_product_12_51_port, 
      predigest_product_12_50_port, predigest_product_12_49_port, 
      predigest_product_12_48_port, predigest_product_12_47_port, 
      predigest_product_12_46_port, predigest_product_12_45_port, 
      predigest_product_12_44_port, predigest_product_12_43_port, 
      predigest_product_12_42_port, predigest_product_12_41_port, 
      predigest_product_12_40_port, predigest_product_12_39_port, 
      predigest_product_12_38_port, predigest_product_12_37_port, 
      predigest_product_12_36_port, predigest_product_12_35_port, 
      predigest_product_12_34_port, predigest_product_12_33_port, 
      predigest_product_12_32_port, predigest_product_12_31_port, 
      predigest_product_12_30_port, predigest_product_12_29_port, 
      predigest_product_12_28_port, predigest_product_12_27_port, 
      predigest_product_12_26_port, predigest_product_12_25_port, 
      predigest_product_12_24_port, predigest_product_12_23_port, 
      predigest_product_12_22_port, predigest_product_12_21_port, 
      predigest_product_12_20_port, predigest_product_12_19_port, 
      predigest_product_12_18_port, predigest_product_12_17_port, 
      predigest_product_12_16_port, predigest_product_12_15_port, 
      predigest_product_12_14_port, predigest_product_12_13_port, 
      predigest_product_12_12_port, predigest_product_12_11_port, 
      predigest_product_12_10_port, predigest_product_12_9_port, 
      predigest_product_12_8_port, predigest_product_12_7_port, 
      predigest_product_12_6_port, predigest_product_12_5_port, 
      predigest_product_12_4_port, predigest_product_12_3_port, 
      predigest_product_12_2_port, predigest_product_12_1_port, 
      predigest_product_12_0_port, predigest_product_13_63_port, 
      predigest_product_13_62_port, predigest_product_13_61_port, 
      predigest_product_13_60_port, predigest_product_13_59_port, 
      predigest_product_13_58_port, predigest_product_13_57_port, 
      predigest_product_13_56_port, predigest_product_13_55_port, 
      predigest_product_13_54_port, predigest_product_13_53_port, 
      predigest_product_13_52_port, predigest_product_13_51_port, 
      predigest_product_13_50_port, predigest_product_13_49_port, 
      predigest_product_13_48_port, predigest_product_13_47_port, 
      predigest_product_13_46_port, predigest_product_13_45_port, 
      predigest_product_13_44_port, predigest_product_13_43_port, 
      predigest_product_13_42_port, predigest_product_13_41_port, 
      predigest_product_13_40_port, predigest_product_13_39_port, 
      predigest_product_13_38_port, predigest_product_13_37_port, 
      predigest_product_13_36_port, predigest_product_13_35_port, 
      predigest_product_13_34_port, predigest_product_13_33_port, 
      predigest_product_13_32_port, predigest_product_13_31_port, 
      predigest_product_13_30_port, predigest_product_13_29_port, 
      predigest_product_13_28_port, predigest_product_13_27_port, 
      predigest_product_13_26_port, predigest_product_13_25_port, 
      predigest_product_13_24_port, predigest_product_13_23_port, 
      predigest_product_13_22_port, predigest_product_13_21_port, 
      predigest_product_13_20_port, predigest_product_13_19_port, 
      predigest_product_13_18_port, predigest_product_13_17_port, 
      predigest_product_13_16_port, predigest_product_13_15_port, 
      predigest_product_13_14_port, predigest_product_13_13_port, 
      predigest_product_13_12_port, predigest_product_13_11_port, 
      predigest_product_13_10_port, predigest_product_13_9_port, 
      predigest_product_13_8_port, predigest_product_13_7_port, 
      predigest_product_13_6_port, predigest_product_13_5_port, 
      predigest_product_13_4_port, predigest_product_13_3_port, 
      predigest_product_13_2_port, predigest_product_13_1_port, 
      predigest_product_13_0_port, predigest_product_14_63_port, 
      predigest_product_14_62_port, predigest_product_14_61_port, 
      predigest_product_14_60_port, predigest_product_14_59_port, 
      predigest_product_14_58_port, predigest_product_14_57_port, 
      predigest_product_14_56_port, predigest_product_14_55_port, 
      predigest_product_14_54_port, predigest_product_14_53_port, 
      predigest_product_14_52_port, predigest_product_14_51_port, 
      predigest_product_14_50_port, predigest_product_14_49_port, 
      predigest_product_14_48_port, predigest_product_14_47_port, 
      predigest_product_14_46_port, predigest_product_14_45_port, 
      predigest_product_14_44_port, predigest_product_14_43_port, 
      predigest_product_14_42_port, predigest_product_14_41_port, 
      predigest_product_14_40_port, predigest_product_14_39_port, 
      predigest_product_14_38_port, predigest_product_14_37_port, 
      predigest_product_14_36_port, predigest_product_14_35_port, 
      predigest_product_14_34_port, predigest_product_14_33_port, 
      predigest_product_14_32_port, predigest_product_14_31_port, 
      predigest_product_14_30_port, predigest_product_14_29_port, 
      predigest_product_14_28_port, predigest_product_14_27_port, 
      predigest_product_14_26_port, predigest_product_14_25_port, 
      predigest_product_14_24_port, predigest_product_14_23_port, 
      predigest_product_14_22_port, predigest_product_14_21_port, 
      predigest_product_14_20_port, predigest_product_14_19_port, 
      predigest_product_14_18_port, predigest_product_14_17_port, 
      predigest_product_14_16_port, predigest_product_14_15_port, 
      predigest_product_14_14_port, predigest_product_14_13_port, 
      predigest_product_14_12_port, predigest_product_14_11_port, 
      predigest_product_14_10_port, predigest_product_14_9_port, 
      predigest_product_14_8_port, predigest_product_14_7_port, 
      predigest_product_14_6_port, predigest_product_14_5_port, 
      predigest_product_14_4_port, predigest_product_14_3_port, 
      predigest_product_14_2_port, predigest_product_14_1_port, 
      predigest_product_14_0_port, n33, n34, n35, n36, n37, n38, n39, n40, n41,
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106 : std_logic;

begin
   
   X_Logic0_port <= '0';
   ENC_0_0 : BOOTH_ENCODER_3BIT_4 port map( B(2) => B(1), B(1) => B(0), B(0) =>
                           X_Logic0_port, ENCODED(2) => 
                           muxs_encoded_signals_0_2_port, ENCODED(1) => 
                           muxs_encoded_signals_0_1_port, ENCODED(0) => 
                           muxs_encoded_signals_0_0_port);
   MUX_00_0 : MUX51_GENERIC_NBIT64_0 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(31), IN1(51) 
                           => A(31), IN1(50) => A(31), IN1(49) => A(31), 
                           IN1(48) => A(31), IN1(47) => A(31), IN1(46) => A(31)
                           , IN1(45) => A(31), IN1(44) => A(31), IN1(43) => 
                           A(31), IN1(42) => A(31), IN1(41) => A(31), IN1(40) 
                           => A(31), IN1(39) => A(31), IN1(38) => A(31), 
                           IN1(37) => A(31), IN1(36) => A(31), IN1(35) => A(31)
                           , IN1(34) => A(31), IN1(33) => A(31), IN1(32) => 
                           A(31), IN1(31) => A(31), IN1(30) => A(30), IN1(29) 
                           => A(29), IN1(28) => A(28), IN1(27) => A(27), 
                           IN1(26) => A(26), IN1(25) => A(25), IN1(24) => A(24)
                           , IN1(23) => A(23), IN1(22) => A(22), IN1(21) => 
                           A(21), IN1(20) => A(20), IN1(19) => A(19), IN1(18) 
                           => A(18), IN1(17) => A(17), IN1(16) => A(16), 
                           IN1(15) => A(15), IN1(14) => A(14), IN1(13) => A(13)
                           , IN1(12) => A(12), IN1(11) => A(11), IN1(10) => 
                           A(10), IN1(9) => A(9), IN1(8) => A(8), IN1(7) => 
                           A(7), IN1(6) => A(6), IN1(5) => A(5), IN1(4) => A(4)
                           , IN1(3) => A(3), IN1(2) => A(2), IN1(1) => A(1), 
                           IN1(0) => A(0), IN2(63) => negative_a_63_port, 
                           IN2(62) => negative_a_62_port, IN2(61) => 
                           negative_a_61_port, IN2(60) => negative_a_60_port, 
                           IN2(59) => negative_a_59_port, IN2(58) => 
                           negative_a_58_port, IN2(57) => negative_a_57_port, 
                           IN2(56) => negative_a_56_port, IN2(55) => 
                           negative_a_55_port, IN2(54) => negative_a_54_port, 
                           IN2(53) => negative_a_53_port, IN2(52) => 
                           negative_a_52_port, IN2(51) => negative_a_51_port, 
                           IN2(50) => negative_a_50_port, IN2(49) => 
                           negative_a_49_port, IN2(48) => negative_a_48_port, 
                           IN2(47) => negative_a_47_port, IN2(46) => 
                           negative_a_46_port, IN2(45) => negative_a_45_port, 
                           IN2(44) => negative_a_44_port, IN2(43) => 
                           negative_a_43_port, IN2(42) => negative_a_42_port, 
                           IN2(41) => negative_a_41_port, IN2(40) => 
                           negative_a_40_port, IN2(39) => negative_a_39_port, 
                           IN2(38) => negative_a_38_port, IN2(37) => 
                           negative_a_37_port, IN2(36) => negative_a_36_port, 
                           IN2(35) => negative_a_35_port, IN2(34) => 
                           negative_a_34_port, IN2(33) => n38, IN2(32) => n35, 
                           IN2(31) => negative_a_31_port, IN2(30) => 
                           negative_a_30_port, IN2(29) => negative_a_29_port, 
                           IN2(28) => negative_a_28_port, IN2(27) => 
                           negative_a_27_port, IN2(26) => negative_a_26_port, 
                           IN2(25) => negative_a_25_port, IN2(24) => 
                           negative_a_24_port, IN2(23) => negative_a_23_port, 
                           IN2(22) => negative_a_22_port, IN2(21) => 
                           negative_a_21_port, IN2(20) => negative_a_20_port, 
                           IN2(19) => negative_a_19_port, IN2(18) => 
                           negative_a_18_port, IN2(17) => negative_a_17_port, 
                           IN2(16) => negative_a_16_port, IN2(15) => 
                           negative_a_15_port, IN2(14) => negative_a_14_port, 
                           IN2(13) => negative_a_13_port, IN2(12) => 
                           negative_a_12_port, IN2(11) => negative_a_11_port, 
                           IN2(10) => negative_a_10_port, IN2(9) => 
                           negative_a_9_port, IN2(8) => negative_a_8_port, 
                           IN2(7) => negative_a_7_port, IN2(6) => 
                           negative_a_6_port, IN2(5) => negative_a_5_port, 
                           IN2(4) => negative_a_4_port, IN2(3) => 
                           negative_a_3_port, IN2(2) => negative_a_2_port, 
                           IN2(1) => negative_a_1_port, IN2(0) => 
                           negative_a_0_port, IN3(63) => A(31), IN3(62) => 
                           A(31), IN3(61) => A(31), IN3(60) => A(31), IN3(59) 
                           => A(31), IN3(58) => A(31), IN3(57) => A(31), 
                           IN3(56) => A(31), IN3(55) => A(31), IN3(54) => A(31)
                           , IN3(53) => A(31), IN3(52) => A(31), IN3(51) => 
                           A(31), IN3(50) => A(31), IN3(49) => A(31), IN3(48) 
                           => A(31), IN3(47) => A(31), IN3(46) => A(31), 
                           IN3(45) => A(31), IN3(44) => A(31), IN3(43) => A(31)
                           , IN3(42) => A(31), IN3(41) => A(31), IN3(40) => 
                           A(31), IN3(39) => A(31), IN3(38) => A(31), IN3(37) 
                           => A(31), IN3(36) => A(31), IN3(35) => A(31), 
                           IN3(34) => A(31), IN3(33) => A(31), IN3(32) => A(31)
                           , IN3(31) => A(30), IN3(30) => A(29), IN3(29) => 
                           A(28), IN3(28) => A(27), IN3(27) => A(26), IN3(26) 
                           => A(25), IN3(25) => A(24), IN3(24) => A(23), 
                           IN3(23) => A(22), IN3(22) => A(21), IN3(21) => A(20)
                           , IN3(20) => A(19), IN3(19) => A(18), IN3(18) => 
                           A(17), IN3(17) => A(16), IN3(16) => A(15), IN3(15) 
                           => A(14), IN3(14) => A(13), IN3(13) => A(12), 
                           IN3(12) => A(11), IN3(11) => A(10), IN3(10) => A(9),
                           IN3(9) => A(8), IN3(8) => A(7), IN3(7) => A(6), 
                           IN3(6) => A(5), IN3(5) => A(4), IN3(4) => A(3), 
                           IN3(3) => A(2), IN3(2) => A(1), IN3(1) => A(0), 
                           IN3(0) => X_Logic0_port, IN4(63) => 
                           negative_a_62_port, IN4(62) => negative_a_61_port, 
                           IN4(61) => negative_a_60_port, IN4(60) => 
                           negative_a_59_port, IN4(59) => negative_a_58_port, 
                           IN4(58) => negative_a_57_port, IN4(57) => 
                           negative_a_56_port, IN4(56) => negative_a_55_port, 
                           IN4(55) => negative_a_54_port, IN4(54) => 
                           negative_a_53_port, IN4(53) => negative_a_52_port, 
                           IN4(52) => negative_a_51_port, IN4(51) => 
                           negative_a_50_port, IN4(50) => negative_a_49_port, 
                           IN4(49) => negative_a_48_port, IN4(48) => 
                           negative_a_47_port, IN4(47) => negative_a_46_port, 
                           IN4(46) => negative_a_45_port, IN4(45) => 
                           negative_a_44_port, IN4(44) => negative_a_43_port, 
                           IN4(43) => negative_a_42_port, IN4(42) => 
                           negative_a_41_port, IN4(41) => negative_a_40_port, 
                           IN4(40) => negative_a_39_port, IN4(39) => 
                           negative_a_38_port, IN4(38) => negative_a_37_port, 
                           IN4(37) => negative_a_36_port, IN4(36) => 
                           negative_a_35_port, IN4(35) => negative_a_34_port, 
                           IN4(34) => n38, IN4(33) => n35, IN4(32) => 
                           negative_a_31_port, IN4(31) => negative_a_30_port, 
                           IN4(30) => negative_a_29_port, IN4(29) => 
                           negative_a_28_port, IN4(28) => negative_a_27_port, 
                           IN4(27) => negative_a_26_port, IN4(26) => 
                           negative_a_25_port, IN4(25) => negative_a_24_port, 
                           IN4(24) => negative_a_23_port, IN4(23) => 
                           negative_a_22_port, IN4(22) => negative_a_21_port, 
                           IN4(21) => negative_a_20_port, IN4(20) => 
                           negative_a_19_port, IN4(19) => negative_a_18_port, 
                           IN4(18) => negative_a_17_port, IN4(17) => 
                           negative_a_16_port, IN4(16) => negative_a_15_port, 
                           IN4(15) => negative_a_14_port, IN4(14) => 
                           negative_a_13_port, IN4(13) => negative_a_12_port, 
                           IN4(12) => negative_a_11_port, IN4(11) => 
                           negative_a_10_port, IN4(10) => negative_a_9_port, 
                           IN4(9) => negative_a_8_port, IN4(8) => 
                           negative_a_7_port, IN4(7) => negative_a_6_port, 
                           IN4(6) => negative_a_5_port, IN4(5) => 
                           negative_a_4_port, IN4(4) => negative_a_3_port, 
                           IN4(3) => negative_a_2_port, IN4(2) => 
                           negative_a_1_port, IN4(1) => negative_a_0_port, 
                           IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_0_2_port, S(1) => 
                           muxs_encoded_signals_0_1_port, S(0) => 
                           muxs_encoded_signals_0_0_port, O(63) => 
                           out_imux_0_63_port, O(62) => out_imux_0_62_port, 
                           O(61) => out_imux_0_61_port, O(60) => 
                           out_imux_0_60_port, O(59) => out_imux_0_59_port, 
                           O(58) => out_imux_0_58_port, O(57) => 
                           out_imux_0_57_port, O(56) => out_imux_0_56_port, 
                           O(55) => out_imux_0_55_port, O(54) => 
                           out_imux_0_54_port, O(53) => out_imux_0_53_port, 
                           O(52) => out_imux_0_52_port, O(51) => 
                           out_imux_0_51_port, O(50) => out_imux_0_50_port, 
                           O(49) => out_imux_0_49_port, O(48) => 
                           out_imux_0_48_port, O(47) => out_imux_0_47_port, 
                           O(46) => out_imux_0_46_port, O(45) => 
                           out_imux_0_45_port, O(44) => out_imux_0_44_port, 
                           O(43) => out_imux_0_43_port, O(42) => 
                           out_imux_0_42_port, O(41) => out_imux_0_41_port, 
                           O(40) => out_imux_0_40_port, O(39) => 
                           out_imux_0_39_port, O(38) => out_imux_0_38_port, 
                           O(37) => out_imux_0_37_port, O(36) => 
                           out_imux_0_36_port, O(35) => out_imux_0_35_port, 
                           O(34) => out_imux_0_34_port, O(33) => 
                           out_imux_0_33_port, O(32) => out_imux_0_32_port, 
                           O(31) => out_imux_0_31_port, O(30) => 
                           out_imux_0_30_port, O(29) => out_imux_0_29_port, 
                           O(28) => out_imux_0_28_port, O(27) => 
                           out_imux_0_27_port, O(26) => out_imux_0_26_port, 
                           O(25) => out_imux_0_25_port, O(24) => 
                           out_imux_0_24_port, O(23) => out_imux_0_23_port, 
                           O(22) => out_imux_0_22_port, O(21) => 
                           out_imux_0_21_port, O(20) => out_imux_0_20_port, 
                           O(19) => out_imux_0_19_port, O(18) => 
                           out_imux_0_18_port, O(17) => out_imux_0_17_port, 
                           O(16) => out_imux_0_16_port, O(15) => 
                           out_imux_0_15_port, O(14) => out_imux_0_14_port, 
                           O(13) => out_imux_0_13_port, O(12) => 
                           out_imux_0_12_port, O(11) => out_imux_0_11_port, 
                           O(10) => out_imux_0_10_port, O(9) => 
                           out_imux_0_9_port, O(8) => out_imux_0_8_port, O(7) 
                           => out_imux_0_7_port, O(6) => out_imux_0_6_port, 
                           O(5) => out_imux_0_5_port, O(4) => out_imux_0_4_port
                           , O(3) => out_imux_0_3_port, O(2) => 
                           out_imux_0_2_port, O(1) => out_imux_0_1_port, O(0) 
                           => out_imux_0_0_port);
   ENC_i_1 : BOOTH_ENCODER_3BIT_19 port map( B(2) => B(3), B(1) => B(2), B(0) 
                           => B(1), ENCODED(2) => muxs_encoded_signals_1_2_port
                           , ENCODED(1) => muxs_encoded_signals_1_1_port, 
                           ENCODED(0) => muxs_encoded_signals_1_0_port);
   MUX_i_1 : MUX51_GENERIC_NBIT64_15 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(31), IN1(51) 
                           => A(31), IN1(50) => A(31), IN1(49) => A(31), 
                           IN1(48) => A(31), IN1(47) => A(31), IN1(46) => A(31)
                           , IN1(45) => A(31), IN1(44) => A(31), IN1(43) => 
                           A(31), IN1(42) => A(31), IN1(41) => A(31), IN1(40) 
                           => A(31), IN1(39) => A(31), IN1(38) => A(31), 
                           IN1(37) => A(31), IN1(36) => A(31), IN1(35) => A(31)
                           , IN1(34) => A(31), IN1(33) => A(31), IN1(32) => 
                           A(30), IN1(31) => A(29), IN1(30) => A(28), IN1(29) 
                           => A(27), IN1(28) => A(26), IN1(27) => A(25), 
                           IN1(26) => A(24), IN1(25) => A(23), IN1(24) => A(22)
                           , IN1(23) => A(21), IN1(22) => A(20), IN1(21) => 
                           A(19), IN1(20) => A(18), IN1(19) => A(17), IN1(18) 
                           => A(16), IN1(17) => A(15), IN1(16) => A(14), 
                           IN1(15) => A(13), IN1(14) => A(12), IN1(13) => A(11)
                           , IN1(12) => A(10), IN1(11) => A(9), IN1(10) => A(8)
                           , IN1(9) => A(7), IN1(8) => A(6), IN1(7) => A(5), 
                           IN1(6) => A(4), IN1(5) => A(3), IN1(4) => A(2), 
                           IN1(3) => A(1), IN1(2) => A(0), IN1(1) => 
                           X_Logic0_port, IN1(0) => X_Logic0_port, IN2(63) => 
                           negative_a_61_port, IN2(62) => negative_a_60_port, 
                           IN2(61) => negative_a_59_port, IN2(60) => 
                           negative_a_58_port, IN2(59) => negative_a_57_port, 
                           IN2(58) => negative_a_56_port, IN2(57) => 
                           negative_a_55_port, IN2(56) => negative_a_54_port, 
                           IN2(55) => negative_a_53_port, IN2(54) => 
                           negative_a_52_port, IN2(53) => negative_a_51_port, 
                           IN2(52) => negative_a_50_port, IN2(51) => 
                           negative_a_49_port, IN2(50) => negative_a_48_port, 
                           IN2(49) => negative_a_47_port, IN2(48) => 
                           negative_a_46_port, IN2(47) => negative_a_45_port, 
                           IN2(46) => negative_a_44_port, IN2(45) => 
                           negative_a_43_port, IN2(44) => negative_a_42_port, 
                           IN2(43) => negative_a_41_port, IN2(42) => 
                           negative_a_40_port, IN2(41) => negative_a_39_port, 
                           IN2(40) => negative_a_38_port, IN2(39) => 
                           negative_a_37_port, IN2(38) => negative_a_36_port, 
                           IN2(37) => negative_a_35_port, IN2(36) => 
                           negative_a_34_port, IN2(35) => n36, IN2(34) => n33, 
                           IN2(33) => negative_a_31_port, IN2(32) => 
                           negative_a_30_port, IN2(31) => negative_a_29_port, 
                           IN2(30) => negative_a_28_port, IN2(29) => 
                           negative_a_27_port, IN2(28) => negative_a_26_port, 
                           IN2(27) => negative_a_25_port, IN2(26) => 
                           negative_a_24_port, IN2(25) => negative_a_23_port, 
                           IN2(24) => negative_a_22_port, IN2(23) => 
                           negative_a_21_port, IN2(22) => negative_a_20_port, 
                           IN2(21) => negative_a_19_port, IN2(20) => 
                           negative_a_18_port, IN2(19) => negative_a_17_port, 
                           IN2(18) => negative_a_16_port, IN2(17) => 
                           negative_a_15_port, IN2(16) => negative_a_14_port, 
                           IN2(15) => negative_a_13_port, IN2(14) => 
                           negative_a_12_port, IN2(13) => negative_a_11_port, 
                           IN2(12) => negative_a_10_port, IN2(11) => 
                           negative_a_9_port, IN2(10) => negative_a_8_port, 
                           IN2(9) => negative_a_7_port, IN2(8) => 
                           negative_a_6_port, IN2(7) => negative_a_5_port, 
                           IN2(6) => negative_a_4_port, IN2(5) => 
                           negative_a_3_port, IN2(4) => negative_a_2_port, 
                           IN2(3) => negative_a_1_port, IN2(2) => 
                           negative_a_0_port, IN2(1) => X_Logic0_port, IN2(0) 
                           => X_Logic0_port, IN3(63) => A(31), IN3(62) => A(31)
                           , IN3(61) => A(31), IN3(60) => A(31), IN3(59) => 
                           A(31), IN3(58) => A(31), IN3(57) => A(31), IN3(56) 
                           => A(31), IN3(55) => A(31), IN3(54) => A(31), 
                           IN3(53) => A(31), IN3(52) => A(31), IN3(51) => A(31)
                           , IN3(50) => A(31), IN3(49) => A(31), IN3(48) => 
                           A(31), IN3(47) => A(31), IN3(46) => A(31), IN3(45) 
                           => A(31), IN3(44) => A(31), IN3(43) => A(31), 
                           IN3(42) => A(31), IN3(41) => A(31), IN3(40) => A(31)
                           , IN3(39) => A(31), IN3(38) => A(31), IN3(37) => 
                           A(31), IN3(36) => A(31), IN3(35) => A(31), IN3(34) 
                           => A(31), IN3(33) => A(30), IN3(32) => A(29), 
                           IN3(31) => A(28), IN3(30) => A(27), IN3(29) => A(26)
                           , IN3(28) => A(25), IN3(27) => A(24), IN3(26) => 
                           A(23), IN3(25) => A(22), IN3(24) => A(21), IN3(23) 
                           => A(20), IN3(22) => A(19), IN3(21) => A(18), 
                           IN3(20) => A(17), IN3(19) => A(16), IN3(18) => A(15)
                           , IN3(17) => A(14), IN3(16) => A(13), IN3(15) => 
                           A(12), IN3(14) => A(11), IN3(13) => A(10), IN3(12) 
                           => A(9), IN3(11) => A(8), IN3(10) => A(7), IN3(9) =>
                           A(6), IN3(8) => A(5), IN3(7) => A(4), IN3(6) => A(3)
                           , IN3(5) => A(2), IN3(4) => A(1), IN3(3) => A(0), 
                           IN3(2) => X_Logic0_port, IN3(1) => X_Logic0_port, 
                           IN3(0) => X_Logic0_port, IN4(63) => 
                           negative_a_60_port, IN4(62) => negative_a_59_port, 
                           IN4(61) => negative_a_58_port, IN4(60) => 
                           negative_a_57_port, IN4(59) => negative_a_56_port, 
                           IN4(58) => negative_a_55_port, IN4(57) => 
                           negative_a_54_port, IN4(56) => negative_a_53_port, 
                           IN4(55) => negative_a_52_port, IN4(54) => 
                           negative_a_51_port, IN4(53) => negative_a_50_port, 
                           IN4(52) => negative_a_49_port, IN4(51) => 
                           negative_a_48_port, IN4(50) => negative_a_47_port, 
                           IN4(49) => negative_a_46_port, IN4(48) => 
                           negative_a_45_port, IN4(47) => negative_a_44_port, 
                           IN4(46) => negative_a_43_port, IN4(45) => 
                           negative_a_42_port, IN4(44) => negative_a_41_port, 
                           IN4(43) => negative_a_40_port, IN4(42) => 
                           negative_a_39_port, IN4(41) => negative_a_38_port, 
                           IN4(40) => negative_a_37_port, IN4(39) => 
                           negative_a_36_port, IN4(38) => negative_a_35_port, 
                           IN4(37) => negative_a_34_port, IN4(36) => n36, 
                           IN4(35) => n33, IN4(34) => negative_a_31_port, 
                           IN4(33) => negative_a_30_port, IN4(32) => 
                           negative_a_29_port, IN4(31) => negative_a_28_port, 
                           IN4(30) => negative_a_27_port, IN4(29) => 
                           negative_a_26_port, IN4(28) => negative_a_25_port, 
                           IN4(27) => negative_a_24_port, IN4(26) => 
                           negative_a_23_port, IN4(25) => negative_a_22_port, 
                           IN4(24) => negative_a_21_port, IN4(23) => 
                           negative_a_20_port, IN4(22) => negative_a_19_port, 
                           IN4(21) => negative_a_18_port, IN4(20) => 
                           negative_a_17_port, IN4(19) => negative_a_16_port, 
                           IN4(18) => negative_a_15_port, IN4(17) => 
                           negative_a_14_port, IN4(16) => negative_a_13_port, 
                           IN4(15) => negative_a_12_port, IN4(14) => 
                           negative_a_11_port, IN4(13) => negative_a_10_port, 
                           IN4(12) => negative_a_9_port, IN4(11) => 
                           negative_a_8_port, IN4(10) => negative_a_7_port, 
                           IN4(9) => negative_a_6_port, IN4(8) => 
                           negative_a_5_port, IN4(7) => negative_a_4_port, 
                           IN4(6) => negative_a_3_port, IN4(5) => 
                           negative_a_2_port, IN4(4) => negative_a_1_port, 
                           IN4(3) => negative_a_0_port, IN4(2) => X_Logic0_port
                           , IN4(1) => X_Logic0_port, IN4(0) => X_Logic0_port, 
                           S(2) => muxs_encoded_signals_1_2_port, S(1) => 
                           muxs_encoded_signals_1_1_port, S(0) => 
                           muxs_encoded_signals_1_0_port, O(63) => 
                           out_imux_1_63_port, O(62) => out_imux_1_62_port, 
                           O(61) => out_imux_1_61_port, O(60) => 
                           out_imux_1_60_port, O(59) => out_imux_1_59_port, 
                           O(58) => out_imux_1_58_port, O(57) => 
                           out_imux_1_57_port, O(56) => out_imux_1_56_port, 
                           O(55) => out_imux_1_55_port, O(54) => 
                           out_imux_1_54_port, O(53) => out_imux_1_53_port, 
                           O(52) => out_imux_1_52_port, O(51) => 
                           out_imux_1_51_port, O(50) => out_imux_1_50_port, 
                           O(49) => out_imux_1_49_port, O(48) => 
                           out_imux_1_48_port, O(47) => out_imux_1_47_port, 
                           O(46) => out_imux_1_46_port, O(45) => 
                           out_imux_1_45_port, O(44) => out_imux_1_44_port, 
                           O(43) => out_imux_1_43_port, O(42) => 
                           out_imux_1_42_port, O(41) => out_imux_1_41_port, 
                           O(40) => out_imux_1_40_port, O(39) => 
                           out_imux_1_39_port, O(38) => out_imux_1_38_port, 
                           O(37) => out_imux_1_37_port, O(36) => 
                           out_imux_1_36_port, O(35) => out_imux_1_35_port, 
                           O(34) => out_imux_1_34_port, O(33) => 
                           out_imux_1_33_port, O(32) => out_imux_1_32_port, 
                           O(31) => out_imux_1_31_port, O(30) => 
                           out_imux_1_30_port, O(29) => out_imux_1_29_port, 
                           O(28) => out_imux_1_28_port, O(27) => 
                           out_imux_1_27_port, O(26) => out_imux_1_26_port, 
                           O(25) => out_imux_1_25_port, O(24) => 
                           out_imux_1_24_port, O(23) => out_imux_1_23_port, 
                           O(22) => out_imux_1_22_port, O(21) => 
                           out_imux_1_21_port, O(20) => out_imux_1_20_port, 
                           O(19) => out_imux_1_19_port, O(18) => 
                           out_imux_1_18_port, O(17) => out_imux_1_17_port, 
                           O(16) => out_imux_1_16_port, O(15) => 
                           out_imux_1_15_port, O(14) => out_imux_1_14_port, 
                           O(13) => out_imux_1_13_port, O(12) => 
                           out_imux_1_12_port, O(11) => out_imux_1_11_port, 
                           O(10) => out_imux_1_10_port, O(9) => 
                           out_imux_1_9_port, O(8) => out_imux_1_8_port, O(7) 
                           => out_imux_1_7_port, O(6) => out_imux_1_6_port, 
                           O(5) => out_imux_1_5_port, O(4) => out_imux_1_4_port
                           , O(3) => out_imux_1_3_port, O(2) => 
                           out_imux_1_2_port, O(1) => out_imux_1_1_port, O(0) 
                           => out_imux_1_0_port);
   ADD64_i_1 : RCA_GENERIC_NBIT64_0 port map( A(63) => out_imux_0_63_port, 
                           A(62) => out_imux_0_62_port, A(61) => 
                           out_imux_0_61_port, A(60) => out_imux_0_60_port, 
                           A(59) => out_imux_0_59_port, A(58) => 
                           out_imux_0_58_port, A(57) => out_imux_0_57_port, 
                           A(56) => out_imux_0_56_port, A(55) => 
                           out_imux_0_55_port, A(54) => out_imux_0_54_port, 
                           A(53) => out_imux_0_53_port, A(52) => 
                           out_imux_0_52_port, A(51) => out_imux_0_51_port, 
                           A(50) => out_imux_0_50_port, A(49) => 
                           out_imux_0_49_port, A(48) => out_imux_0_48_port, 
                           A(47) => out_imux_0_47_port, A(46) => 
                           out_imux_0_46_port, A(45) => out_imux_0_45_port, 
                           A(44) => out_imux_0_44_port, A(43) => 
                           out_imux_0_43_port, A(42) => out_imux_0_42_port, 
                           A(41) => out_imux_0_41_port, A(40) => 
                           out_imux_0_40_port, A(39) => out_imux_0_39_port, 
                           A(38) => out_imux_0_38_port, A(37) => 
                           out_imux_0_37_port, A(36) => out_imux_0_36_port, 
                           A(35) => out_imux_0_35_port, A(34) => 
                           out_imux_0_34_port, A(33) => out_imux_0_33_port, 
                           A(32) => out_imux_0_32_port, A(31) => 
                           out_imux_0_31_port, A(30) => out_imux_0_30_port, 
                           A(29) => out_imux_0_29_port, A(28) => 
                           out_imux_0_28_port, A(27) => out_imux_0_27_port, 
                           A(26) => out_imux_0_26_port, A(25) => 
                           out_imux_0_25_port, A(24) => out_imux_0_24_port, 
                           A(23) => out_imux_0_23_port, A(22) => 
                           out_imux_0_22_port, A(21) => out_imux_0_21_port, 
                           A(20) => out_imux_0_20_port, A(19) => 
                           out_imux_0_19_port, A(18) => out_imux_0_18_port, 
                           A(17) => out_imux_0_17_port, A(16) => 
                           out_imux_0_16_port, A(15) => out_imux_0_15_port, 
                           A(14) => out_imux_0_14_port, A(13) => 
                           out_imux_0_13_port, A(12) => out_imux_0_12_port, 
                           A(11) => out_imux_0_11_port, A(10) => 
                           out_imux_0_10_port, A(9) => out_imux_0_9_port, A(8) 
                           => out_imux_0_8_port, A(7) => out_imux_0_7_port, 
                           A(6) => out_imux_0_6_port, A(5) => out_imux_0_5_port
                           , A(4) => out_imux_0_4_port, A(3) => 
                           out_imux_0_3_port, A(2) => out_imux_0_2_port, A(1) 
                           => out_imux_0_1_port, A(0) => out_imux_0_0_port, 
                           B(63) => out_imux_1_63_port, B(62) => 
                           out_imux_1_62_port, B(61) => out_imux_1_61_port, 
                           B(60) => out_imux_1_60_port, B(59) => 
                           out_imux_1_59_port, B(58) => out_imux_1_58_port, 
                           B(57) => out_imux_1_57_port, B(56) => 
                           out_imux_1_56_port, B(55) => out_imux_1_55_port, 
                           B(54) => out_imux_1_54_port, B(53) => 
                           out_imux_1_53_port, B(52) => out_imux_1_52_port, 
                           B(51) => out_imux_1_51_port, B(50) => 
                           out_imux_1_50_port, B(49) => out_imux_1_49_port, 
                           B(48) => out_imux_1_48_port, B(47) => 
                           out_imux_1_47_port, B(46) => out_imux_1_46_port, 
                           B(45) => out_imux_1_45_port, B(44) => 
                           out_imux_1_44_port, B(43) => out_imux_1_43_port, 
                           B(42) => out_imux_1_42_port, B(41) => 
                           out_imux_1_41_port, B(40) => out_imux_1_40_port, 
                           B(39) => out_imux_1_39_port, B(38) => 
                           out_imux_1_38_port, B(37) => out_imux_1_37_port, 
                           B(36) => out_imux_1_36_port, B(35) => 
                           out_imux_1_35_port, B(34) => out_imux_1_34_port, 
                           B(33) => out_imux_1_33_port, B(32) => 
                           out_imux_1_32_port, B(31) => out_imux_1_31_port, 
                           B(30) => out_imux_1_30_port, B(29) => 
                           out_imux_1_29_port, B(28) => out_imux_1_28_port, 
                           B(27) => out_imux_1_27_port, B(26) => 
                           out_imux_1_26_port, B(25) => out_imux_1_25_port, 
                           B(24) => out_imux_1_24_port, B(23) => 
                           out_imux_1_23_port, B(22) => out_imux_1_22_port, 
                           B(21) => out_imux_1_21_port, B(20) => 
                           out_imux_1_20_port, B(19) => out_imux_1_19_port, 
                           B(18) => out_imux_1_18_port, B(17) => 
                           out_imux_1_17_port, B(16) => out_imux_1_16_port, 
                           B(15) => out_imux_1_15_port, B(14) => 
                           out_imux_1_14_port, B(13) => out_imux_1_13_port, 
                           B(12) => out_imux_1_12_port, B(11) => 
                           out_imux_1_11_port, B(10) => out_imux_1_10_port, 
                           B(9) => out_imux_1_9_port, B(8) => out_imux_1_8_port
                           , B(7) => out_imux_1_7_port, B(6) => 
                           out_imux_1_6_port, B(5) => out_imux_1_5_port, B(4) 
                           => out_imux_1_4_port, B(3) => out_imux_1_3_port, 
                           B(2) => out_imux_1_2_port, B(1) => out_imux_1_1_port
                           , B(0) => out_imux_1_0_port, Ci => X_Logic0_port, 
                           S(63) => predigest_product_1_63_port, S(62) => 
                           predigest_product_1_62_port, S(61) => 
                           predigest_product_1_61_port, S(60) => 
                           predigest_product_1_60_port, S(59) => 
                           predigest_product_1_59_port, S(58) => 
                           predigest_product_1_58_port, S(57) => 
                           predigest_product_1_57_port, S(56) => 
                           predigest_product_1_56_port, S(55) => 
                           predigest_product_1_55_port, S(54) => 
                           predigest_product_1_54_port, S(53) => 
                           predigest_product_1_53_port, S(52) => 
                           predigest_product_1_52_port, S(51) => 
                           predigest_product_1_51_port, S(50) => 
                           predigest_product_1_50_port, S(49) => 
                           predigest_product_1_49_port, S(48) => 
                           predigest_product_1_48_port, S(47) => 
                           predigest_product_1_47_port, S(46) => 
                           predigest_product_1_46_port, S(45) => 
                           predigest_product_1_45_port, S(44) => 
                           predigest_product_1_44_port, S(43) => 
                           predigest_product_1_43_port, S(42) => 
                           predigest_product_1_42_port, S(41) => 
                           predigest_product_1_41_port, S(40) => 
                           predigest_product_1_40_port, S(39) => 
                           predigest_product_1_39_port, S(38) => 
                           predigest_product_1_38_port, S(37) => 
                           predigest_product_1_37_port, S(36) => 
                           predigest_product_1_36_port, S(35) => 
                           predigest_product_1_35_port, S(34) => 
                           predigest_product_1_34_port, S(33) => 
                           predigest_product_1_33_port, S(32) => 
                           predigest_product_1_32_port, S(31) => 
                           predigest_product_1_31_port, S(30) => 
                           predigest_product_1_30_port, S(29) => 
                           predigest_product_1_29_port, S(28) => 
                           predigest_product_1_28_port, S(27) => 
                           predigest_product_1_27_port, S(26) => 
                           predigest_product_1_26_port, S(25) => 
                           predigest_product_1_25_port, S(24) => 
                           predigest_product_1_24_port, S(23) => 
                           predigest_product_1_23_port, S(22) => 
                           predigest_product_1_22_port, S(21) => 
                           predigest_product_1_21_port, S(20) => 
                           predigest_product_1_20_port, S(19) => 
                           predigest_product_1_19_port, S(18) => 
                           predigest_product_1_18_port, S(17) => 
                           predigest_product_1_17_port, S(16) => 
                           predigest_product_1_16_port, S(15) => 
                           predigest_product_1_15_port, S(14) => 
                           predigest_product_1_14_port, S(13) => 
                           predigest_product_1_13_port, S(12) => 
                           predigest_product_1_12_port, S(11) => 
                           predigest_product_1_11_port, S(10) => 
                           predigest_product_1_10_port, S(9) => 
                           predigest_product_1_9_port, S(8) => 
                           predigest_product_1_8_port, S(7) => 
                           predigest_product_1_7_port, S(6) => 
                           predigest_product_1_6_port, S(5) => 
                           predigest_product_1_5_port, S(4) => 
                           predigest_product_1_4_port, S(3) => 
                           predigest_product_1_3_port, S(2) => 
                           predigest_product_1_2_port, S(1) => 
                           predigest_product_1_1_port, S(0) => 
                           predigest_product_1_0_port, Co => n_1092);
   ENC_i_2 : BOOTH_ENCODER_3BIT_18 port map( B(2) => B(5), B(1) => B(4), B(0) 
                           => B(3), ENCODED(2) => muxs_encoded_signals_2_2_port
                           , ENCODED(1) => muxs_encoded_signals_2_1_port, 
                           ENCODED(0) => muxs_encoded_signals_2_0_port);
   MUX_i_2 : MUX51_GENERIC_NBIT64_14 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(31), IN1(51) 
                           => A(31), IN1(50) => A(31), IN1(49) => A(31), 
                           IN1(48) => A(31), IN1(47) => A(31), IN1(46) => A(31)
                           , IN1(45) => A(31), IN1(44) => A(31), IN1(43) => 
                           A(31), IN1(42) => A(31), IN1(41) => A(31), IN1(40) 
                           => A(31), IN1(39) => A(31), IN1(38) => A(31), 
                           IN1(37) => A(31), IN1(36) => A(31), IN1(35) => A(31)
                           , IN1(34) => A(30), IN1(33) => A(29), IN1(32) => 
                           A(28), IN1(31) => A(27), IN1(30) => A(26), IN1(29) 
                           => A(25), IN1(28) => A(24), IN1(27) => A(23), 
                           IN1(26) => A(22), IN1(25) => A(21), IN1(24) => A(20)
                           , IN1(23) => A(19), IN1(22) => A(18), IN1(21) => 
                           A(17), IN1(20) => A(16), IN1(19) => A(15), IN1(18) 
                           => A(14), IN1(17) => A(13), IN1(16) => A(12), 
                           IN1(15) => A(11), IN1(14) => A(10), IN1(13) => A(9),
                           IN1(12) => A(8), IN1(11) => A(7), IN1(10) => A(6), 
                           IN1(9) => A(5), IN1(8) => A(4), IN1(7) => A(3), 
                           IN1(6) => A(2), IN1(5) => A(1), IN1(4) => A(0), 
                           IN1(3) => X_Logic0_port, IN1(2) => X_Logic0_port, 
                           IN1(1) => X_Logic0_port, IN1(0) => X_Logic0_port, 
                           IN2(63) => negative_a_59_port, IN2(62) => 
                           negative_a_58_port, IN2(61) => negative_a_57_port, 
                           IN2(60) => negative_a_56_port, IN2(59) => 
                           negative_a_55_port, IN2(58) => negative_a_54_port, 
                           IN2(57) => negative_a_53_port, IN2(56) => 
                           negative_a_52_port, IN2(55) => negative_a_51_port, 
                           IN2(54) => negative_a_50_port, IN2(53) => 
                           negative_a_49_port, IN2(52) => negative_a_48_port, 
                           IN2(51) => negative_a_47_port, IN2(50) => 
                           negative_a_46_port, IN2(49) => negative_a_45_port, 
                           IN2(48) => negative_a_44_port, IN2(47) => 
                           negative_a_43_port, IN2(46) => negative_a_42_port, 
                           IN2(45) => negative_a_41_port, IN2(44) => 
                           negative_a_40_port, IN2(43) => negative_a_39_port, 
                           IN2(42) => negative_a_38_port, IN2(41) => 
                           negative_a_37_port, IN2(40) => negative_a_36_port, 
                           IN2(39) => negative_a_35_port, IN2(38) => 
                           negative_a_34_port, IN2(37) => n36, IN2(36) => n33, 
                           IN2(35) => negative_a_31_port, IN2(34) => 
                           negative_a_30_port, IN2(33) => negative_a_29_port, 
                           IN2(32) => negative_a_28_port, IN2(31) => 
                           negative_a_27_port, IN2(30) => negative_a_26_port, 
                           IN2(29) => negative_a_25_port, IN2(28) => 
                           negative_a_24_port, IN2(27) => negative_a_23_port, 
                           IN2(26) => negative_a_22_port, IN2(25) => 
                           negative_a_21_port, IN2(24) => negative_a_20_port, 
                           IN2(23) => negative_a_19_port, IN2(22) => 
                           negative_a_18_port, IN2(21) => negative_a_17_port, 
                           IN2(20) => negative_a_16_port, IN2(19) => 
                           negative_a_15_port, IN2(18) => negative_a_14_port, 
                           IN2(17) => negative_a_13_port, IN2(16) => 
                           negative_a_12_port, IN2(15) => negative_a_11_port, 
                           IN2(14) => negative_a_10_port, IN2(13) => 
                           negative_a_9_port, IN2(12) => negative_a_8_port, 
                           IN2(11) => negative_a_7_port, IN2(10) => 
                           negative_a_6_port, IN2(9) => negative_a_5_port, 
                           IN2(8) => negative_a_4_port, IN2(7) => 
                           negative_a_3_port, IN2(6) => negative_a_2_port, 
                           IN2(5) => negative_a_1_port, IN2(4) => 
                           negative_a_0_port, IN2(3) => X_Logic0_port, IN2(2) 
                           => X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) =>
                           X_Logic0_port, IN3(63) => A(31), IN3(62) => A(31), 
                           IN3(61) => A(31), IN3(60) => A(31), IN3(59) => A(31)
                           , IN3(58) => A(31), IN3(57) => A(31), IN3(56) => 
                           A(31), IN3(55) => A(31), IN3(54) => A(31), IN3(53) 
                           => A(31), IN3(52) => A(31), IN3(51) => A(31), 
                           IN3(50) => A(31), IN3(49) => A(31), IN3(48) => A(31)
                           , IN3(47) => A(31), IN3(46) => A(31), IN3(45) => 
                           A(31), IN3(44) => A(31), IN3(43) => A(31), IN3(42) 
                           => A(31), IN3(41) => A(31), IN3(40) => A(31), 
                           IN3(39) => A(31), IN3(38) => A(31), IN3(37) => A(31)
                           , IN3(36) => A(31), IN3(35) => A(30), IN3(34) => 
                           A(29), IN3(33) => A(28), IN3(32) => A(27), IN3(31) 
                           => A(26), IN3(30) => A(25), IN3(29) => A(24), 
                           IN3(28) => A(23), IN3(27) => A(22), IN3(26) => A(21)
                           , IN3(25) => A(20), IN3(24) => A(19), IN3(23) => 
                           A(18), IN3(22) => A(17), IN3(21) => A(16), IN3(20) 
                           => A(15), IN3(19) => A(14), IN3(18) => A(13), 
                           IN3(17) => A(12), IN3(16) => A(11), IN3(15) => A(10)
                           , IN3(14) => A(9), IN3(13) => A(8), IN3(12) => A(7),
                           IN3(11) => A(6), IN3(10) => A(5), IN3(9) => A(4), 
                           IN3(8) => A(3), IN3(7) => A(2), IN3(6) => A(1), 
                           IN3(5) => A(0), IN3(4) => X_Logic0_port, IN3(3) => 
                           X_Logic0_port, IN3(2) => X_Logic0_port, IN3(1) => 
                           X_Logic0_port, IN3(0) => X_Logic0_port, IN4(63) => 
                           negative_a_58_port, IN4(62) => negative_a_57_port, 
                           IN4(61) => negative_a_56_port, IN4(60) => 
                           negative_a_55_port, IN4(59) => negative_a_54_port, 
                           IN4(58) => negative_a_53_port, IN4(57) => 
                           negative_a_52_port, IN4(56) => negative_a_51_port, 
                           IN4(55) => negative_a_50_port, IN4(54) => 
                           negative_a_49_port, IN4(53) => negative_a_48_port, 
                           IN4(52) => negative_a_47_port, IN4(51) => 
                           negative_a_46_port, IN4(50) => negative_a_45_port, 
                           IN4(49) => negative_a_44_port, IN4(48) => 
                           negative_a_43_port, IN4(47) => negative_a_42_port, 
                           IN4(46) => negative_a_41_port, IN4(45) => 
                           negative_a_40_port, IN4(44) => negative_a_39_port, 
                           IN4(43) => negative_a_38_port, IN4(42) => 
                           negative_a_37_port, IN4(41) => negative_a_36_port, 
                           IN4(40) => negative_a_35_port, IN4(39) => 
                           negative_a_34_port, IN4(38) => n36, IN4(37) => n33, 
                           IN4(36) => negative_a_31_port, IN4(35) => 
                           negative_a_30_port, IN4(34) => negative_a_29_port, 
                           IN4(33) => negative_a_28_port, IN4(32) => 
                           negative_a_27_port, IN4(31) => negative_a_26_port, 
                           IN4(30) => negative_a_25_port, IN4(29) => 
                           negative_a_24_port, IN4(28) => negative_a_23_port, 
                           IN4(27) => negative_a_22_port, IN4(26) => 
                           negative_a_21_port, IN4(25) => negative_a_20_port, 
                           IN4(24) => negative_a_19_port, IN4(23) => 
                           negative_a_18_port, IN4(22) => negative_a_17_port, 
                           IN4(21) => negative_a_16_port, IN4(20) => 
                           negative_a_15_port, IN4(19) => negative_a_14_port, 
                           IN4(18) => negative_a_13_port, IN4(17) => 
                           negative_a_12_port, IN4(16) => negative_a_11_port, 
                           IN4(15) => negative_a_10_port, IN4(14) => 
                           negative_a_9_port, IN4(13) => negative_a_8_port, 
                           IN4(12) => negative_a_7_port, IN4(11) => 
                           negative_a_6_port, IN4(10) => negative_a_5_port, 
                           IN4(9) => negative_a_4_port, IN4(8) => 
                           negative_a_3_port, IN4(7) => negative_a_2_port, 
                           IN4(6) => negative_a_1_port, IN4(5) => 
                           negative_a_0_port, IN4(4) => X_Logic0_port, IN4(3) 
                           => X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) =>
                           X_Logic0_port, IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_2_2_port, S(1) => 
                           muxs_encoded_signals_2_1_port, S(0) => 
                           muxs_encoded_signals_2_0_port, O(63) => 
                           out_imux_2_63_port, O(62) => out_imux_2_62_port, 
                           O(61) => out_imux_2_61_port, O(60) => 
                           out_imux_2_60_port, O(59) => out_imux_2_59_port, 
                           O(58) => out_imux_2_58_port, O(57) => 
                           out_imux_2_57_port, O(56) => out_imux_2_56_port, 
                           O(55) => out_imux_2_55_port, O(54) => 
                           out_imux_2_54_port, O(53) => out_imux_2_53_port, 
                           O(52) => out_imux_2_52_port, O(51) => 
                           out_imux_2_51_port, O(50) => out_imux_2_50_port, 
                           O(49) => out_imux_2_49_port, O(48) => 
                           out_imux_2_48_port, O(47) => out_imux_2_47_port, 
                           O(46) => out_imux_2_46_port, O(45) => 
                           out_imux_2_45_port, O(44) => out_imux_2_44_port, 
                           O(43) => out_imux_2_43_port, O(42) => 
                           out_imux_2_42_port, O(41) => out_imux_2_41_port, 
                           O(40) => out_imux_2_40_port, O(39) => 
                           out_imux_2_39_port, O(38) => out_imux_2_38_port, 
                           O(37) => out_imux_2_37_port, O(36) => 
                           out_imux_2_36_port, O(35) => out_imux_2_35_port, 
                           O(34) => out_imux_2_34_port, O(33) => 
                           out_imux_2_33_port, O(32) => out_imux_2_32_port, 
                           O(31) => out_imux_2_31_port, O(30) => 
                           out_imux_2_30_port, O(29) => out_imux_2_29_port, 
                           O(28) => out_imux_2_28_port, O(27) => 
                           out_imux_2_27_port, O(26) => out_imux_2_26_port, 
                           O(25) => out_imux_2_25_port, O(24) => 
                           out_imux_2_24_port, O(23) => out_imux_2_23_port, 
                           O(22) => out_imux_2_22_port, O(21) => 
                           out_imux_2_21_port, O(20) => out_imux_2_20_port, 
                           O(19) => out_imux_2_19_port, O(18) => 
                           out_imux_2_18_port, O(17) => out_imux_2_17_port, 
                           O(16) => out_imux_2_16_port, O(15) => 
                           out_imux_2_15_port, O(14) => out_imux_2_14_port, 
                           O(13) => out_imux_2_13_port, O(12) => 
                           out_imux_2_12_port, O(11) => out_imux_2_11_port, 
                           O(10) => out_imux_2_10_port, O(9) => 
                           out_imux_2_9_port, O(8) => out_imux_2_8_port, O(7) 
                           => out_imux_2_7_port, O(6) => out_imux_2_6_port, 
                           O(5) => out_imux_2_5_port, O(4) => out_imux_2_4_port
                           , O(3) => out_imux_2_3_port, O(2) => 
                           out_imux_2_2_port, O(1) => out_imux_2_1_port, O(0) 
                           => out_imux_2_0_port);
   ADD64_i_2 : RCA_GENERIC_NBIT64_14 port map( A(63) => 
                           predigest_product_1_63_port, A(62) => 
                           predigest_product_1_62_port, A(61) => 
                           predigest_product_1_61_port, A(60) => 
                           predigest_product_1_60_port, A(59) => 
                           predigest_product_1_59_port, A(58) => 
                           predigest_product_1_58_port, A(57) => 
                           predigest_product_1_57_port, A(56) => 
                           predigest_product_1_56_port, A(55) => 
                           predigest_product_1_55_port, A(54) => 
                           predigest_product_1_54_port, A(53) => 
                           predigest_product_1_53_port, A(52) => 
                           predigest_product_1_52_port, A(51) => 
                           predigest_product_1_51_port, A(50) => 
                           predigest_product_1_50_port, A(49) => 
                           predigest_product_1_49_port, A(48) => 
                           predigest_product_1_48_port, A(47) => 
                           predigest_product_1_47_port, A(46) => 
                           predigest_product_1_46_port, A(45) => 
                           predigest_product_1_45_port, A(44) => 
                           predigest_product_1_44_port, A(43) => 
                           predigest_product_1_43_port, A(42) => 
                           predigest_product_1_42_port, A(41) => 
                           predigest_product_1_41_port, A(40) => 
                           predigest_product_1_40_port, A(39) => 
                           predigest_product_1_39_port, A(38) => 
                           predigest_product_1_38_port, A(37) => 
                           predigest_product_1_37_port, A(36) => 
                           predigest_product_1_36_port, A(35) => 
                           predigest_product_1_35_port, A(34) => 
                           predigest_product_1_34_port, A(33) => 
                           predigest_product_1_33_port, A(32) => 
                           predigest_product_1_32_port, A(31) => 
                           predigest_product_1_31_port, A(30) => 
                           predigest_product_1_30_port, A(29) => 
                           predigest_product_1_29_port, A(28) => 
                           predigest_product_1_28_port, A(27) => 
                           predigest_product_1_27_port, A(26) => 
                           predigest_product_1_26_port, A(25) => 
                           predigest_product_1_25_port, A(24) => 
                           predigest_product_1_24_port, A(23) => 
                           predigest_product_1_23_port, A(22) => 
                           predigest_product_1_22_port, A(21) => 
                           predigest_product_1_21_port, A(20) => 
                           predigest_product_1_20_port, A(19) => 
                           predigest_product_1_19_port, A(18) => 
                           predigest_product_1_18_port, A(17) => 
                           predigest_product_1_17_port, A(16) => 
                           predigest_product_1_16_port, A(15) => 
                           predigest_product_1_15_port, A(14) => 
                           predigest_product_1_14_port, A(13) => 
                           predigest_product_1_13_port, A(12) => 
                           predigest_product_1_12_port, A(11) => 
                           predigest_product_1_11_port, A(10) => 
                           predigest_product_1_10_port, A(9) => 
                           predigest_product_1_9_port, A(8) => 
                           predigest_product_1_8_port, A(7) => 
                           predigest_product_1_7_port, A(6) => 
                           predigest_product_1_6_port, A(5) => 
                           predigest_product_1_5_port, A(4) => 
                           predigest_product_1_4_port, A(3) => 
                           predigest_product_1_3_port, A(2) => 
                           predigest_product_1_2_port, A(1) => 
                           predigest_product_1_1_port, A(0) => 
                           predigest_product_1_0_port, B(63) => 
                           out_imux_2_63_port, B(62) => out_imux_2_62_port, 
                           B(61) => out_imux_2_61_port, B(60) => 
                           out_imux_2_60_port, B(59) => out_imux_2_59_port, 
                           B(58) => out_imux_2_58_port, B(57) => 
                           out_imux_2_57_port, B(56) => out_imux_2_56_port, 
                           B(55) => out_imux_2_55_port, B(54) => 
                           out_imux_2_54_port, B(53) => out_imux_2_53_port, 
                           B(52) => out_imux_2_52_port, B(51) => 
                           out_imux_2_51_port, B(50) => out_imux_2_50_port, 
                           B(49) => out_imux_2_49_port, B(48) => 
                           out_imux_2_48_port, B(47) => out_imux_2_47_port, 
                           B(46) => out_imux_2_46_port, B(45) => 
                           out_imux_2_45_port, B(44) => out_imux_2_44_port, 
                           B(43) => out_imux_2_43_port, B(42) => 
                           out_imux_2_42_port, B(41) => out_imux_2_41_port, 
                           B(40) => out_imux_2_40_port, B(39) => 
                           out_imux_2_39_port, B(38) => out_imux_2_38_port, 
                           B(37) => out_imux_2_37_port, B(36) => 
                           out_imux_2_36_port, B(35) => out_imux_2_35_port, 
                           B(34) => out_imux_2_34_port, B(33) => 
                           out_imux_2_33_port, B(32) => out_imux_2_32_port, 
                           B(31) => out_imux_2_31_port, B(30) => 
                           out_imux_2_30_port, B(29) => out_imux_2_29_port, 
                           B(28) => out_imux_2_28_port, B(27) => 
                           out_imux_2_27_port, B(26) => out_imux_2_26_port, 
                           B(25) => out_imux_2_25_port, B(24) => 
                           out_imux_2_24_port, B(23) => out_imux_2_23_port, 
                           B(22) => out_imux_2_22_port, B(21) => 
                           out_imux_2_21_port, B(20) => out_imux_2_20_port, 
                           B(19) => out_imux_2_19_port, B(18) => 
                           out_imux_2_18_port, B(17) => out_imux_2_17_port, 
                           B(16) => out_imux_2_16_port, B(15) => 
                           out_imux_2_15_port, B(14) => out_imux_2_14_port, 
                           B(13) => out_imux_2_13_port, B(12) => 
                           out_imux_2_12_port, B(11) => out_imux_2_11_port, 
                           B(10) => out_imux_2_10_port, B(9) => 
                           out_imux_2_9_port, B(8) => out_imux_2_8_port, B(7) 
                           => out_imux_2_7_port, B(6) => out_imux_2_6_port, 
                           B(5) => out_imux_2_5_port, B(4) => out_imux_2_4_port
                           , B(3) => out_imux_2_3_port, B(2) => 
                           out_imux_2_2_port, B(1) => out_imux_2_1_port, B(0) 
                           => out_imux_2_0_port, Ci => X_Logic0_port, S(63) => 
                           predigest_product_2_63_port, S(62) => 
                           predigest_product_2_62_port, S(61) => 
                           predigest_product_2_61_port, S(60) => 
                           predigest_product_2_60_port, S(59) => 
                           predigest_product_2_59_port, S(58) => 
                           predigest_product_2_58_port, S(57) => 
                           predigest_product_2_57_port, S(56) => 
                           predigest_product_2_56_port, S(55) => 
                           predigest_product_2_55_port, S(54) => 
                           predigest_product_2_54_port, S(53) => 
                           predigest_product_2_53_port, S(52) => 
                           predigest_product_2_52_port, S(51) => 
                           predigest_product_2_51_port, S(50) => 
                           predigest_product_2_50_port, S(49) => 
                           predigest_product_2_49_port, S(48) => 
                           predigest_product_2_48_port, S(47) => 
                           predigest_product_2_47_port, S(46) => 
                           predigest_product_2_46_port, S(45) => 
                           predigest_product_2_45_port, S(44) => 
                           predigest_product_2_44_port, S(43) => 
                           predigest_product_2_43_port, S(42) => 
                           predigest_product_2_42_port, S(41) => 
                           predigest_product_2_41_port, S(40) => 
                           predigest_product_2_40_port, S(39) => 
                           predigest_product_2_39_port, S(38) => 
                           predigest_product_2_38_port, S(37) => 
                           predigest_product_2_37_port, S(36) => 
                           predigest_product_2_36_port, S(35) => 
                           predigest_product_2_35_port, S(34) => 
                           predigest_product_2_34_port, S(33) => 
                           predigest_product_2_33_port, S(32) => 
                           predigest_product_2_32_port, S(31) => 
                           predigest_product_2_31_port, S(30) => 
                           predigest_product_2_30_port, S(29) => 
                           predigest_product_2_29_port, S(28) => 
                           predigest_product_2_28_port, S(27) => 
                           predigest_product_2_27_port, S(26) => 
                           predigest_product_2_26_port, S(25) => 
                           predigest_product_2_25_port, S(24) => 
                           predigest_product_2_24_port, S(23) => 
                           predigest_product_2_23_port, S(22) => 
                           predigest_product_2_22_port, S(21) => 
                           predigest_product_2_21_port, S(20) => 
                           predigest_product_2_20_port, S(19) => 
                           predigest_product_2_19_port, S(18) => 
                           predigest_product_2_18_port, S(17) => 
                           predigest_product_2_17_port, S(16) => 
                           predigest_product_2_16_port, S(15) => 
                           predigest_product_2_15_port, S(14) => 
                           predigest_product_2_14_port, S(13) => 
                           predigest_product_2_13_port, S(12) => 
                           predigest_product_2_12_port, S(11) => 
                           predigest_product_2_11_port, S(10) => 
                           predigest_product_2_10_port, S(9) => 
                           predigest_product_2_9_port, S(8) => 
                           predigest_product_2_8_port, S(7) => 
                           predigest_product_2_7_port, S(6) => 
                           predigest_product_2_6_port, S(5) => 
                           predigest_product_2_5_port, S(4) => 
                           predigest_product_2_4_port, S(3) => 
                           predigest_product_2_3_port, S(2) => 
                           predigest_product_2_2_port, S(1) => 
                           predigest_product_2_1_port, S(0) => 
                           predigest_product_2_0_port, Co => n_1093);
   ENC_i_3 : BOOTH_ENCODER_3BIT_17 port map( B(2) => B(7), B(1) => B(6), B(0) 
                           => B(5), ENCODED(2) => muxs_encoded_signals_3_2_port
                           , ENCODED(1) => muxs_encoded_signals_3_1_port, 
                           ENCODED(0) => muxs_encoded_signals_3_0_port);
   MUX_i_3 : MUX51_GENERIC_NBIT64_13 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(31), IN1(51) 
                           => A(31), IN1(50) => A(31), IN1(49) => A(31), 
                           IN1(48) => A(31), IN1(47) => A(31), IN1(46) => A(31)
                           , IN1(45) => A(31), IN1(44) => A(31), IN1(43) => 
                           A(31), IN1(42) => A(31), IN1(41) => A(31), IN1(40) 
                           => A(31), IN1(39) => A(31), IN1(38) => A(31), 
                           IN1(37) => A(31), IN1(36) => A(30), IN1(35) => A(29)
                           , IN1(34) => A(28), IN1(33) => A(27), IN1(32) => 
                           A(26), IN1(31) => A(25), IN1(30) => A(24), IN1(29) 
                           => A(23), IN1(28) => A(22), IN1(27) => A(21), 
                           IN1(26) => A(20), IN1(25) => A(19), IN1(24) => A(18)
                           , IN1(23) => A(17), IN1(22) => A(16), IN1(21) => 
                           A(15), IN1(20) => A(14), IN1(19) => A(13), IN1(18) 
                           => A(12), IN1(17) => A(11), IN1(16) => A(10), 
                           IN1(15) => A(9), IN1(14) => A(8), IN1(13) => A(7), 
                           IN1(12) => A(6), IN1(11) => A(5), IN1(10) => A(4), 
                           IN1(9) => A(3), IN1(8) => A(2), IN1(7) => A(1), 
                           IN1(6) => A(0), IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(63) => negative_a_57_port, 
                           IN2(62) => negative_a_56_port, IN2(61) => 
                           negative_a_55_port, IN2(60) => negative_a_54_port, 
                           IN2(59) => negative_a_53_port, IN2(58) => 
                           negative_a_52_port, IN2(57) => negative_a_51_port, 
                           IN2(56) => negative_a_50_port, IN2(55) => 
                           negative_a_49_port, IN2(54) => negative_a_48_port, 
                           IN2(53) => negative_a_47_port, IN2(52) => 
                           negative_a_46_port, IN2(51) => negative_a_45_port, 
                           IN2(50) => negative_a_44_port, IN2(49) => 
                           negative_a_43_port, IN2(48) => negative_a_42_port, 
                           IN2(47) => negative_a_41_port, IN2(46) => 
                           negative_a_40_port, IN2(45) => negative_a_39_port, 
                           IN2(44) => negative_a_38_port, IN2(43) => 
                           negative_a_37_port, IN2(42) => negative_a_36_port, 
                           IN2(41) => negative_a_35_port, IN2(40) => 
                           negative_a_34_port, IN2(39) => n36, IN2(38) => n33, 
                           IN2(37) => negative_a_31_port, IN2(36) => 
                           negative_a_30_port, IN2(35) => negative_a_29_port, 
                           IN2(34) => negative_a_28_port, IN2(33) => 
                           negative_a_27_port, IN2(32) => negative_a_26_port, 
                           IN2(31) => negative_a_25_port, IN2(30) => 
                           negative_a_24_port, IN2(29) => negative_a_23_port, 
                           IN2(28) => negative_a_22_port, IN2(27) => 
                           negative_a_21_port, IN2(26) => negative_a_20_port, 
                           IN2(25) => negative_a_19_port, IN2(24) => 
                           negative_a_18_port, IN2(23) => negative_a_17_port, 
                           IN2(22) => negative_a_16_port, IN2(21) => 
                           negative_a_15_port, IN2(20) => negative_a_14_port, 
                           IN2(19) => negative_a_13_port, IN2(18) => 
                           negative_a_12_port, IN2(17) => negative_a_11_port, 
                           IN2(16) => negative_a_10_port, IN2(15) => 
                           negative_a_9_port, IN2(14) => negative_a_8_port, 
                           IN2(13) => negative_a_7_port, IN2(12) => 
                           negative_a_6_port, IN2(11) => negative_a_5_port, 
                           IN2(10) => negative_a_4_port, IN2(9) => 
                           negative_a_3_port, IN2(8) => negative_a_2_port, 
                           IN2(7) => negative_a_1_port, IN2(6) => 
                           negative_a_0_port, IN2(5) => X_Logic0_port, IN2(4) 
                           => X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) =>
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(63) => A(31), IN3(62) => A(31), 
                           IN3(61) => A(31), IN3(60) => A(31), IN3(59) => A(31)
                           , IN3(58) => A(31), IN3(57) => A(31), IN3(56) => 
                           A(31), IN3(55) => A(31), IN3(54) => A(31), IN3(53) 
                           => A(31), IN3(52) => A(31), IN3(51) => A(31), 
                           IN3(50) => A(31), IN3(49) => A(31), IN3(48) => A(31)
                           , IN3(47) => A(31), IN3(46) => A(31), IN3(45) => 
                           A(31), IN3(44) => A(31), IN3(43) => A(31), IN3(42) 
                           => A(31), IN3(41) => A(31), IN3(40) => A(31), 
                           IN3(39) => A(31), IN3(38) => A(31), IN3(37) => A(30)
                           , IN3(36) => A(29), IN3(35) => A(28), IN3(34) => 
                           A(27), IN3(33) => A(26), IN3(32) => A(25), IN3(31) 
                           => A(24), IN3(30) => A(23), IN3(29) => A(22), 
                           IN3(28) => A(21), IN3(27) => A(20), IN3(26) => A(19)
                           , IN3(25) => A(18), IN3(24) => A(17), IN3(23) => 
                           A(16), IN3(22) => A(15), IN3(21) => A(14), IN3(20) 
                           => A(13), IN3(19) => A(12), IN3(18) => A(11), 
                           IN3(17) => A(10), IN3(16) => A(9), IN3(15) => A(8), 
                           IN3(14) => A(7), IN3(13) => A(6), IN3(12) => A(5), 
                           IN3(11) => A(4), IN3(10) => A(3), IN3(9) => A(2), 
                           IN3(8) => A(1), IN3(7) => A(0), IN3(6) => 
                           X_Logic0_port, IN3(5) => X_Logic0_port, IN3(4) => 
                           X_Logic0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(63) => negative_a_56_port, 
                           IN4(62) => negative_a_55_port, IN4(61) => 
                           negative_a_54_port, IN4(60) => negative_a_53_port, 
                           IN4(59) => negative_a_52_port, IN4(58) => 
                           negative_a_51_port, IN4(57) => negative_a_50_port, 
                           IN4(56) => negative_a_49_port, IN4(55) => 
                           negative_a_48_port, IN4(54) => negative_a_47_port, 
                           IN4(53) => negative_a_46_port, IN4(52) => 
                           negative_a_45_port, IN4(51) => negative_a_44_port, 
                           IN4(50) => negative_a_43_port, IN4(49) => 
                           negative_a_42_port, IN4(48) => negative_a_41_port, 
                           IN4(47) => negative_a_40_port, IN4(46) => 
                           negative_a_39_port, IN4(45) => negative_a_38_port, 
                           IN4(44) => negative_a_37_port, IN4(43) => 
                           negative_a_36_port, IN4(42) => negative_a_35_port, 
                           IN4(41) => negative_a_34_port, IN4(40) => n36, 
                           IN4(39) => n33, IN4(38) => negative_a_31_port, 
                           IN4(37) => negative_a_30_port, IN4(36) => 
                           negative_a_29_port, IN4(35) => negative_a_28_port, 
                           IN4(34) => negative_a_27_port, IN4(33) => 
                           negative_a_26_port, IN4(32) => negative_a_25_port, 
                           IN4(31) => negative_a_24_port, IN4(30) => 
                           negative_a_23_port, IN4(29) => negative_a_22_port, 
                           IN4(28) => negative_a_21_port, IN4(27) => 
                           negative_a_20_port, IN4(26) => negative_a_19_port, 
                           IN4(25) => negative_a_18_port, IN4(24) => 
                           negative_a_17_port, IN4(23) => negative_a_16_port, 
                           IN4(22) => negative_a_15_port, IN4(21) => 
                           negative_a_14_port, IN4(20) => negative_a_13_port, 
                           IN4(19) => negative_a_12_port, IN4(18) => 
                           negative_a_11_port, IN4(17) => negative_a_10_port, 
                           IN4(16) => negative_a_9_port, IN4(15) => 
                           negative_a_8_port, IN4(14) => negative_a_7_port, 
                           IN4(13) => negative_a_6_port, IN4(12) => 
                           negative_a_5_port, IN4(11) => negative_a_4_port, 
                           IN4(10) => negative_a_3_port, IN4(9) => 
                           negative_a_2_port, IN4(8) => negative_a_1_port, 
                           IN4(7) => negative_a_0_port, IN4(6) => X_Logic0_port
                           , IN4(5) => X_Logic0_port, IN4(4) => X_Logic0_port, 
                           IN4(3) => X_Logic0_port, IN4(2) => X_Logic0_port, 
                           IN4(1) => X_Logic0_port, IN4(0) => X_Logic0_port, 
                           S(2) => muxs_encoded_signals_3_2_port, S(1) => 
                           muxs_encoded_signals_3_1_port, S(0) => 
                           muxs_encoded_signals_3_0_port, O(63) => 
                           out_imux_3_63_port, O(62) => out_imux_3_62_port, 
                           O(61) => out_imux_3_61_port, O(60) => 
                           out_imux_3_60_port, O(59) => out_imux_3_59_port, 
                           O(58) => out_imux_3_58_port, O(57) => 
                           out_imux_3_57_port, O(56) => out_imux_3_56_port, 
                           O(55) => out_imux_3_55_port, O(54) => 
                           out_imux_3_54_port, O(53) => out_imux_3_53_port, 
                           O(52) => out_imux_3_52_port, O(51) => 
                           out_imux_3_51_port, O(50) => out_imux_3_50_port, 
                           O(49) => out_imux_3_49_port, O(48) => 
                           out_imux_3_48_port, O(47) => out_imux_3_47_port, 
                           O(46) => out_imux_3_46_port, O(45) => 
                           out_imux_3_45_port, O(44) => out_imux_3_44_port, 
                           O(43) => out_imux_3_43_port, O(42) => 
                           out_imux_3_42_port, O(41) => out_imux_3_41_port, 
                           O(40) => out_imux_3_40_port, O(39) => 
                           out_imux_3_39_port, O(38) => out_imux_3_38_port, 
                           O(37) => out_imux_3_37_port, O(36) => 
                           out_imux_3_36_port, O(35) => out_imux_3_35_port, 
                           O(34) => out_imux_3_34_port, O(33) => 
                           out_imux_3_33_port, O(32) => out_imux_3_32_port, 
                           O(31) => out_imux_3_31_port, O(30) => 
                           out_imux_3_30_port, O(29) => out_imux_3_29_port, 
                           O(28) => out_imux_3_28_port, O(27) => 
                           out_imux_3_27_port, O(26) => out_imux_3_26_port, 
                           O(25) => out_imux_3_25_port, O(24) => 
                           out_imux_3_24_port, O(23) => out_imux_3_23_port, 
                           O(22) => out_imux_3_22_port, O(21) => 
                           out_imux_3_21_port, O(20) => out_imux_3_20_port, 
                           O(19) => out_imux_3_19_port, O(18) => 
                           out_imux_3_18_port, O(17) => out_imux_3_17_port, 
                           O(16) => out_imux_3_16_port, O(15) => 
                           out_imux_3_15_port, O(14) => out_imux_3_14_port, 
                           O(13) => out_imux_3_13_port, O(12) => 
                           out_imux_3_12_port, O(11) => out_imux_3_11_port, 
                           O(10) => out_imux_3_10_port, O(9) => 
                           out_imux_3_9_port, O(8) => out_imux_3_8_port, O(7) 
                           => out_imux_3_7_port, O(6) => out_imux_3_6_port, 
                           O(5) => out_imux_3_5_port, O(4) => out_imux_3_4_port
                           , O(3) => out_imux_3_3_port, O(2) => 
                           out_imux_3_2_port, O(1) => out_imux_3_1_port, O(0) 
                           => out_imux_3_0_port);
   ADD64_i_3 : RCA_GENERIC_NBIT64_13 port map( A(63) => 
                           predigest_product_2_63_port, A(62) => 
                           predigest_product_2_62_port, A(61) => 
                           predigest_product_2_61_port, A(60) => 
                           predigest_product_2_60_port, A(59) => 
                           predigest_product_2_59_port, A(58) => 
                           predigest_product_2_58_port, A(57) => 
                           predigest_product_2_57_port, A(56) => 
                           predigest_product_2_56_port, A(55) => 
                           predigest_product_2_55_port, A(54) => 
                           predigest_product_2_54_port, A(53) => 
                           predigest_product_2_53_port, A(52) => 
                           predigest_product_2_52_port, A(51) => 
                           predigest_product_2_51_port, A(50) => 
                           predigest_product_2_50_port, A(49) => 
                           predigest_product_2_49_port, A(48) => 
                           predigest_product_2_48_port, A(47) => 
                           predigest_product_2_47_port, A(46) => 
                           predigest_product_2_46_port, A(45) => 
                           predigest_product_2_45_port, A(44) => 
                           predigest_product_2_44_port, A(43) => 
                           predigest_product_2_43_port, A(42) => 
                           predigest_product_2_42_port, A(41) => 
                           predigest_product_2_41_port, A(40) => 
                           predigest_product_2_40_port, A(39) => 
                           predigest_product_2_39_port, A(38) => 
                           predigest_product_2_38_port, A(37) => 
                           predigest_product_2_37_port, A(36) => 
                           predigest_product_2_36_port, A(35) => 
                           predigest_product_2_35_port, A(34) => 
                           predigest_product_2_34_port, A(33) => 
                           predigest_product_2_33_port, A(32) => 
                           predigest_product_2_32_port, A(31) => 
                           predigest_product_2_31_port, A(30) => 
                           predigest_product_2_30_port, A(29) => 
                           predigest_product_2_29_port, A(28) => 
                           predigest_product_2_28_port, A(27) => 
                           predigest_product_2_27_port, A(26) => 
                           predigest_product_2_26_port, A(25) => 
                           predigest_product_2_25_port, A(24) => 
                           predigest_product_2_24_port, A(23) => 
                           predigest_product_2_23_port, A(22) => 
                           predigest_product_2_22_port, A(21) => 
                           predigest_product_2_21_port, A(20) => 
                           predigest_product_2_20_port, A(19) => 
                           predigest_product_2_19_port, A(18) => 
                           predigest_product_2_18_port, A(17) => 
                           predigest_product_2_17_port, A(16) => 
                           predigest_product_2_16_port, A(15) => 
                           predigest_product_2_15_port, A(14) => 
                           predigest_product_2_14_port, A(13) => 
                           predigest_product_2_13_port, A(12) => 
                           predigest_product_2_12_port, A(11) => 
                           predigest_product_2_11_port, A(10) => 
                           predigest_product_2_10_port, A(9) => 
                           predigest_product_2_9_port, A(8) => 
                           predigest_product_2_8_port, A(7) => 
                           predigest_product_2_7_port, A(6) => 
                           predigest_product_2_6_port, A(5) => 
                           predigest_product_2_5_port, A(4) => 
                           predigest_product_2_4_port, A(3) => 
                           predigest_product_2_3_port, A(2) => 
                           predigest_product_2_2_port, A(1) => 
                           predigest_product_2_1_port, A(0) => 
                           predigest_product_2_0_port, B(63) => 
                           out_imux_3_63_port, B(62) => out_imux_3_62_port, 
                           B(61) => out_imux_3_61_port, B(60) => 
                           out_imux_3_60_port, B(59) => out_imux_3_59_port, 
                           B(58) => out_imux_3_58_port, B(57) => 
                           out_imux_3_57_port, B(56) => out_imux_3_56_port, 
                           B(55) => out_imux_3_55_port, B(54) => 
                           out_imux_3_54_port, B(53) => out_imux_3_53_port, 
                           B(52) => out_imux_3_52_port, B(51) => 
                           out_imux_3_51_port, B(50) => out_imux_3_50_port, 
                           B(49) => out_imux_3_49_port, B(48) => 
                           out_imux_3_48_port, B(47) => out_imux_3_47_port, 
                           B(46) => out_imux_3_46_port, B(45) => 
                           out_imux_3_45_port, B(44) => out_imux_3_44_port, 
                           B(43) => out_imux_3_43_port, B(42) => 
                           out_imux_3_42_port, B(41) => out_imux_3_41_port, 
                           B(40) => out_imux_3_40_port, B(39) => 
                           out_imux_3_39_port, B(38) => out_imux_3_38_port, 
                           B(37) => out_imux_3_37_port, B(36) => 
                           out_imux_3_36_port, B(35) => out_imux_3_35_port, 
                           B(34) => out_imux_3_34_port, B(33) => 
                           out_imux_3_33_port, B(32) => out_imux_3_32_port, 
                           B(31) => out_imux_3_31_port, B(30) => 
                           out_imux_3_30_port, B(29) => out_imux_3_29_port, 
                           B(28) => out_imux_3_28_port, B(27) => 
                           out_imux_3_27_port, B(26) => out_imux_3_26_port, 
                           B(25) => out_imux_3_25_port, B(24) => 
                           out_imux_3_24_port, B(23) => out_imux_3_23_port, 
                           B(22) => out_imux_3_22_port, B(21) => 
                           out_imux_3_21_port, B(20) => out_imux_3_20_port, 
                           B(19) => out_imux_3_19_port, B(18) => 
                           out_imux_3_18_port, B(17) => out_imux_3_17_port, 
                           B(16) => out_imux_3_16_port, B(15) => 
                           out_imux_3_15_port, B(14) => out_imux_3_14_port, 
                           B(13) => out_imux_3_13_port, B(12) => 
                           out_imux_3_12_port, B(11) => out_imux_3_11_port, 
                           B(10) => out_imux_3_10_port, B(9) => 
                           out_imux_3_9_port, B(8) => out_imux_3_8_port, B(7) 
                           => out_imux_3_7_port, B(6) => out_imux_3_6_port, 
                           B(5) => out_imux_3_5_port, B(4) => out_imux_3_4_port
                           , B(3) => out_imux_3_3_port, B(2) => 
                           out_imux_3_2_port, B(1) => out_imux_3_1_port, B(0) 
                           => out_imux_3_0_port, Ci => X_Logic0_port, S(63) => 
                           predigest_product_3_63_port, S(62) => 
                           predigest_product_3_62_port, S(61) => 
                           predigest_product_3_61_port, S(60) => 
                           predigest_product_3_60_port, S(59) => 
                           predigest_product_3_59_port, S(58) => 
                           predigest_product_3_58_port, S(57) => 
                           predigest_product_3_57_port, S(56) => 
                           predigest_product_3_56_port, S(55) => 
                           predigest_product_3_55_port, S(54) => 
                           predigest_product_3_54_port, S(53) => 
                           predigest_product_3_53_port, S(52) => 
                           predigest_product_3_52_port, S(51) => 
                           predigest_product_3_51_port, S(50) => 
                           predigest_product_3_50_port, S(49) => 
                           predigest_product_3_49_port, S(48) => 
                           predigest_product_3_48_port, S(47) => 
                           predigest_product_3_47_port, S(46) => 
                           predigest_product_3_46_port, S(45) => 
                           predigest_product_3_45_port, S(44) => 
                           predigest_product_3_44_port, S(43) => 
                           predigest_product_3_43_port, S(42) => 
                           predigest_product_3_42_port, S(41) => 
                           predigest_product_3_41_port, S(40) => 
                           predigest_product_3_40_port, S(39) => 
                           predigest_product_3_39_port, S(38) => 
                           predigest_product_3_38_port, S(37) => 
                           predigest_product_3_37_port, S(36) => 
                           predigest_product_3_36_port, S(35) => 
                           predigest_product_3_35_port, S(34) => 
                           predigest_product_3_34_port, S(33) => 
                           predigest_product_3_33_port, S(32) => 
                           predigest_product_3_32_port, S(31) => 
                           predigest_product_3_31_port, S(30) => 
                           predigest_product_3_30_port, S(29) => 
                           predigest_product_3_29_port, S(28) => 
                           predigest_product_3_28_port, S(27) => 
                           predigest_product_3_27_port, S(26) => 
                           predigest_product_3_26_port, S(25) => 
                           predigest_product_3_25_port, S(24) => 
                           predigest_product_3_24_port, S(23) => 
                           predigest_product_3_23_port, S(22) => 
                           predigest_product_3_22_port, S(21) => 
                           predigest_product_3_21_port, S(20) => 
                           predigest_product_3_20_port, S(19) => 
                           predigest_product_3_19_port, S(18) => 
                           predigest_product_3_18_port, S(17) => 
                           predigest_product_3_17_port, S(16) => 
                           predigest_product_3_16_port, S(15) => 
                           predigest_product_3_15_port, S(14) => 
                           predigest_product_3_14_port, S(13) => 
                           predigest_product_3_13_port, S(12) => 
                           predigest_product_3_12_port, S(11) => 
                           predigest_product_3_11_port, S(10) => 
                           predigest_product_3_10_port, S(9) => 
                           predigest_product_3_9_port, S(8) => 
                           predigest_product_3_8_port, S(7) => 
                           predigest_product_3_7_port, S(6) => 
                           predigest_product_3_6_port, S(5) => 
                           predigest_product_3_5_port, S(4) => 
                           predigest_product_3_4_port, S(3) => 
                           predigest_product_3_3_port, S(2) => 
                           predigest_product_3_2_port, S(1) => 
                           predigest_product_3_1_port, S(0) => 
                           predigest_product_3_0_port, Co => n_1094);
   ENC_i_4 : BOOTH_ENCODER_3BIT_16 port map( B(2) => B(9), B(1) => B(8), B(0) 
                           => B(7), ENCODED(2) => muxs_encoded_signals_4_2_port
                           , ENCODED(1) => muxs_encoded_signals_4_1_port, 
                           ENCODED(0) => muxs_encoded_signals_4_0_port);
   MUX_i_4 : MUX51_GENERIC_NBIT64_12 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(31), IN1(51) 
                           => A(31), IN1(50) => A(31), IN1(49) => A(31), 
                           IN1(48) => A(31), IN1(47) => A(31), IN1(46) => A(31)
                           , IN1(45) => A(31), IN1(44) => A(31), IN1(43) => 
                           A(31), IN1(42) => A(31), IN1(41) => A(31), IN1(40) 
                           => A(31), IN1(39) => A(31), IN1(38) => A(30), 
                           IN1(37) => A(29), IN1(36) => A(28), IN1(35) => A(27)
                           , IN1(34) => A(26), IN1(33) => A(25), IN1(32) => 
                           A(24), IN1(31) => A(23), IN1(30) => A(22), IN1(29) 
                           => A(21), IN1(28) => A(20), IN1(27) => A(19), 
                           IN1(26) => A(18), IN1(25) => A(17), IN1(24) => A(16)
                           , IN1(23) => A(15), IN1(22) => A(14), IN1(21) => 
                           A(13), IN1(20) => A(12), IN1(19) => A(11), IN1(18) 
                           => A(10), IN1(17) => A(9), IN1(16) => A(8), IN1(15) 
                           => A(7), IN1(14) => A(6), IN1(13) => A(5), IN1(12) 
                           => A(4), IN1(11) => A(3), IN1(10) => A(2), IN1(9) =>
                           A(1), IN1(8) => A(0), IN1(7) => X_Logic0_port, 
                           IN1(6) => X_Logic0_port, IN1(5) => X_Logic0_port, 
                           IN1(4) => X_Logic0_port, IN1(3) => X_Logic0_port, 
                           IN1(2) => X_Logic0_port, IN1(1) => X_Logic0_port, 
                           IN1(0) => X_Logic0_port, IN2(63) => 
                           negative_a_55_port, IN2(62) => negative_a_54_port, 
                           IN2(61) => negative_a_53_port, IN2(60) => 
                           negative_a_52_port, IN2(59) => negative_a_51_port, 
                           IN2(58) => negative_a_50_port, IN2(57) => 
                           negative_a_49_port, IN2(56) => negative_a_48_port, 
                           IN2(55) => negative_a_47_port, IN2(54) => 
                           negative_a_46_port, IN2(53) => negative_a_45_port, 
                           IN2(52) => negative_a_44_port, IN2(51) => 
                           negative_a_43_port, IN2(50) => negative_a_42_port, 
                           IN2(49) => negative_a_41_port, IN2(48) => 
                           negative_a_40_port, IN2(47) => negative_a_39_port, 
                           IN2(46) => negative_a_38_port, IN2(45) => 
                           negative_a_37_port, IN2(44) => negative_a_36_port, 
                           IN2(43) => negative_a_35_port, IN2(42) => 
                           negative_a_34_port, IN2(41) => n36, IN2(40) => n33, 
                           IN2(39) => negative_a_31_port, IN2(38) => 
                           negative_a_30_port, IN2(37) => negative_a_29_port, 
                           IN2(36) => negative_a_28_port, IN2(35) => 
                           negative_a_27_port, IN2(34) => negative_a_26_port, 
                           IN2(33) => negative_a_25_port, IN2(32) => 
                           negative_a_24_port, IN2(31) => negative_a_23_port, 
                           IN2(30) => negative_a_22_port, IN2(29) => 
                           negative_a_21_port, IN2(28) => negative_a_20_port, 
                           IN2(27) => negative_a_19_port, IN2(26) => 
                           negative_a_18_port, IN2(25) => negative_a_17_port, 
                           IN2(24) => negative_a_16_port, IN2(23) => 
                           negative_a_15_port, IN2(22) => negative_a_14_port, 
                           IN2(21) => negative_a_13_port, IN2(20) => 
                           negative_a_12_port, IN2(19) => negative_a_11_port, 
                           IN2(18) => negative_a_10_port, IN2(17) => 
                           negative_a_9_port, IN2(16) => negative_a_8_port, 
                           IN2(15) => negative_a_7_port, IN2(14) => 
                           negative_a_6_port, IN2(13) => negative_a_5_port, 
                           IN2(12) => negative_a_4_port, IN2(11) => 
                           negative_a_3_port, IN2(10) => negative_a_2_port, 
                           IN2(9) => negative_a_1_port, IN2(8) => 
                           negative_a_0_port, IN2(7) => X_Logic0_port, IN2(6) 
                           => X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) =>
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(63) => A(31), IN3(62) => A(31), 
                           IN3(61) => A(31), IN3(60) => A(31), IN3(59) => A(31)
                           , IN3(58) => A(31), IN3(57) => A(31), IN3(56) => 
                           A(31), IN3(55) => A(31), IN3(54) => A(31), IN3(53) 
                           => A(31), IN3(52) => A(31), IN3(51) => A(31), 
                           IN3(50) => A(31), IN3(49) => A(31), IN3(48) => A(31)
                           , IN3(47) => A(31), IN3(46) => A(31), IN3(45) => 
                           A(31), IN3(44) => A(31), IN3(43) => A(31), IN3(42) 
                           => A(31), IN3(41) => A(31), IN3(40) => A(31), 
                           IN3(39) => A(30), IN3(38) => A(29), IN3(37) => A(28)
                           , IN3(36) => A(27), IN3(35) => A(26), IN3(34) => 
                           A(25), IN3(33) => A(24), IN3(32) => A(23), IN3(31) 
                           => A(22), IN3(30) => A(21), IN3(29) => A(20), 
                           IN3(28) => A(19), IN3(27) => A(18), IN3(26) => A(17)
                           , IN3(25) => A(16), IN3(24) => A(15), IN3(23) => 
                           A(14), IN3(22) => A(13), IN3(21) => A(12), IN3(20) 
                           => A(11), IN3(19) => A(10), IN3(18) => A(9), IN3(17)
                           => A(8), IN3(16) => A(7), IN3(15) => A(6), IN3(14) 
                           => A(5), IN3(13) => A(4), IN3(12) => A(3), IN3(11) 
                           => A(2), IN3(10) => A(1), IN3(9) => A(0), IN3(8) => 
                           X_Logic0_port, IN3(7) => X_Logic0_port, IN3(6) => 
                           X_Logic0_port, IN3(5) => X_Logic0_port, IN3(4) => 
                           X_Logic0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(63) => negative_a_54_port, 
                           IN4(62) => negative_a_53_port, IN4(61) => 
                           negative_a_52_port, IN4(60) => negative_a_51_port, 
                           IN4(59) => negative_a_50_port, IN4(58) => 
                           negative_a_49_port, IN4(57) => negative_a_48_port, 
                           IN4(56) => negative_a_47_port, IN4(55) => 
                           negative_a_46_port, IN4(54) => negative_a_45_port, 
                           IN4(53) => negative_a_44_port, IN4(52) => 
                           negative_a_43_port, IN4(51) => negative_a_42_port, 
                           IN4(50) => negative_a_41_port, IN4(49) => 
                           negative_a_40_port, IN4(48) => negative_a_39_port, 
                           IN4(47) => negative_a_38_port, IN4(46) => 
                           negative_a_37_port, IN4(45) => negative_a_36_port, 
                           IN4(44) => negative_a_35_port, IN4(43) => 
                           negative_a_34_port, IN4(42) => n36, IN4(41) => n33, 
                           IN4(40) => negative_a_31_port, IN4(39) => 
                           negative_a_30_port, IN4(38) => negative_a_29_port, 
                           IN4(37) => negative_a_28_port, IN4(36) => 
                           negative_a_27_port, IN4(35) => negative_a_26_port, 
                           IN4(34) => negative_a_25_port, IN4(33) => 
                           negative_a_24_port, IN4(32) => negative_a_23_port, 
                           IN4(31) => negative_a_22_port, IN4(30) => 
                           negative_a_21_port, IN4(29) => negative_a_20_port, 
                           IN4(28) => negative_a_19_port, IN4(27) => 
                           negative_a_18_port, IN4(26) => negative_a_17_port, 
                           IN4(25) => negative_a_16_port, IN4(24) => 
                           negative_a_15_port, IN4(23) => negative_a_14_port, 
                           IN4(22) => negative_a_13_port, IN4(21) => 
                           negative_a_12_port, IN4(20) => negative_a_11_port, 
                           IN4(19) => negative_a_10_port, IN4(18) => 
                           negative_a_9_port, IN4(17) => negative_a_8_port, 
                           IN4(16) => negative_a_7_port, IN4(15) => 
                           negative_a_6_port, IN4(14) => negative_a_5_port, 
                           IN4(13) => negative_a_4_port, IN4(12) => 
                           negative_a_3_port, IN4(11) => negative_a_2_port, 
                           IN4(10) => negative_a_1_port, IN4(9) => 
                           negative_a_0_port, IN4(8) => X_Logic0_port, IN4(7) 
                           => X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) =>
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_4_2_port, S(1) => 
                           muxs_encoded_signals_4_1_port, S(0) => 
                           muxs_encoded_signals_4_0_port, O(63) => 
                           out_imux_4_63_port, O(62) => out_imux_4_62_port, 
                           O(61) => out_imux_4_61_port, O(60) => 
                           out_imux_4_60_port, O(59) => out_imux_4_59_port, 
                           O(58) => out_imux_4_58_port, O(57) => 
                           out_imux_4_57_port, O(56) => out_imux_4_56_port, 
                           O(55) => out_imux_4_55_port, O(54) => 
                           out_imux_4_54_port, O(53) => out_imux_4_53_port, 
                           O(52) => out_imux_4_52_port, O(51) => 
                           out_imux_4_51_port, O(50) => out_imux_4_50_port, 
                           O(49) => out_imux_4_49_port, O(48) => 
                           out_imux_4_48_port, O(47) => out_imux_4_47_port, 
                           O(46) => out_imux_4_46_port, O(45) => 
                           out_imux_4_45_port, O(44) => out_imux_4_44_port, 
                           O(43) => out_imux_4_43_port, O(42) => 
                           out_imux_4_42_port, O(41) => out_imux_4_41_port, 
                           O(40) => out_imux_4_40_port, O(39) => 
                           out_imux_4_39_port, O(38) => out_imux_4_38_port, 
                           O(37) => out_imux_4_37_port, O(36) => 
                           out_imux_4_36_port, O(35) => out_imux_4_35_port, 
                           O(34) => out_imux_4_34_port, O(33) => 
                           out_imux_4_33_port, O(32) => out_imux_4_32_port, 
                           O(31) => out_imux_4_31_port, O(30) => 
                           out_imux_4_30_port, O(29) => out_imux_4_29_port, 
                           O(28) => out_imux_4_28_port, O(27) => 
                           out_imux_4_27_port, O(26) => out_imux_4_26_port, 
                           O(25) => out_imux_4_25_port, O(24) => 
                           out_imux_4_24_port, O(23) => out_imux_4_23_port, 
                           O(22) => out_imux_4_22_port, O(21) => 
                           out_imux_4_21_port, O(20) => out_imux_4_20_port, 
                           O(19) => out_imux_4_19_port, O(18) => 
                           out_imux_4_18_port, O(17) => out_imux_4_17_port, 
                           O(16) => out_imux_4_16_port, O(15) => 
                           out_imux_4_15_port, O(14) => out_imux_4_14_port, 
                           O(13) => out_imux_4_13_port, O(12) => 
                           out_imux_4_12_port, O(11) => out_imux_4_11_port, 
                           O(10) => out_imux_4_10_port, O(9) => 
                           out_imux_4_9_port, O(8) => out_imux_4_8_port, O(7) 
                           => out_imux_4_7_port, O(6) => out_imux_4_6_port, 
                           O(5) => out_imux_4_5_port, O(4) => out_imux_4_4_port
                           , O(3) => out_imux_4_3_port, O(2) => 
                           out_imux_4_2_port, O(1) => out_imux_4_1_port, O(0) 
                           => out_imux_4_0_port);
   ADD64_i_4 : RCA_GENERIC_NBIT64_12 port map( A(63) => 
                           predigest_product_3_63_port, A(62) => 
                           predigest_product_3_62_port, A(61) => 
                           predigest_product_3_61_port, A(60) => 
                           predigest_product_3_60_port, A(59) => 
                           predigest_product_3_59_port, A(58) => 
                           predigest_product_3_58_port, A(57) => 
                           predigest_product_3_57_port, A(56) => 
                           predigest_product_3_56_port, A(55) => 
                           predigest_product_3_55_port, A(54) => 
                           predigest_product_3_54_port, A(53) => 
                           predigest_product_3_53_port, A(52) => 
                           predigest_product_3_52_port, A(51) => 
                           predigest_product_3_51_port, A(50) => 
                           predigest_product_3_50_port, A(49) => 
                           predigest_product_3_49_port, A(48) => 
                           predigest_product_3_48_port, A(47) => 
                           predigest_product_3_47_port, A(46) => 
                           predigest_product_3_46_port, A(45) => 
                           predigest_product_3_45_port, A(44) => 
                           predigest_product_3_44_port, A(43) => 
                           predigest_product_3_43_port, A(42) => 
                           predigest_product_3_42_port, A(41) => 
                           predigest_product_3_41_port, A(40) => 
                           predigest_product_3_40_port, A(39) => 
                           predigest_product_3_39_port, A(38) => 
                           predigest_product_3_38_port, A(37) => 
                           predigest_product_3_37_port, A(36) => 
                           predigest_product_3_36_port, A(35) => 
                           predigest_product_3_35_port, A(34) => 
                           predigest_product_3_34_port, A(33) => 
                           predigest_product_3_33_port, A(32) => 
                           predigest_product_3_32_port, A(31) => 
                           predigest_product_3_31_port, A(30) => 
                           predigest_product_3_30_port, A(29) => 
                           predigest_product_3_29_port, A(28) => 
                           predigest_product_3_28_port, A(27) => 
                           predigest_product_3_27_port, A(26) => 
                           predigest_product_3_26_port, A(25) => 
                           predigest_product_3_25_port, A(24) => 
                           predigest_product_3_24_port, A(23) => 
                           predigest_product_3_23_port, A(22) => 
                           predigest_product_3_22_port, A(21) => 
                           predigest_product_3_21_port, A(20) => 
                           predigest_product_3_20_port, A(19) => 
                           predigest_product_3_19_port, A(18) => 
                           predigest_product_3_18_port, A(17) => 
                           predigest_product_3_17_port, A(16) => 
                           predigest_product_3_16_port, A(15) => 
                           predigest_product_3_15_port, A(14) => 
                           predigest_product_3_14_port, A(13) => 
                           predigest_product_3_13_port, A(12) => 
                           predigest_product_3_12_port, A(11) => 
                           predigest_product_3_11_port, A(10) => 
                           predigest_product_3_10_port, A(9) => 
                           predigest_product_3_9_port, A(8) => 
                           predigest_product_3_8_port, A(7) => 
                           predigest_product_3_7_port, A(6) => 
                           predigest_product_3_6_port, A(5) => 
                           predigest_product_3_5_port, A(4) => 
                           predigest_product_3_4_port, A(3) => 
                           predigest_product_3_3_port, A(2) => 
                           predigest_product_3_2_port, A(1) => 
                           predigest_product_3_1_port, A(0) => 
                           predigest_product_3_0_port, B(63) => 
                           out_imux_4_63_port, B(62) => out_imux_4_62_port, 
                           B(61) => out_imux_4_61_port, B(60) => 
                           out_imux_4_60_port, B(59) => out_imux_4_59_port, 
                           B(58) => out_imux_4_58_port, B(57) => 
                           out_imux_4_57_port, B(56) => out_imux_4_56_port, 
                           B(55) => out_imux_4_55_port, B(54) => 
                           out_imux_4_54_port, B(53) => out_imux_4_53_port, 
                           B(52) => out_imux_4_52_port, B(51) => 
                           out_imux_4_51_port, B(50) => out_imux_4_50_port, 
                           B(49) => out_imux_4_49_port, B(48) => 
                           out_imux_4_48_port, B(47) => out_imux_4_47_port, 
                           B(46) => out_imux_4_46_port, B(45) => 
                           out_imux_4_45_port, B(44) => out_imux_4_44_port, 
                           B(43) => out_imux_4_43_port, B(42) => 
                           out_imux_4_42_port, B(41) => out_imux_4_41_port, 
                           B(40) => out_imux_4_40_port, B(39) => 
                           out_imux_4_39_port, B(38) => out_imux_4_38_port, 
                           B(37) => out_imux_4_37_port, B(36) => 
                           out_imux_4_36_port, B(35) => out_imux_4_35_port, 
                           B(34) => out_imux_4_34_port, B(33) => 
                           out_imux_4_33_port, B(32) => out_imux_4_32_port, 
                           B(31) => out_imux_4_31_port, B(30) => 
                           out_imux_4_30_port, B(29) => out_imux_4_29_port, 
                           B(28) => out_imux_4_28_port, B(27) => 
                           out_imux_4_27_port, B(26) => out_imux_4_26_port, 
                           B(25) => out_imux_4_25_port, B(24) => 
                           out_imux_4_24_port, B(23) => out_imux_4_23_port, 
                           B(22) => out_imux_4_22_port, B(21) => 
                           out_imux_4_21_port, B(20) => out_imux_4_20_port, 
                           B(19) => out_imux_4_19_port, B(18) => 
                           out_imux_4_18_port, B(17) => out_imux_4_17_port, 
                           B(16) => out_imux_4_16_port, B(15) => 
                           out_imux_4_15_port, B(14) => out_imux_4_14_port, 
                           B(13) => out_imux_4_13_port, B(12) => 
                           out_imux_4_12_port, B(11) => out_imux_4_11_port, 
                           B(10) => out_imux_4_10_port, B(9) => 
                           out_imux_4_9_port, B(8) => out_imux_4_8_port, B(7) 
                           => out_imux_4_7_port, B(6) => out_imux_4_6_port, 
                           B(5) => out_imux_4_5_port, B(4) => out_imux_4_4_port
                           , B(3) => out_imux_4_3_port, B(2) => 
                           out_imux_4_2_port, B(1) => out_imux_4_1_port, B(0) 
                           => out_imux_4_0_port, Ci => X_Logic0_port, S(63) => 
                           predigest_product_4_63_port, S(62) => 
                           predigest_product_4_62_port, S(61) => 
                           predigest_product_4_61_port, S(60) => 
                           predigest_product_4_60_port, S(59) => 
                           predigest_product_4_59_port, S(58) => 
                           predigest_product_4_58_port, S(57) => 
                           predigest_product_4_57_port, S(56) => 
                           predigest_product_4_56_port, S(55) => 
                           predigest_product_4_55_port, S(54) => 
                           predigest_product_4_54_port, S(53) => 
                           predigest_product_4_53_port, S(52) => 
                           predigest_product_4_52_port, S(51) => 
                           predigest_product_4_51_port, S(50) => 
                           predigest_product_4_50_port, S(49) => 
                           predigest_product_4_49_port, S(48) => 
                           predigest_product_4_48_port, S(47) => 
                           predigest_product_4_47_port, S(46) => 
                           predigest_product_4_46_port, S(45) => 
                           predigest_product_4_45_port, S(44) => 
                           predigest_product_4_44_port, S(43) => 
                           predigest_product_4_43_port, S(42) => 
                           predigest_product_4_42_port, S(41) => 
                           predigest_product_4_41_port, S(40) => 
                           predigest_product_4_40_port, S(39) => 
                           predigest_product_4_39_port, S(38) => 
                           predigest_product_4_38_port, S(37) => 
                           predigest_product_4_37_port, S(36) => 
                           predigest_product_4_36_port, S(35) => 
                           predigest_product_4_35_port, S(34) => 
                           predigest_product_4_34_port, S(33) => 
                           predigest_product_4_33_port, S(32) => 
                           predigest_product_4_32_port, S(31) => 
                           predigest_product_4_31_port, S(30) => 
                           predigest_product_4_30_port, S(29) => 
                           predigest_product_4_29_port, S(28) => 
                           predigest_product_4_28_port, S(27) => 
                           predigest_product_4_27_port, S(26) => 
                           predigest_product_4_26_port, S(25) => 
                           predigest_product_4_25_port, S(24) => 
                           predigest_product_4_24_port, S(23) => 
                           predigest_product_4_23_port, S(22) => 
                           predigest_product_4_22_port, S(21) => 
                           predigest_product_4_21_port, S(20) => 
                           predigest_product_4_20_port, S(19) => 
                           predigest_product_4_19_port, S(18) => 
                           predigest_product_4_18_port, S(17) => 
                           predigest_product_4_17_port, S(16) => 
                           predigest_product_4_16_port, S(15) => 
                           predigest_product_4_15_port, S(14) => 
                           predigest_product_4_14_port, S(13) => 
                           predigest_product_4_13_port, S(12) => 
                           predigest_product_4_12_port, S(11) => 
                           predigest_product_4_11_port, S(10) => 
                           predigest_product_4_10_port, S(9) => 
                           predigest_product_4_9_port, S(8) => 
                           predigest_product_4_8_port, S(7) => 
                           predigest_product_4_7_port, S(6) => 
                           predigest_product_4_6_port, S(5) => 
                           predigest_product_4_5_port, S(4) => 
                           predigest_product_4_4_port, S(3) => 
                           predigest_product_4_3_port, S(2) => 
                           predigest_product_4_2_port, S(1) => 
                           predigest_product_4_1_port, S(0) => 
                           predigest_product_4_0_port, Co => n_1095);
   ENC_i_5 : BOOTH_ENCODER_3BIT_15 port map( B(2) => B(11), B(1) => B(10), B(0)
                           => B(9), ENCODED(2) => muxs_encoded_signals_5_2_port
                           , ENCODED(1) => muxs_encoded_signals_5_1_port, 
                           ENCODED(0) => muxs_encoded_signals_5_0_port);
   MUX_i_5 : MUX51_GENERIC_NBIT64_11 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(31), IN1(51) 
                           => A(31), IN1(50) => A(31), IN1(49) => A(31), 
                           IN1(48) => A(31), IN1(47) => A(31), IN1(46) => A(31)
                           , IN1(45) => A(31), IN1(44) => A(31), IN1(43) => 
                           A(31), IN1(42) => A(31), IN1(41) => A(31), IN1(40) 
                           => A(30), IN1(39) => A(29), IN1(38) => A(28), 
                           IN1(37) => A(27), IN1(36) => A(26), IN1(35) => A(25)
                           , IN1(34) => A(24), IN1(33) => A(23), IN1(32) => 
                           A(22), IN1(31) => A(21), IN1(30) => A(20), IN1(29) 
                           => A(19), IN1(28) => A(18), IN1(27) => A(17), 
                           IN1(26) => A(16), IN1(25) => A(15), IN1(24) => A(14)
                           , IN1(23) => A(13), IN1(22) => A(12), IN1(21) => 
                           A(11), IN1(20) => A(10), IN1(19) => A(9), IN1(18) =>
                           A(8), IN1(17) => A(7), IN1(16) => A(6), IN1(15) => 
                           A(5), IN1(14) => A(4), IN1(13) => A(3), IN1(12) => 
                           A(2), IN1(11) => A(1), IN1(10) => A(0), IN1(9) => 
                           X_Logic0_port, IN1(8) => X_Logic0_port, IN1(7) => 
                           X_Logic0_port, IN1(6) => X_Logic0_port, IN1(5) => 
                           X_Logic0_port, IN1(4) => X_Logic0_port, IN1(3) => 
                           X_Logic0_port, IN1(2) => X_Logic0_port, IN1(1) => 
                           X_Logic0_port, IN1(0) => X_Logic0_port, IN2(63) => 
                           negative_a_53_port, IN2(62) => negative_a_52_port, 
                           IN2(61) => negative_a_51_port, IN2(60) => 
                           negative_a_50_port, IN2(59) => negative_a_49_port, 
                           IN2(58) => negative_a_48_port, IN2(57) => 
                           negative_a_47_port, IN2(56) => negative_a_46_port, 
                           IN2(55) => negative_a_45_port, IN2(54) => 
                           negative_a_44_port, IN2(53) => negative_a_43_port, 
                           IN2(52) => negative_a_42_port, IN2(51) => 
                           negative_a_41_port, IN2(50) => negative_a_40_port, 
                           IN2(49) => negative_a_39_port, IN2(48) => 
                           negative_a_38_port, IN2(47) => negative_a_37_port, 
                           IN2(46) => negative_a_36_port, IN2(45) => 
                           negative_a_35_port, IN2(44) => negative_a_34_port, 
                           IN2(43) => n36, IN2(42) => n33, IN2(41) => 
                           negative_a_31_port, IN2(40) => negative_a_30_port, 
                           IN2(39) => negative_a_29_port, IN2(38) => 
                           negative_a_28_port, IN2(37) => negative_a_27_port, 
                           IN2(36) => negative_a_26_port, IN2(35) => 
                           negative_a_25_port, IN2(34) => negative_a_24_port, 
                           IN2(33) => negative_a_23_port, IN2(32) => 
                           negative_a_22_port, IN2(31) => negative_a_21_port, 
                           IN2(30) => negative_a_20_port, IN2(29) => 
                           negative_a_19_port, IN2(28) => negative_a_18_port, 
                           IN2(27) => negative_a_17_port, IN2(26) => 
                           negative_a_16_port, IN2(25) => negative_a_15_port, 
                           IN2(24) => negative_a_14_port, IN2(23) => 
                           negative_a_13_port, IN2(22) => negative_a_12_port, 
                           IN2(21) => negative_a_11_port, IN2(20) => 
                           negative_a_10_port, IN2(19) => negative_a_9_port, 
                           IN2(18) => negative_a_8_port, IN2(17) => 
                           negative_a_7_port, IN2(16) => negative_a_6_port, 
                           IN2(15) => negative_a_5_port, IN2(14) => 
                           negative_a_4_port, IN2(13) => negative_a_3_port, 
                           IN2(12) => negative_a_2_port, IN2(11) => 
                           negative_a_1_port, IN2(10) => negative_a_0_port, 
                           IN2(9) => X_Logic0_port, IN2(8) => X_Logic0_port, 
                           IN2(7) => X_Logic0_port, IN2(6) => X_Logic0_port, 
                           IN2(5) => X_Logic0_port, IN2(4) => X_Logic0_port, 
                           IN2(3) => X_Logic0_port, IN2(2) => X_Logic0_port, 
                           IN2(1) => X_Logic0_port, IN2(0) => X_Logic0_port, 
                           IN3(63) => A(31), IN3(62) => A(31), IN3(61) => A(31)
                           , IN3(60) => A(31), IN3(59) => A(31), IN3(58) => 
                           A(31), IN3(57) => A(31), IN3(56) => A(31), IN3(55) 
                           => A(31), IN3(54) => A(31), IN3(53) => A(31), 
                           IN3(52) => A(31), IN3(51) => A(31), IN3(50) => A(31)
                           , IN3(49) => A(31), IN3(48) => A(31), IN3(47) => 
                           A(31), IN3(46) => A(31), IN3(45) => A(31), IN3(44) 
                           => A(31), IN3(43) => A(31), IN3(42) => A(31), 
                           IN3(41) => A(30), IN3(40) => A(29), IN3(39) => A(28)
                           , IN3(38) => A(27), IN3(37) => A(26), IN3(36) => 
                           A(25), IN3(35) => A(24), IN3(34) => A(23), IN3(33) 
                           => A(22), IN3(32) => A(21), IN3(31) => A(20), 
                           IN3(30) => A(19), IN3(29) => A(18), IN3(28) => A(17)
                           , IN3(27) => A(16), IN3(26) => A(15), IN3(25) => 
                           A(14), IN3(24) => A(13), IN3(23) => A(12), IN3(22) 
                           => A(11), IN3(21) => A(10), IN3(20) => A(9), IN3(19)
                           => A(8), IN3(18) => A(7), IN3(17) => A(6), IN3(16) 
                           => A(5), IN3(15) => A(4), IN3(14) => A(3), IN3(13) 
                           => A(2), IN3(12) => A(1), IN3(11) => A(0), IN3(10) 
                           => X_Logic0_port, IN3(9) => X_Logic0_port, IN3(8) =>
                           X_Logic0_port, IN3(7) => X_Logic0_port, IN3(6) => 
                           X_Logic0_port, IN3(5) => X_Logic0_port, IN3(4) => 
                           X_Logic0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(63) => negative_a_52_port, 
                           IN4(62) => negative_a_51_port, IN4(61) => 
                           negative_a_50_port, IN4(60) => negative_a_49_port, 
                           IN4(59) => negative_a_48_port, IN4(58) => 
                           negative_a_47_port, IN4(57) => negative_a_46_port, 
                           IN4(56) => negative_a_45_port, IN4(55) => 
                           negative_a_44_port, IN4(54) => negative_a_43_port, 
                           IN4(53) => negative_a_42_port, IN4(52) => 
                           negative_a_41_port, IN4(51) => negative_a_40_port, 
                           IN4(50) => negative_a_39_port, IN4(49) => 
                           negative_a_38_port, IN4(48) => negative_a_37_port, 
                           IN4(47) => negative_a_36_port, IN4(46) => 
                           negative_a_35_port, IN4(45) => negative_a_34_port, 
                           IN4(44) => n36, IN4(43) => n33, IN4(42) => 
                           negative_a_31_port, IN4(41) => negative_a_30_port, 
                           IN4(40) => negative_a_29_port, IN4(39) => 
                           negative_a_28_port, IN4(38) => negative_a_27_port, 
                           IN4(37) => negative_a_26_port, IN4(36) => 
                           negative_a_25_port, IN4(35) => negative_a_24_port, 
                           IN4(34) => negative_a_23_port, IN4(33) => 
                           negative_a_22_port, IN4(32) => negative_a_21_port, 
                           IN4(31) => negative_a_20_port, IN4(30) => 
                           negative_a_19_port, IN4(29) => negative_a_18_port, 
                           IN4(28) => negative_a_17_port, IN4(27) => 
                           negative_a_16_port, IN4(26) => negative_a_15_port, 
                           IN4(25) => negative_a_14_port, IN4(24) => 
                           negative_a_13_port, IN4(23) => negative_a_12_port, 
                           IN4(22) => negative_a_11_port, IN4(21) => 
                           negative_a_10_port, IN4(20) => negative_a_9_port, 
                           IN4(19) => negative_a_8_port, IN4(18) => 
                           negative_a_7_port, IN4(17) => negative_a_6_port, 
                           IN4(16) => negative_a_5_port, IN4(15) => 
                           negative_a_4_port, IN4(14) => negative_a_3_port, 
                           IN4(13) => negative_a_2_port, IN4(12) => 
                           negative_a_1_port, IN4(11) => negative_a_0_port, 
                           IN4(10) => X_Logic0_port, IN4(9) => X_Logic0_port, 
                           IN4(8) => X_Logic0_port, IN4(7) => X_Logic0_port, 
                           IN4(6) => X_Logic0_port, IN4(5) => X_Logic0_port, 
                           IN4(4) => X_Logic0_port, IN4(3) => X_Logic0_port, 
                           IN4(2) => X_Logic0_port, IN4(1) => X_Logic0_port, 
                           IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_5_2_port, S(1) => 
                           muxs_encoded_signals_5_1_port, S(0) => 
                           muxs_encoded_signals_5_0_port, O(63) => 
                           out_imux_5_63_port, O(62) => out_imux_5_62_port, 
                           O(61) => out_imux_5_61_port, O(60) => 
                           out_imux_5_60_port, O(59) => out_imux_5_59_port, 
                           O(58) => out_imux_5_58_port, O(57) => 
                           out_imux_5_57_port, O(56) => out_imux_5_56_port, 
                           O(55) => out_imux_5_55_port, O(54) => 
                           out_imux_5_54_port, O(53) => out_imux_5_53_port, 
                           O(52) => out_imux_5_52_port, O(51) => 
                           out_imux_5_51_port, O(50) => out_imux_5_50_port, 
                           O(49) => out_imux_5_49_port, O(48) => 
                           out_imux_5_48_port, O(47) => out_imux_5_47_port, 
                           O(46) => out_imux_5_46_port, O(45) => 
                           out_imux_5_45_port, O(44) => out_imux_5_44_port, 
                           O(43) => out_imux_5_43_port, O(42) => 
                           out_imux_5_42_port, O(41) => out_imux_5_41_port, 
                           O(40) => out_imux_5_40_port, O(39) => 
                           out_imux_5_39_port, O(38) => out_imux_5_38_port, 
                           O(37) => out_imux_5_37_port, O(36) => 
                           out_imux_5_36_port, O(35) => out_imux_5_35_port, 
                           O(34) => out_imux_5_34_port, O(33) => 
                           out_imux_5_33_port, O(32) => out_imux_5_32_port, 
                           O(31) => out_imux_5_31_port, O(30) => 
                           out_imux_5_30_port, O(29) => out_imux_5_29_port, 
                           O(28) => out_imux_5_28_port, O(27) => 
                           out_imux_5_27_port, O(26) => out_imux_5_26_port, 
                           O(25) => out_imux_5_25_port, O(24) => 
                           out_imux_5_24_port, O(23) => out_imux_5_23_port, 
                           O(22) => out_imux_5_22_port, O(21) => 
                           out_imux_5_21_port, O(20) => out_imux_5_20_port, 
                           O(19) => out_imux_5_19_port, O(18) => 
                           out_imux_5_18_port, O(17) => out_imux_5_17_port, 
                           O(16) => out_imux_5_16_port, O(15) => 
                           out_imux_5_15_port, O(14) => out_imux_5_14_port, 
                           O(13) => out_imux_5_13_port, O(12) => 
                           out_imux_5_12_port, O(11) => out_imux_5_11_port, 
                           O(10) => out_imux_5_10_port, O(9) => 
                           out_imux_5_9_port, O(8) => out_imux_5_8_port, O(7) 
                           => out_imux_5_7_port, O(6) => out_imux_5_6_port, 
                           O(5) => out_imux_5_5_port, O(4) => out_imux_5_4_port
                           , O(3) => out_imux_5_3_port, O(2) => 
                           out_imux_5_2_port, O(1) => out_imux_5_1_port, O(0) 
                           => out_imux_5_0_port);
   ADD64_i_5 : RCA_GENERIC_NBIT64_11 port map( A(63) => 
                           predigest_product_4_63_port, A(62) => 
                           predigest_product_4_62_port, A(61) => 
                           predigest_product_4_61_port, A(60) => 
                           predigest_product_4_60_port, A(59) => 
                           predigest_product_4_59_port, A(58) => 
                           predigest_product_4_58_port, A(57) => 
                           predigest_product_4_57_port, A(56) => 
                           predigest_product_4_56_port, A(55) => 
                           predigest_product_4_55_port, A(54) => 
                           predigest_product_4_54_port, A(53) => 
                           predigest_product_4_53_port, A(52) => 
                           predigest_product_4_52_port, A(51) => 
                           predigest_product_4_51_port, A(50) => 
                           predigest_product_4_50_port, A(49) => 
                           predigest_product_4_49_port, A(48) => 
                           predigest_product_4_48_port, A(47) => 
                           predigest_product_4_47_port, A(46) => 
                           predigest_product_4_46_port, A(45) => 
                           predigest_product_4_45_port, A(44) => 
                           predigest_product_4_44_port, A(43) => 
                           predigest_product_4_43_port, A(42) => 
                           predigest_product_4_42_port, A(41) => 
                           predigest_product_4_41_port, A(40) => 
                           predigest_product_4_40_port, A(39) => 
                           predigest_product_4_39_port, A(38) => 
                           predigest_product_4_38_port, A(37) => 
                           predigest_product_4_37_port, A(36) => 
                           predigest_product_4_36_port, A(35) => 
                           predigest_product_4_35_port, A(34) => 
                           predigest_product_4_34_port, A(33) => 
                           predigest_product_4_33_port, A(32) => 
                           predigest_product_4_32_port, A(31) => 
                           predigest_product_4_31_port, A(30) => 
                           predigest_product_4_30_port, A(29) => 
                           predigest_product_4_29_port, A(28) => 
                           predigest_product_4_28_port, A(27) => 
                           predigest_product_4_27_port, A(26) => 
                           predigest_product_4_26_port, A(25) => 
                           predigest_product_4_25_port, A(24) => 
                           predigest_product_4_24_port, A(23) => 
                           predigest_product_4_23_port, A(22) => 
                           predigest_product_4_22_port, A(21) => 
                           predigest_product_4_21_port, A(20) => 
                           predigest_product_4_20_port, A(19) => 
                           predigest_product_4_19_port, A(18) => 
                           predigest_product_4_18_port, A(17) => 
                           predigest_product_4_17_port, A(16) => 
                           predigest_product_4_16_port, A(15) => 
                           predigest_product_4_15_port, A(14) => 
                           predigest_product_4_14_port, A(13) => 
                           predigest_product_4_13_port, A(12) => 
                           predigest_product_4_12_port, A(11) => 
                           predigest_product_4_11_port, A(10) => 
                           predigest_product_4_10_port, A(9) => 
                           predigest_product_4_9_port, A(8) => 
                           predigest_product_4_8_port, A(7) => 
                           predigest_product_4_7_port, A(6) => 
                           predigest_product_4_6_port, A(5) => 
                           predigest_product_4_5_port, A(4) => 
                           predigest_product_4_4_port, A(3) => 
                           predigest_product_4_3_port, A(2) => 
                           predigest_product_4_2_port, A(1) => 
                           predigest_product_4_1_port, A(0) => 
                           predigest_product_4_0_port, B(63) => 
                           out_imux_5_63_port, B(62) => out_imux_5_62_port, 
                           B(61) => out_imux_5_61_port, B(60) => 
                           out_imux_5_60_port, B(59) => out_imux_5_59_port, 
                           B(58) => out_imux_5_58_port, B(57) => 
                           out_imux_5_57_port, B(56) => out_imux_5_56_port, 
                           B(55) => out_imux_5_55_port, B(54) => 
                           out_imux_5_54_port, B(53) => out_imux_5_53_port, 
                           B(52) => out_imux_5_52_port, B(51) => 
                           out_imux_5_51_port, B(50) => out_imux_5_50_port, 
                           B(49) => out_imux_5_49_port, B(48) => 
                           out_imux_5_48_port, B(47) => out_imux_5_47_port, 
                           B(46) => out_imux_5_46_port, B(45) => 
                           out_imux_5_45_port, B(44) => out_imux_5_44_port, 
                           B(43) => out_imux_5_43_port, B(42) => 
                           out_imux_5_42_port, B(41) => out_imux_5_41_port, 
                           B(40) => out_imux_5_40_port, B(39) => 
                           out_imux_5_39_port, B(38) => out_imux_5_38_port, 
                           B(37) => out_imux_5_37_port, B(36) => 
                           out_imux_5_36_port, B(35) => out_imux_5_35_port, 
                           B(34) => out_imux_5_34_port, B(33) => 
                           out_imux_5_33_port, B(32) => out_imux_5_32_port, 
                           B(31) => out_imux_5_31_port, B(30) => 
                           out_imux_5_30_port, B(29) => out_imux_5_29_port, 
                           B(28) => out_imux_5_28_port, B(27) => 
                           out_imux_5_27_port, B(26) => out_imux_5_26_port, 
                           B(25) => out_imux_5_25_port, B(24) => 
                           out_imux_5_24_port, B(23) => out_imux_5_23_port, 
                           B(22) => out_imux_5_22_port, B(21) => 
                           out_imux_5_21_port, B(20) => out_imux_5_20_port, 
                           B(19) => out_imux_5_19_port, B(18) => 
                           out_imux_5_18_port, B(17) => out_imux_5_17_port, 
                           B(16) => out_imux_5_16_port, B(15) => 
                           out_imux_5_15_port, B(14) => out_imux_5_14_port, 
                           B(13) => out_imux_5_13_port, B(12) => 
                           out_imux_5_12_port, B(11) => out_imux_5_11_port, 
                           B(10) => out_imux_5_10_port, B(9) => 
                           out_imux_5_9_port, B(8) => out_imux_5_8_port, B(7) 
                           => out_imux_5_7_port, B(6) => out_imux_5_6_port, 
                           B(5) => out_imux_5_5_port, B(4) => out_imux_5_4_port
                           , B(3) => out_imux_5_3_port, B(2) => 
                           out_imux_5_2_port, B(1) => out_imux_5_1_port, B(0) 
                           => out_imux_5_0_port, Ci => X_Logic0_port, S(63) => 
                           predigest_product_5_63_port, S(62) => 
                           predigest_product_5_62_port, S(61) => 
                           predigest_product_5_61_port, S(60) => 
                           predigest_product_5_60_port, S(59) => 
                           predigest_product_5_59_port, S(58) => 
                           predigest_product_5_58_port, S(57) => 
                           predigest_product_5_57_port, S(56) => 
                           predigest_product_5_56_port, S(55) => 
                           predigest_product_5_55_port, S(54) => 
                           predigest_product_5_54_port, S(53) => 
                           predigest_product_5_53_port, S(52) => 
                           predigest_product_5_52_port, S(51) => 
                           predigest_product_5_51_port, S(50) => 
                           predigest_product_5_50_port, S(49) => 
                           predigest_product_5_49_port, S(48) => 
                           predigest_product_5_48_port, S(47) => 
                           predigest_product_5_47_port, S(46) => 
                           predigest_product_5_46_port, S(45) => 
                           predigest_product_5_45_port, S(44) => 
                           predigest_product_5_44_port, S(43) => 
                           predigest_product_5_43_port, S(42) => 
                           predigest_product_5_42_port, S(41) => 
                           predigest_product_5_41_port, S(40) => 
                           predigest_product_5_40_port, S(39) => 
                           predigest_product_5_39_port, S(38) => 
                           predigest_product_5_38_port, S(37) => 
                           predigest_product_5_37_port, S(36) => 
                           predigest_product_5_36_port, S(35) => 
                           predigest_product_5_35_port, S(34) => 
                           predigest_product_5_34_port, S(33) => 
                           predigest_product_5_33_port, S(32) => 
                           predigest_product_5_32_port, S(31) => 
                           predigest_product_5_31_port, S(30) => 
                           predigest_product_5_30_port, S(29) => 
                           predigest_product_5_29_port, S(28) => 
                           predigest_product_5_28_port, S(27) => 
                           predigest_product_5_27_port, S(26) => 
                           predigest_product_5_26_port, S(25) => 
                           predigest_product_5_25_port, S(24) => 
                           predigest_product_5_24_port, S(23) => 
                           predigest_product_5_23_port, S(22) => 
                           predigest_product_5_22_port, S(21) => 
                           predigest_product_5_21_port, S(20) => 
                           predigest_product_5_20_port, S(19) => 
                           predigest_product_5_19_port, S(18) => 
                           predigest_product_5_18_port, S(17) => 
                           predigest_product_5_17_port, S(16) => 
                           predigest_product_5_16_port, S(15) => 
                           predigest_product_5_15_port, S(14) => 
                           predigest_product_5_14_port, S(13) => 
                           predigest_product_5_13_port, S(12) => 
                           predigest_product_5_12_port, S(11) => 
                           predigest_product_5_11_port, S(10) => 
                           predigest_product_5_10_port, S(9) => 
                           predigest_product_5_9_port, S(8) => 
                           predigest_product_5_8_port, S(7) => 
                           predigest_product_5_7_port, S(6) => 
                           predigest_product_5_6_port, S(5) => 
                           predigest_product_5_5_port, S(4) => 
                           predigest_product_5_4_port, S(3) => 
                           predigest_product_5_3_port, S(2) => 
                           predigest_product_5_2_port, S(1) => 
                           predigest_product_5_1_port, S(0) => 
                           predigest_product_5_0_port, Co => n_1096);
   ENC_i_6 : BOOTH_ENCODER_3BIT_14 port map( B(2) => B(13), B(1) => B(12), B(0)
                           => B(11), ENCODED(2) => 
                           muxs_encoded_signals_6_2_port, ENCODED(1) => 
                           muxs_encoded_signals_6_1_port, ENCODED(0) => 
                           muxs_encoded_signals_6_0_port);
   MUX_i_6 : MUX51_GENERIC_NBIT64_10 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(31), IN1(51) 
                           => A(31), IN1(50) => A(31), IN1(49) => A(31), 
                           IN1(48) => A(31), IN1(47) => A(31), IN1(46) => A(31)
                           , IN1(45) => A(31), IN1(44) => A(31), IN1(43) => 
                           A(31), IN1(42) => A(30), IN1(41) => A(29), IN1(40) 
                           => A(28), IN1(39) => A(27), IN1(38) => A(26), 
                           IN1(37) => A(25), IN1(36) => A(24), IN1(35) => A(23)
                           , IN1(34) => A(22), IN1(33) => A(21), IN1(32) => 
                           A(20), IN1(31) => A(19), IN1(30) => A(18), IN1(29) 
                           => A(17), IN1(28) => A(16), IN1(27) => A(15), 
                           IN1(26) => A(14), IN1(25) => A(13), IN1(24) => A(12)
                           , IN1(23) => A(11), IN1(22) => A(10), IN1(21) => 
                           A(9), IN1(20) => A(8), IN1(19) => A(7), IN1(18) => 
                           A(6), IN1(17) => A(5), IN1(16) => A(4), IN1(15) => 
                           A(3), IN1(14) => A(2), IN1(13) => A(1), IN1(12) => 
                           A(0), IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(63) => negative_a_51_port, 
                           IN2(62) => negative_a_50_port, IN2(61) => 
                           negative_a_49_port, IN2(60) => negative_a_48_port, 
                           IN2(59) => negative_a_47_port, IN2(58) => 
                           negative_a_46_port, IN2(57) => negative_a_45_port, 
                           IN2(56) => negative_a_44_port, IN2(55) => 
                           negative_a_43_port, IN2(54) => negative_a_42_port, 
                           IN2(53) => negative_a_41_port, IN2(52) => 
                           negative_a_40_port, IN2(51) => negative_a_39_port, 
                           IN2(50) => negative_a_38_port, IN2(49) => 
                           negative_a_37_port, IN2(48) => negative_a_36_port, 
                           IN2(47) => negative_a_35_port, IN2(46) => 
                           negative_a_34_port, IN2(45) => n37, IN2(44) => n34, 
                           IN2(43) => negative_a_31_port, IN2(42) => 
                           negative_a_30_port, IN2(41) => negative_a_29_port, 
                           IN2(40) => negative_a_28_port, IN2(39) => 
                           negative_a_27_port, IN2(38) => negative_a_26_port, 
                           IN2(37) => negative_a_25_port, IN2(36) => 
                           negative_a_24_port, IN2(35) => negative_a_23_port, 
                           IN2(34) => negative_a_22_port, IN2(33) => 
                           negative_a_21_port, IN2(32) => negative_a_20_port, 
                           IN2(31) => negative_a_19_port, IN2(30) => 
                           negative_a_18_port, IN2(29) => negative_a_17_port, 
                           IN2(28) => negative_a_16_port, IN2(27) => 
                           negative_a_15_port, IN2(26) => negative_a_14_port, 
                           IN2(25) => negative_a_13_port, IN2(24) => 
                           negative_a_12_port, IN2(23) => negative_a_11_port, 
                           IN2(22) => negative_a_10_port, IN2(21) => 
                           negative_a_9_port, IN2(20) => negative_a_8_port, 
                           IN2(19) => negative_a_7_port, IN2(18) => 
                           negative_a_6_port, IN2(17) => negative_a_5_port, 
                           IN2(16) => negative_a_4_port, IN2(15) => 
                           negative_a_3_port, IN2(14) => negative_a_2_port, 
                           IN2(13) => negative_a_1_port, IN2(12) => 
                           negative_a_0_port, IN2(11) => X_Logic0_port, IN2(10)
                           => X_Logic0_port, IN2(9) => X_Logic0_port, IN2(8) =>
                           X_Logic0_port, IN2(7) => X_Logic0_port, IN2(6) => 
                           X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) => 
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(63) => A(31), IN3(62) => A(31), 
                           IN3(61) => A(31), IN3(60) => A(31), IN3(59) => A(31)
                           , IN3(58) => A(31), IN3(57) => A(31), IN3(56) => 
                           A(31), IN3(55) => A(31), IN3(54) => A(31), IN3(53) 
                           => A(31), IN3(52) => A(31), IN3(51) => A(31), 
                           IN3(50) => A(31), IN3(49) => A(31), IN3(48) => A(31)
                           , IN3(47) => A(31), IN3(46) => A(31), IN3(45) => 
                           A(31), IN3(44) => A(31), IN3(43) => A(30), IN3(42) 
                           => A(29), IN3(41) => A(28), IN3(40) => A(27), 
                           IN3(39) => A(26), IN3(38) => A(25), IN3(37) => A(24)
                           , IN3(36) => A(23), IN3(35) => A(22), IN3(34) => 
                           A(21), IN3(33) => A(20), IN3(32) => A(19), IN3(31) 
                           => A(18), IN3(30) => A(17), IN3(29) => A(16), 
                           IN3(28) => A(15), IN3(27) => A(14), IN3(26) => A(13)
                           , IN3(25) => A(12), IN3(24) => A(11), IN3(23) => 
                           A(10), IN3(22) => A(9), IN3(21) => A(8), IN3(20) => 
                           A(7), IN3(19) => A(6), IN3(18) => A(5), IN3(17) => 
                           A(4), IN3(16) => A(3), IN3(15) => A(2), IN3(14) => 
                           A(1), IN3(13) => A(0), IN3(12) => X_Logic0_port, 
                           IN3(11) => X_Logic0_port, IN3(10) => X_Logic0_port, 
                           IN3(9) => X_Logic0_port, IN3(8) => X_Logic0_port, 
                           IN3(7) => X_Logic0_port, IN3(6) => X_Logic0_port, 
                           IN3(5) => X_Logic0_port, IN3(4) => X_Logic0_port, 
                           IN3(3) => X_Logic0_port, IN3(2) => X_Logic0_port, 
                           IN3(1) => X_Logic0_port, IN3(0) => X_Logic0_port, 
                           IN4(63) => negative_a_50_port, IN4(62) => 
                           negative_a_49_port, IN4(61) => negative_a_48_port, 
                           IN4(60) => negative_a_47_port, IN4(59) => 
                           negative_a_46_port, IN4(58) => negative_a_45_port, 
                           IN4(57) => negative_a_44_port, IN4(56) => 
                           negative_a_43_port, IN4(55) => negative_a_42_port, 
                           IN4(54) => negative_a_41_port, IN4(53) => 
                           negative_a_40_port, IN4(52) => negative_a_39_port, 
                           IN4(51) => negative_a_38_port, IN4(50) => 
                           negative_a_37_port, IN4(49) => negative_a_36_port, 
                           IN4(48) => negative_a_35_port, IN4(47) => 
                           negative_a_34_port, IN4(46) => n36, IN4(45) => n33, 
                           IN4(44) => negative_a_31_port, IN4(43) => 
                           negative_a_30_port, IN4(42) => negative_a_29_port, 
                           IN4(41) => negative_a_28_port, IN4(40) => 
                           negative_a_27_port, IN4(39) => negative_a_26_port, 
                           IN4(38) => negative_a_25_port, IN4(37) => 
                           negative_a_24_port, IN4(36) => negative_a_23_port, 
                           IN4(35) => negative_a_22_port, IN4(34) => 
                           negative_a_21_port, IN4(33) => negative_a_20_port, 
                           IN4(32) => negative_a_19_port, IN4(31) => 
                           negative_a_18_port, IN4(30) => negative_a_17_port, 
                           IN4(29) => negative_a_16_port, IN4(28) => 
                           negative_a_15_port, IN4(27) => negative_a_14_port, 
                           IN4(26) => negative_a_13_port, IN4(25) => 
                           negative_a_12_port, IN4(24) => negative_a_11_port, 
                           IN4(23) => negative_a_10_port, IN4(22) => 
                           negative_a_9_port, IN4(21) => negative_a_8_port, 
                           IN4(20) => negative_a_7_port, IN4(19) => 
                           negative_a_6_port, IN4(18) => negative_a_5_port, 
                           IN4(17) => negative_a_4_port, IN4(16) => 
                           negative_a_3_port, IN4(15) => negative_a_2_port, 
                           IN4(14) => negative_a_1_port, IN4(13) => 
                           negative_a_0_port, IN4(12) => X_Logic0_port, IN4(11)
                           => X_Logic0_port, IN4(10) => X_Logic0_port, IN4(9) 
                           => X_Logic0_port, IN4(8) => X_Logic0_port, IN4(7) =>
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_6_2_port, S(1) => 
                           muxs_encoded_signals_6_1_port, S(0) => 
                           muxs_encoded_signals_6_0_port, O(63) => 
                           out_imux_6_63_port, O(62) => out_imux_6_62_port, 
                           O(61) => out_imux_6_61_port, O(60) => 
                           out_imux_6_60_port, O(59) => out_imux_6_59_port, 
                           O(58) => out_imux_6_58_port, O(57) => 
                           out_imux_6_57_port, O(56) => out_imux_6_56_port, 
                           O(55) => out_imux_6_55_port, O(54) => 
                           out_imux_6_54_port, O(53) => out_imux_6_53_port, 
                           O(52) => out_imux_6_52_port, O(51) => 
                           out_imux_6_51_port, O(50) => out_imux_6_50_port, 
                           O(49) => out_imux_6_49_port, O(48) => 
                           out_imux_6_48_port, O(47) => out_imux_6_47_port, 
                           O(46) => out_imux_6_46_port, O(45) => 
                           out_imux_6_45_port, O(44) => out_imux_6_44_port, 
                           O(43) => out_imux_6_43_port, O(42) => 
                           out_imux_6_42_port, O(41) => out_imux_6_41_port, 
                           O(40) => out_imux_6_40_port, O(39) => 
                           out_imux_6_39_port, O(38) => out_imux_6_38_port, 
                           O(37) => out_imux_6_37_port, O(36) => 
                           out_imux_6_36_port, O(35) => out_imux_6_35_port, 
                           O(34) => out_imux_6_34_port, O(33) => 
                           out_imux_6_33_port, O(32) => out_imux_6_32_port, 
                           O(31) => out_imux_6_31_port, O(30) => 
                           out_imux_6_30_port, O(29) => out_imux_6_29_port, 
                           O(28) => out_imux_6_28_port, O(27) => 
                           out_imux_6_27_port, O(26) => out_imux_6_26_port, 
                           O(25) => out_imux_6_25_port, O(24) => 
                           out_imux_6_24_port, O(23) => out_imux_6_23_port, 
                           O(22) => out_imux_6_22_port, O(21) => 
                           out_imux_6_21_port, O(20) => out_imux_6_20_port, 
                           O(19) => out_imux_6_19_port, O(18) => 
                           out_imux_6_18_port, O(17) => out_imux_6_17_port, 
                           O(16) => out_imux_6_16_port, O(15) => 
                           out_imux_6_15_port, O(14) => out_imux_6_14_port, 
                           O(13) => out_imux_6_13_port, O(12) => 
                           out_imux_6_12_port, O(11) => out_imux_6_11_port, 
                           O(10) => out_imux_6_10_port, O(9) => 
                           out_imux_6_9_port, O(8) => out_imux_6_8_port, O(7) 
                           => out_imux_6_7_port, O(6) => out_imux_6_6_port, 
                           O(5) => out_imux_6_5_port, O(4) => out_imux_6_4_port
                           , O(3) => out_imux_6_3_port, O(2) => 
                           out_imux_6_2_port, O(1) => out_imux_6_1_port, O(0) 
                           => out_imux_6_0_port);
   ADD64_i_6 : RCA_GENERIC_NBIT64_10 port map( A(63) => 
                           predigest_product_5_63_port, A(62) => 
                           predigest_product_5_62_port, A(61) => 
                           predigest_product_5_61_port, A(60) => 
                           predigest_product_5_60_port, A(59) => 
                           predigest_product_5_59_port, A(58) => 
                           predigest_product_5_58_port, A(57) => 
                           predigest_product_5_57_port, A(56) => 
                           predigest_product_5_56_port, A(55) => 
                           predigest_product_5_55_port, A(54) => 
                           predigest_product_5_54_port, A(53) => 
                           predigest_product_5_53_port, A(52) => 
                           predigest_product_5_52_port, A(51) => 
                           predigest_product_5_51_port, A(50) => 
                           predigest_product_5_50_port, A(49) => 
                           predigest_product_5_49_port, A(48) => 
                           predigest_product_5_48_port, A(47) => 
                           predigest_product_5_47_port, A(46) => 
                           predigest_product_5_46_port, A(45) => 
                           predigest_product_5_45_port, A(44) => 
                           predigest_product_5_44_port, A(43) => 
                           predigest_product_5_43_port, A(42) => 
                           predigest_product_5_42_port, A(41) => 
                           predigest_product_5_41_port, A(40) => 
                           predigest_product_5_40_port, A(39) => 
                           predigest_product_5_39_port, A(38) => 
                           predigest_product_5_38_port, A(37) => 
                           predigest_product_5_37_port, A(36) => 
                           predigest_product_5_36_port, A(35) => 
                           predigest_product_5_35_port, A(34) => 
                           predigest_product_5_34_port, A(33) => 
                           predigest_product_5_33_port, A(32) => 
                           predigest_product_5_32_port, A(31) => 
                           predigest_product_5_31_port, A(30) => 
                           predigest_product_5_30_port, A(29) => 
                           predigest_product_5_29_port, A(28) => 
                           predigest_product_5_28_port, A(27) => 
                           predigest_product_5_27_port, A(26) => 
                           predigest_product_5_26_port, A(25) => 
                           predigest_product_5_25_port, A(24) => 
                           predigest_product_5_24_port, A(23) => 
                           predigest_product_5_23_port, A(22) => 
                           predigest_product_5_22_port, A(21) => 
                           predigest_product_5_21_port, A(20) => 
                           predigest_product_5_20_port, A(19) => 
                           predigest_product_5_19_port, A(18) => 
                           predigest_product_5_18_port, A(17) => 
                           predigest_product_5_17_port, A(16) => 
                           predigest_product_5_16_port, A(15) => 
                           predigest_product_5_15_port, A(14) => 
                           predigest_product_5_14_port, A(13) => 
                           predigest_product_5_13_port, A(12) => 
                           predigest_product_5_12_port, A(11) => 
                           predigest_product_5_11_port, A(10) => 
                           predigest_product_5_10_port, A(9) => 
                           predigest_product_5_9_port, A(8) => 
                           predigest_product_5_8_port, A(7) => 
                           predigest_product_5_7_port, A(6) => 
                           predigest_product_5_6_port, A(5) => 
                           predigest_product_5_5_port, A(4) => 
                           predigest_product_5_4_port, A(3) => 
                           predigest_product_5_3_port, A(2) => 
                           predigest_product_5_2_port, A(1) => 
                           predigest_product_5_1_port, A(0) => 
                           predigest_product_5_0_port, B(63) => 
                           out_imux_6_63_port, B(62) => out_imux_6_62_port, 
                           B(61) => out_imux_6_61_port, B(60) => 
                           out_imux_6_60_port, B(59) => out_imux_6_59_port, 
                           B(58) => out_imux_6_58_port, B(57) => 
                           out_imux_6_57_port, B(56) => out_imux_6_56_port, 
                           B(55) => out_imux_6_55_port, B(54) => 
                           out_imux_6_54_port, B(53) => out_imux_6_53_port, 
                           B(52) => out_imux_6_52_port, B(51) => 
                           out_imux_6_51_port, B(50) => out_imux_6_50_port, 
                           B(49) => out_imux_6_49_port, B(48) => 
                           out_imux_6_48_port, B(47) => out_imux_6_47_port, 
                           B(46) => out_imux_6_46_port, B(45) => 
                           out_imux_6_45_port, B(44) => out_imux_6_44_port, 
                           B(43) => out_imux_6_43_port, B(42) => 
                           out_imux_6_42_port, B(41) => out_imux_6_41_port, 
                           B(40) => out_imux_6_40_port, B(39) => 
                           out_imux_6_39_port, B(38) => out_imux_6_38_port, 
                           B(37) => out_imux_6_37_port, B(36) => 
                           out_imux_6_36_port, B(35) => out_imux_6_35_port, 
                           B(34) => out_imux_6_34_port, B(33) => 
                           out_imux_6_33_port, B(32) => out_imux_6_32_port, 
                           B(31) => out_imux_6_31_port, B(30) => 
                           out_imux_6_30_port, B(29) => out_imux_6_29_port, 
                           B(28) => out_imux_6_28_port, B(27) => 
                           out_imux_6_27_port, B(26) => out_imux_6_26_port, 
                           B(25) => out_imux_6_25_port, B(24) => 
                           out_imux_6_24_port, B(23) => out_imux_6_23_port, 
                           B(22) => out_imux_6_22_port, B(21) => 
                           out_imux_6_21_port, B(20) => out_imux_6_20_port, 
                           B(19) => out_imux_6_19_port, B(18) => 
                           out_imux_6_18_port, B(17) => out_imux_6_17_port, 
                           B(16) => out_imux_6_16_port, B(15) => 
                           out_imux_6_15_port, B(14) => out_imux_6_14_port, 
                           B(13) => out_imux_6_13_port, B(12) => 
                           out_imux_6_12_port, B(11) => out_imux_6_11_port, 
                           B(10) => out_imux_6_10_port, B(9) => 
                           out_imux_6_9_port, B(8) => out_imux_6_8_port, B(7) 
                           => out_imux_6_7_port, B(6) => out_imux_6_6_port, 
                           B(5) => out_imux_6_5_port, B(4) => out_imux_6_4_port
                           , B(3) => out_imux_6_3_port, B(2) => 
                           out_imux_6_2_port, B(1) => out_imux_6_1_port, B(0) 
                           => out_imux_6_0_port, Ci => X_Logic0_port, S(63) => 
                           predigest_product_6_63_port, S(62) => 
                           predigest_product_6_62_port, S(61) => 
                           predigest_product_6_61_port, S(60) => 
                           predigest_product_6_60_port, S(59) => 
                           predigest_product_6_59_port, S(58) => 
                           predigest_product_6_58_port, S(57) => 
                           predigest_product_6_57_port, S(56) => 
                           predigest_product_6_56_port, S(55) => 
                           predigest_product_6_55_port, S(54) => 
                           predigest_product_6_54_port, S(53) => 
                           predigest_product_6_53_port, S(52) => 
                           predigest_product_6_52_port, S(51) => 
                           predigest_product_6_51_port, S(50) => 
                           predigest_product_6_50_port, S(49) => 
                           predigest_product_6_49_port, S(48) => 
                           predigest_product_6_48_port, S(47) => 
                           predigest_product_6_47_port, S(46) => 
                           predigest_product_6_46_port, S(45) => 
                           predigest_product_6_45_port, S(44) => 
                           predigest_product_6_44_port, S(43) => 
                           predigest_product_6_43_port, S(42) => 
                           predigest_product_6_42_port, S(41) => 
                           predigest_product_6_41_port, S(40) => 
                           predigest_product_6_40_port, S(39) => 
                           predigest_product_6_39_port, S(38) => 
                           predigest_product_6_38_port, S(37) => 
                           predigest_product_6_37_port, S(36) => 
                           predigest_product_6_36_port, S(35) => 
                           predigest_product_6_35_port, S(34) => 
                           predigest_product_6_34_port, S(33) => 
                           predigest_product_6_33_port, S(32) => 
                           predigest_product_6_32_port, S(31) => 
                           predigest_product_6_31_port, S(30) => 
                           predigest_product_6_30_port, S(29) => 
                           predigest_product_6_29_port, S(28) => 
                           predigest_product_6_28_port, S(27) => 
                           predigest_product_6_27_port, S(26) => 
                           predigest_product_6_26_port, S(25) => 
                           predigest_product_6_25_port, S(24) => 
                           predigest_product_6_24_port, S(23) => 
                           predigest_product_6_23_port, S(22) => 
                           predigest_product_6_22_port, S(21) => 
                           predigest_product_6_21_port, S(20) => 
                           predigest_product_6_20_port, S(19) => 
                           predigest_product_6_19_port, S(18) => 
                           predigest_product_6_18_port, S(17) => 
                           predigest_product_6_17_port, S(16) => 
                           predigest_product_6_16_port, S(15) => 
                           predigest_product_6_15_port, S(14) => 
                           predigest_product_6_14_port, S(13) => 
                           predigest_product_6_13_port, S(12) => 
                           predigest_product_6_12_port, S(11) => 
                           predigest_product_6_11_port, S(10) => 
                           predigest_product_6_10_port, S(9) => 
                           predigest_product_6_9_port, S(8) => 
                           predigest_product_6_8_port, S(7) => 
                           predigest_product_6_7_port, S(6) => 
                           predigest_product_6_6_port, S(5) => 
                           predigest_product_6_5_port, S(4) => 
                           predigest_product_6_4_port, S(3) => 
                           predigest_product_6_3_port, S(2) => 
                           predigest_product_6_2_port, S(1) => 
                           predigest_product_6_1_port, S(0) => 
                           predigest_product_6_0_port, Co => n_1097);
   ENC_i_7 : BOOTH_ENCODER_3BIT_13 port map( B(2) => B(15), B(1) => B(14), B(0)
                           => B(13), ENCODED(2) => 
                           muxs_encoded_signals_7_2_port, ENCODED(1) => 
                           muxs_encoded_signals_7_1_port, ENCODED(0) => 
                           muxs_encoded_signals_7_0_port);
   MUX_i_7 : MUX51_GENERIC_NBIT64_9 port map( IN0(63) => X_Logic0_port, IN0(62)
                           => X_Logic0_port, IN0(61) => X_Logic0_port, IN0(60) 
                           => X_Logic0_port, IN0(59) => X_Logic0_port, IN0(58) 
                           => X_Logic0_port, IN0(57) => X_Logic0_port, IN0(56) 
                           => X_Logic0_port, IN0(55) => X_Logic0_port, IN0(54) 
                           => X_Logic0_port, IN0(53) => X_Logic0_port, IN0(52) 
                           => X_Logic0_port, IN0(51) => X_Logic0_port, IN0(50) 
                           => X_Logic0_port, IN0(49) => X_Logic0_port, IN0(48) 
                           => X_Logic0_port, IN0(47) => X_Logic0_port, IN0(46) 
                           => X_Logic0_port, IN0(45) => X_Logic0_port, IN0(44) 
                           => X_Logic0_port, IN0(43) => X_Logic0_port, IN0(42) 
                           => X_Logic0_port, IN0(41) => X_Logic0_port, IN0(40) 
                           => X_Logic0_port, IN0(39) => X_Logic0_port, IN0(38) 
                           => X_Logic0_port, IN0(37) => X_Logic0_port, IN0(36) 
                           => X_Logic0_port, IN0(35) => X_Logic0_port, IN0(34) 
                           => X_Logic0_port, IN0(33) => X_Logic0_port, IN0(32) 
                           => X_Logic0_port, IN0(31) => X_Logic0_port, IN0(30) 
                           => X_Logic0_port, IN0(29) => X_Logic0_port, IN0(28) 
                           => X_Logic0_port, IN0(27) => X_Logic0_port, IN0(26) 
                           => X_Logic0_port, IN0(25) => X_Logic0_port, IN0(24) 
                           => X_Logic0_port, IN0(23) => X_Logic0_port, IN0(22) 
                           => X_Logic0_port, IN0(21) => X_Logic0_port, IN0(20) 
                           => X_Logic0_port, IN0(19) => X_Logic0_port, IN0(18) 
                           => X_Logic0_port, IN0(17) => X_Logic0_port, IN0(16) 
                           => X_Logic0_port, IN0(15) => X_Logic0_port, IN0(14) 
                           => X_Logic0_port, IN0(13) => X_Logic0_port, IN0(12) 
                           => X_Logic0_port, IN0(11) => X_Logic0_port, IN0(10) 
                           => X_Logic0_port, IN0(9) => X_Logic0_port, IN0(8) =>
                           X_Logic0_port, IN0(7) => X_Logic0_port, IN0(6) => 
                           X_Logic0_port, IN0(5) => X_Logic0_port, IN0(4) => 
                           X_Logic0_port, IN0(3) => X_Logic0_port, IN0(2) => 
                           X_Logic0_port, IN0(1) => X_Logic0_port, IN0(0) => 
                           X_Logic0_port, IN1(63) => A(31), IN1(62) => A(31), 
                           IN1(61) => A(31), IN1(60) => A(31), IN1(59) => A(31)
                           , IN1(58) => A(31), IN1(57) => A(31), IN1(56) => 
                           A(31), IN1(55) => A(31), IN1(54) => A(31), IN1(53) 
                           => A(31), IN1(52) => A(31), IN1(51) => A(31), 
                           IN1(50) => A(31), IN1(49) => A(31), IN1(48) => A(31)
                           , IN1(47) => A(31), IN1(46) => A(31), IN1(45) => 
                           A(31), IN1(44) => A(30), IN1(43) => A(29), IN1(42) 
                           => A(28), IN1(41) => A(27), IN1(40) => A(26), 
                           IN1(39) => A(25), IN1(38) => A(24), IN1(37) => A(23)
                           , IN1(36) => A(22), IN1(35) => A(21), IN1(34) => 
                           A(20), IN1(33) => A(19), IN1(32) => A(18), IN1(31) 
                           => A(17), IN1(30) => A(16), IN1(29) => A(15), 
                           IN1(28) => A(14), IN1(27) => A(13), IN1(26) => A(12)
                           , IN1(25) => A(11), IN1(24) => A(10), IN1(23) => 
                           A(9), IN1(22) => A(8), IN1(21) => A(7), IN1(20) => 
                           A(6), IN1(19) => A(5), IN1(18) => A(4), IN1(17) => 
                           A(3), IN1(16) => A(2), IN1(15) => A(1), IN1(14) => 
                           A(0), IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(63) => negative_a_49_port, 
                           IN2(62) => negative_a_48_port, IN2(61) => 
                           negative_a_47_port, IN2(60) => negative_a_46_port, 
                           IN2(59) => negative_a_45_port, IN2(58) => 
                           negative_a_44_port, IN2(57) => negative_a_43_port, 
                           IN2(56) => negative_a_42_port, IN2(55) => 
                           negative_a_41_port, IN2(54) => negative_a_40_port, 
                           IN2(53) => negative_a_39_port, IN2(52) => 
                           negative_a_38_port, IN2(51) => negative_a_37_port, 
                           IN2(50) => negative_a_36_port, IN2(49) => 
                           negative_a_35_port, IN2(48) => negative_a_34_port, 
                           IN2(47) => n37, IN2(46) => n34, IN2(45) => 
                           negative_a_31_port, IN2(44) => negative_a_30_port, 
                           IN2(43) => negative_a_29_port, IN2(42) => 
                           negative_a_28_port, IN2(41) => negative_a_27_port, 
                           IN2(40) => negative_a_26_port, IN2(39) => 
                           negative_a_25_port, IN2(38) => negative_a_24_port, 
                           IN2(37) => negative_a_23_port, IN2(36) => 
                           negative_a_22_port, IN2(35) => negative_a_21_port, 
                           IN2(34) => negative_a_20_port, IN2(33) => 
                           negative_a_19_port, IN2(32) => negative_a_18_port, 
                           IN2(31) => negative_a_17_port, IN2(30) => 
                           negative_a_16_port, IN2(29) => negative_a_15_port, 
                           IN2(28) => negative_a_14_port, IN2(27) => 
                           negative_a_13_port, IN2(26) => negative_a_12_port, 
                           IN2(25) => negative_a_11_port, IN2(24) => 
                           negative_a_10_port, IN2(23) => negative_a_9_port, 
                           IN2(22) => negative_a_8_port, IN2(21) => 
                           negative_a_7_port, IN2(20) => negative_a_6_port, 
                           IN2(19) => negative_a_5_port, IN2(18) => 
                           negative_a_4_port, IN2(17) => negative_a_3_port, 
                           IN2(16) => negative_a_2_port, IN2(15) => 
                           negative_a_1_port, IN2(14) => negative_a_0_port, 
                           IN2(13) => X_Logic0_port, IN2(12) => X_Logic0_port, 
                           IN2(11) => X_Logic0_port, IN2(10) => X_Logic0_port, 
                           IN2(9) => X_Logic0_port, IN2(8) => X_Logic0_port, 
                           IN2(7) => X_Logic0_port, IN2(6) => X_Logic0_port, 
                           IN2(5) => X_Logic0_port, IN2(4) => X_Logic0_port, 
                           IN2(3) => X_Logic0_port, IN2(2) => X_Logic0_port, 
                           IN2(1) => X_Logic0_port, IN2(0) => X_Logic0_port, 
                           IN3(63) => A(31), IN3(62) => A(31), IN3(61) => A(31)
                           , IN3(60) => A(31), IN3(59) => A(31), IN3(58) => 
                           A(31), IN3(57) => A(31), IN3(56) => A(31), IN3(55) 
                           => A(31), IN3(54) => A(31), IN3(53) => A(31), 
                           IN3(52) => A(31), IN3(51) => A(31), IN3(50) => A(31)
                           , IN3(49) => A(31), IN3(48) => A(31), IN3(47) => 
                           A(31), IN3(46) => A(31), IN3(45) => A(30), IN3(44) 
                           => A(29), IN3(43) => A(28), IN3(42) => A(27), 
                           IN3(41) => A(26), IN3(40) => A(25), IN3(39) => A(24)
                           , IN3(38) => A(23), IN3(37) => A(22), IN3(36) => 
                           A(21), IN3(35) => A(20), IN3(34) => A(19), IN3(33) 
                           => A(18), IN3(32) => A(17), IN3(31) => A(16), 
                           IN3(30) => A(15), IN3(29) => A(14), IN3(28) => A(13)
                           , IN3(27) => A(12), IN3(26) => A(11), IN3(25) => 
                           A(10), IN3(24) => A(9), IN3(23) => A(8), IN3(22) => 
                           A(7), IN3(21) => A(6), IN3(20) => A(5), IN3(19) => 
                           A(4), IN3(18) => A(3), IN3(17) => A(2), IN3(16) => 
                           A(1), IN3(15) => A(0), IN3(14) => X_Logic0_port, 
                           IN3(13) => X_Logic0_port, IN3(12) => X_Logic0_port, 
                           IN3(11) => X_Logic0_port, IN3(10) => X_Logic0_port, 
                           IN3(9) => X_Logic0_port, IN3(8) => X_Logic0_port, 
                           IN3(7) => X_Logic0_port, IN3(6) => X_Logic0_port, 
                           IN3(5) => X_Logic0_port, IN3(4) => X_Logic0_port, 
                           IN3(3) => X_Logic0_port, IN3(2) => X_Logic0_port, 
                           IN3(1) => X_Logic0_port, IN3(0) => X_Logic0_port, 
                           IN4(63) => negative_a_48_port, IN4(62) => 
                           negative_a_47_port, IN4(61) => negative_a_46_port, 
                           IN4(60) => negative_a_45_port, IN4(59) => 
                           negative_a_44_port, IN4(58) => negative_a_43_port, 
                           IN4(57) => negative_a_42_port, IN4(56) => 
                           negative_a_41_port, IN4(55) => negative_a_40_port, 
                           IN4(54) => negative_a_39_port, IN4(53) => 
                           negative_a_38_port, IN4(52) => negative_a_37_port, 
                           IN4(51) => negative_a_36_port, IN4(50) => 
                           negative_a_35_port, IN4(49) => negative_a_34_port, 
                           IN4(48) => n37, IN4(47) => n34, IN4(46) => 
                           negative_a_31_port, IN4(45) => negative_a_30_port, 
                           IN4(44) => negative_a_29_port, IN4(43) => 
                           negative_a_28_port, IN4(42) => negative_a_27_port, 
                           IN4(41) => negative_a_26_port, IN4(40) => 
                           negative_a_25_port, IN4(39) => negative_a_24_port, 
                           IN4(38) => negative_a_23_port, IN4(37) => 
                           negative_a_22_port, IN4(36) => negative_a_21_port, 
                           IN4(35) => negative_a_20_port, IN4(34) => 
                           negative_a_19_port, IN4(33) => negative_a_18_port, 
                           IN4(32) => negative_a_17_port, IN4(31) => 
                           negative_a_16_port, IN4(30) => negative_a_15_port, 
                           IN4(29) => negative_a_14_port, IN4(28) => 
                           negative_a_13_port, IN4(27) => negative_a_12_port, 
                           IN4(26) => negative_a_11_port, IN4(25) => 
                           negative_a_10_port, IN4(24) => negative_a_9_port, 
                           IN4(23) => negative_a_8_port, IN4(22) => 
                           negative_a_7_port, IN4(21) => negative_a_6_port, 
                           IN4(20) => negative_a_5_port, IN4(19) => 
                           negative_a_4_port, IN4(18) => negative_a_3_port, 
                           IN4(17) => negative_a_2_port, IN4(16) => 
                           negative_a_1_port, IN4(15) => negative_a_0_port, 
                           IN4(14) => X_Logic0_port, IN4(13) => X_Logic0_port, 
                           IN4(12) => X_Logic0_port, IN4(11) => X_Logic0_port, 
                           IN4(10) => X_Logic0_port, IN4(9) => X_Logic0_port, 
                           IN4(8) => X_Logic0_port, IN4(7) => X_Logic0_port, 
                           IN4(6) => X_Logic0_port, IN4(5) => X_Logic0_port, 
                           IN4(4) => X_Logic0_port, IN4(3) => X_Logic0_port, 
                           IN4(2) => X_Logic0_port, IN4(1) => X_Logic0_port, 
                           IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_7_2_port, S(1) => 
                           muxs_encoded_signals_7_1_port, S(0) => 
                           muxs_encoded_signals_7_0_port, O(63) => 
                           out_imux_7_63_port, O(62) => out_imux_7_62_port, 
                           O(61) => out_imux_7_61_port, O(60) => 
                           out_imux_7_60_port, O(59) => out_imux_7_59_port, 
                           O(58) => out_imux_7_58_port, O(57) => 
                           out_imux_7_57_port, O(56) => out_imux_7_56_port, 
                           O(55) => out_imux_7_55_port, O(54) => 
                           out_imux_7_54_port, O(53) => out_imux_7_53_port, 
                           O(52) => out_imux_7_52_port, O(51) => 
                           out_imux_7_51_port, O(50) => out_imux_7_50_port, 
                           O(49) => out_imux_7_49_port, O(48) => 
                           out_imux_7_48_port, O(47) => out_imux_7_47_port, 
                           O(46) => out_imux_7_46_port, O(45) => 
                           out_imux_7_45_port, O(44) => out_imux_7_44_port, 
                           O(43) => out_imux_7_43_port, O(42) => 
                           out_imux_7_42_port, O(41) => out_imux_7_41_port, 
                           O(40) => out_imux_7_40_port, O(39) => 
                           out_imux_7_39_port, O(38) => out_imux_7_38_port, 
                           O(37) => out_imux_7_37_port, O(36) => 
                           out_imux_7_36_port, O(35) => out_imux_7_35_port, 
                           O(34) => out_imux_7_34_port, O(33) => 
                           out_imux_7_33_port, O(32) => out_imux_7_32_port, 
                           O(31) => out_imux_7_31_port, O(30) => 
                           out_imux_7_30_port, O(29) => out_imux_7_29_port, 
                           O(28) => out_imux_7_28_port, O(27) => 
                           out_imux_7_27_port, O(26) => out_imux_7_26_port, 
                           O(25) => out_imux_7_25_port, O(24) => 
                           out_imux_7_24_port, O(23) => out_imux_7_23_port, 
                           O(22) => out_imux_7_22_port, O(21) => 
                           out_imux_7_21_port, O(20) => out_imux_7_20_port, 
                           O(19) => out_imux_7_19_port, O(18) => 
                           out_imux_7_18_port, O(17) => out_imux_7_17_port, 
                           O(16) => out_imux_7_16_port, O(15) => 
                           out_imux_7_15_port, O(14) => out_imux_7_14_port, 
                           O(13) => out_imux_7_13_port, O(12) => 
                           out_imux_7_12_port, O(11) => out_imux_7_11_port, 
                           O(10) => out_imux_7_10_port, O(9) => 
                           out_imux_7_9_port, O(8) => out_imux_7_8_port, O(7) 
                           => out_imux_7_7_port, O(6) => out_imux_7_6_port, 
                           O(5) => out_imux_7_5_port, O(4) => out_imux_7_4_port
                           , O(3) => out_imux_7_3_port, O(2) => 
                           out_imux_7_2_port, O(1) => out_imux_7_1_port, O(0) 
                           => out_imux_7_0_port);
   ADD64_i_7 : RCA_GENERIC_NBIT64_9 port map( A(63) => 
                           predigest_product_6_63_port, A(62) => 
                           predigest_product_6_62_port, A(61) => 
                           predigest_product_6_61_port, A(60) => 
                           predigest_product_6_60_port, A(59) => 
                           predigest_product_6_59_port, A(58) => 
                           predigest_product_6_58_port, A(57) => 
                           predigest_product_6_57_port, A(56) => 
                           predigest_product_6_56_port, A(55) => 
                           predigest_product_6_55_port, A(54) => 
                           predigest_product_6_54_port, A(53) => 
                           predigest_product_6_53_port, A(52) => 
                           predigest_product_6_52_port, A(51) => 
                           predigest_product_6_51_port, A(50) => 
                           predigest_product_6_50_port, A(49) => 
                           predigest_product_6_49_port, A(48) => 
                           predigest_product_6_48_port, A(47) => 
                           predigest_product_6_47_port, A(46) => 
                           predigest_product_6_46_port, A(45) => 
                           predigest_product_6_45_port, A(44) => 
                           predigest_product_6_44_port, A(43) => 
                           predigest_product_6_43_port, A(42) => 
                           predigest_product_6_42_port, A(41) => 
                           predigest_product_6_41_port, A(40) => 
                           predigest_product_6_40_port, A(39) => 
                           predigest_product_6_39_port, A(38) => 
                           predigest_product_6_38_port, A(37) => 
                           predigest_product_6_37_port, A(36) => 
                           predigest_product_6_36_port, A(35) => 
                           predigest_product_6_35_port, A(34) => 
                           predigest_product_6_34_port, A(33) => 
                           predigest_product_6_33_port, A(32) => 
                           predigest_product_6_32_port, A(31) => 
                           predigest_product_6_31_port, A(30) => 
                           predigest_product_6_30_port, A(29) => 
                           predigest_product_6_29_port, A(28) => 
                           predigest_product_6_28_port, A(27) => 
                           predigest_product_6_27_port, A(26) => 
                           predigest_product_6_26_port, A(25) => 
                           predigest_product_6_25_port, A(24) => 
                           predigest_product_6_24_port, A(23) => 
                           predigest_product_6_23_port, A(22) => 
                           predigest_product_6_22_port, A(21) => 
                           predigest_product_6_21_port, A(20) => 
                           predigest_product_6_20_port, A(19) => 
                           predigest_product_6_19_port, A(18) => 
                           predigest_product_6_18_port, A(17) => 
                           predigest_product_6_17_port, A(16) => 
                           predigest_product_6_16_port, A(15) => 
                           predigest_product_6_15_port, A(14) => 
                           predigest_product_6_14_port, A(13) => 
                           predigest_product_6_13_port, A(12) => 
                           predigest_product_6_12_port, A(11) => 
                           predigest_product_6_11_port, A(10) => 
                           predigest_product_6_10_port, A(9) => 
                           predigest_product_6_9_port, A(8) => 
                           predigest_product_6_8_port, A(7) => 
                           predigest_product_6_7_port, A(6) => 
                           predigest_product_6_6_port, A(5) => 
                           predigest_product_6_5_port, A(4) => 
                           predigest_product_6_4_port, A(3) => 
                           predigest_product_6_3_port, A(2) => 
                           predigest_product_6_2_port, A(1) => 
                           predigest_product_6_1_port, A(0) => 
                           predigest_product_6_0_port, B(63) => 
                           out_imux_7_63_port, B(62) => out_imux_7_62_port, 
                           B(61) => out_imux_7_61_port, B(60) => 
                           out_imux_7_60_port, B(59) => out_imux_7_59_port, 
                           B(58) => out_imux_7_58_port, B(57) => 
                           out_imux_7_57_port, B(56) => out_imux_7_56_port, 
                           B(55) => out_imux_7_55_port, B(54) => 
                           out_imux_7_54_port, B(53) => out_imux_7_53_port, 
                           B(52) => out_imux_7_52_port, B(51) => 
                           out_imux_7_51_port, B(50) => out_imux_7_50_port, 
                           B(49) => out_imux_7_49_port, B(48) => 
                           out_imux_7_48_port, B(47) => out_imux_7_47_port, 
                           B(46) => out_imux_7_46_port, B(45) => 
                           out_imux_7_45_port, B(44) => out_imux_7_44_port, 
                           B(43) => out_imux_7_43_port, B(42) => 
                           out_imux_7_42_port, B(41) => out_imux_7_41_port, 
                           B(40) => out_imux_7_40_port, B(39) => 
                           out_imux_7_39_port, B(38) => out_imux_7_38_port, 
                           B(37) => out_imux_7_37_port, B(36) => 
                           out_imux_7_36_port, B(35) => out_imux_7_35_port, 
                           B(34) => out_imux_7_34_port, B(33) => 
                           out_imux_7_33_port, B(32) => out_imux_7_32_port, 
                           B(31) => out_imux_7_31_port, B(30) => 
                           out_imux_7_30_port, B(29) => out_imux_7_29_port, 
                           B(28) => out_imux_7_28_port, B(27) => 
                           out_imux_7_27_port, B(26) => out_imux_7_26_port, 
                           B(25) => out_imux_7_25_port, B(24) => 
                           out_imux_7_24_port, B(23) => out_imux_7_23_port, 
                           B(22) => out_imux_7_22_port, B(21) => 
                           out_imux_7_21_port, B(20) => out_imux_7_20_port, 
                           B(19) => out_imux_7_19_port, B(18) => 
                           out_imux_7_18_port, B(17) => out_imux_7_17_port, 
                           B(16) => out_imux_7_16_port, B(15) => 
                           out_imux_7_15_port, B(14) => out_imux_7_14_port, 
                           B(13) => out_imux_7_13_port, B(12) => 
                           out_imux_7_12_port, B(11) => out_imux_7_11_port, 
                           B(10) => out_imux_7_10_port, B(9) => 
                           out_imux_7_9_port, B(8) => out_imux_7_8_port, B(7) 
                           => out_imux_7_7_port, B(6) => out_imux_7_6_port, 
                           B(5) => out_imux_7_5_port, B(4) => out_imux_7_4_port
                           , B(3) => out_imux_7_3_port, B(2) => 
                           out_imux_7_2_port, B(1) => out_imux_7_1_port, B(0) 
                           => out_imux_7_0_port, Ci => X_Logic0_port, S(63) => 
                           predigest_product_7_63_port, S(62) => 
                           predigest_product_7_62_port, S(61) => 
                           predigest_product_7_61_port, S(60) => 
                           predigest_product_7_60_port, S(59) => 
                           predigest_product_7_59_port, S(58) => 
                           predigest_product_7_58_port, S(57) => 
                           predigest_product_7_57_port, S(56) => 
                           predigest_product_7_56_port, S(55) => 
                           predigest_product_7_55_port, S(54) => 
                           predigest_product_7_54_port, S(53) => 
                           predigest_product_7_53_port, S(52) => 
                           predigest_product_7_52_port, S(51) => 
                           predigest_product_7_51_port, S(50) => 
                           predigest_product_7_50_port, S(49) => 
                           predigest_product_7_49_port, S(48) => 
                           predigest_product_7_48_port, S(47) => 
                           predigest_product_7_47_port, S(46) => 
                           predigest_product_7_46_port, S(45) => 
                           predigest_product_7_45_port, S(44) => 
                           predigest_product_7_44_port, S(43) => 
                           predigest_product_7_43_port, S(42) => 
                           predigest_product_7_42_port, S(41) => 
                           predigest_product_7_41_port, S(40) => 
                           predigest_product_7_40_port, S(39) => 
                           predigest_product_7_39_port, S(38) => 
                           predigest_product_7_38_port, S(37) => 
                           predigest_product_7_37_port, S(36) => 
                           predigest_product_7_36_port, S(35) => 
                           predigest_product_7_35_port, S(34) => 
                           predigest_product_7_34_port, S(33) => 
                           predigest_product_7_33_port, S(32) => 
                           predigest_product_7_32_port, S(31) => 
                           predigest_product_7_31_port, S(30) => 
                           predigest_product_7_30_port, S(29) => 
                           predigest_product_7_29_port, S(28) => 
                           predigest_product_7_28_port, S(27) => 
                           predigest_product_7_27_port, S(26) => 
                           predigest_product_7_26_port, S(25) => 
                           predigest_product_7_25_port, S(24) => 
                           predigest_product_7_24_port, S(23) => 
                           predigest_product_7_23_port, S(22) => 
                           predigest_product_7_22_port, S(21) => 
                           predigest_product_7_21_port, S(20) => 
                           predigest_product_7_20_port, S(19) => 
                           predigest_product_7_19_port, S(18) => 
                           predigest_product_7_18_port, S(17) => 
                           predigest_product_7_17_port, S(16) => 
                           predigest_product_7_16_port, S(15) => 
                           predigest_product_7_15_port, S(14) => 
                           predigest_product_7_14_port, S(13) => 
                           predigest_product_7_13_port, S(12) => 
                           predigest_product_7_12_port, S(11) => 
                           predigest_product_7_11_port, S(10) => 
                           predigest_product_7_10_port, S(9) => 
                           predigest_product_7_9_port, S(8) => 
                           predigest_product_7_8_port, S(7) => 
                           predigest_product_7_7_port, S(6) => 
                           predigest_product_7_6_port, S(5) => 
                           predigest_product_7_5_port, S(4) => 
                           predigest_product_7_4_port, S(3) => 
                           predigest_product_7_3_port, S(2) => 
                           predigest_product_7_2_port, S(1) => 
                           predigest_product_7_1_port, S(0) => 
                           predigest_product_7_0_port, Co => n_1098);
   ENC_i_8 : BOOTH_ENCODER_3BIT_12 port map( B(2) => B(17), B(1) => B(16), B(0)
                           => B(15), ENCODED(2) => 
                           muxs_encoded_signals_8_2_port, ENCODED(1) => 
                           muxs_encoded_signals_8_1_port, ENCODED(0) => 
                           muxs_encoded_signals_8_0_port);
   MUX_i_8 : MUX51_GENERIC_NBIT64_8 port map( IN0(63) => X_Logic0_port, IN0(62)
                           => X_Logic0_port, IN0(61) => X_Logic0_port, IN0(60) 
                           => X_Logic0_port, IN0(59) => X_Logic0_port, IN0(58) 
                           => X_Logic0_port, IN0(57) => X_Logic0_port, IN0(56) 
                           => X_Logic0_port, IN0(55) => X_Logic0_port, IN0(54) 
                           => X_Logic0_port, IN0(53) => X_Logic0_port, IN0(52) 
                           => X_Logic0_port, IN0(51) => X_Logic0_port, IN0(50) 
                           => X_Logic0_port, IN0(49) => X_Logic0_port, IN0(48) 
                           => X_Logic0_port, IN0(47) => X_Logic0_port, IN0(46) 
                           => X_Logic0_port, IN0(45) => X_Logic0_port, IN0(44) 
                           => X_Logic0_port, IN0(43) => X_Logic0_port, IN0(42) 
                           => X_Logic0_port, IN0(41) => X_Logic0_port, IN0(40) 
                           => X_Logic0_port, IN0(39) => X_Logic0_port, IN0(38) 
                           => X_Logic0_port, IN0(37) => X_Logic0_port, IN0(36) 
                           => X_Logic0_port, IN0(35) => X_Logic0_port, IN0(34) 
                           => X_Logic0_port, IN0(33) => X_Logic0_port, IN0(32) 
                           => X_Logic0_port, IN0(31) => X_Logic0_port, IN0(30) 
                           => X_Logic0_port, IN0(29) => X_Logic0_port, IN0(28) 
                           => X_Logic0_port, IN0(27) => X_Logic0_port, IN0(26) 
                           => X_Logic0_port, IN0(25) => X_Logic0_port, IN0(24) 
                           => X_Logic0_port, IN0(23) => X_Logic0_port, IN0(22) 
                           => X_Logic0_port, IN0(21) => X_Logic0_port, IN0(20) 
                           => X_Logic0_port, IN0(19) => X_Logic0_port, IN0(18) 
                           => X_Logic0_port, IN0(17) => X_Logic0_port, IN0(16) 
                           => X_Logic0_port, IN0(15) => X_Logic0_port, IN0(14) 
                           => X_Logic0_port, IN0(13) => X_Logic0_port, IN0(12) 
                           => X_Logic0_port, IN0(11) => X_Logic0_port, IN0(10) 
                           => X_Logic0_port, IN0(9) => X_Logic0_port, IN0(8) =>
                           X_Logic0_port, IN0(7) => X_Logic0_port, IN0(6) => 
                           X_Logic0_port, IN0(5) => X_Logic0_port, IN0(4) => 
                           X_Logic0_port, IN0(3) => X_Logic0_port, IN0(2) => 
                           X_Logic0_port, IN0(1) => X_Logic0_port, IN0(0) => 
                           X_Logic0_port, IN1(63) => A(31), IN1(62) => A(31), 
                           IN1(61) => A(31), IN1(60) => A(31), IN1(59) => A(31)
                           , IN1(58) => A(31), IN1(57) => A(31), IN1(56) => 
                           A(31), IN1(55) => A(31), IN1(54) => A(31), IN1(53) 
                           => A(31), IN1(52) => A(31), IN1(51) => A(31), 
                           IN1(50) => A(31), IN1(49) => A(31), IN1(48) => A(31)
                           , IN1(47) => A(31), IN1(46) => A(30), IN1(45) => 
                           A(29), IN1(44) => A(28), IN1(43) => A(27), IN1(42) 
                           => A(26), IN1(41) => A(25), IN1(40) => A(24), 
                           IN1(39) => A(23), IN1(38) => A(22), IN1(37) => A(21)
                           , IN1(36) => A(20), IN1(35) => A(19), IN1(34) => 
                           A(18), IN1(33) => A(17), IN1(32) => A(16), IN1(31) 
                           => A(15), IN1(30) => A(14), IN1(29) => A(13), 
                           IN1(28) => A(12), IN1(27) => A(11), IN1(26) => A(10)
                           , IN1(25) => A(9), IN1(24) => A(8), IN1(23) => A(7),
                           IN1(22) => A(6), IN1(21) => A(5), IN1(20) => A(4), 
                           IN1(19) => A(3), IN1(18) => A(2), IN1(17) => A(1), 
                           IN1(16) => A(0), IN1(15) => X_Logic0_port, IN1(14) 
                           => X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) 
                           => X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) 
                           => X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) =>
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(63) => negative_a_47_port, 
                           IN2(62) => negative_a_46_port, IN2(61) => 
                           negative_a_45_port, IN2(60) => negative_a_44_port, 
                           IN2(59) => negative_a_43_port, IN2(58) => 
                           negative_a_42_port, IN2(57) => negative_a_41_port, 
                           IN2(56) => negative_a_40_port, IN2(55) => 
                           negative_a_39_port, IN2(54) => negative_a_38_port, 
                           IN2(53) => negative_a_37_port, IN2(52) => 
                           negative_a_36_port, IN2(51) => negative_a_35_port, 
                           IN2(50) => negative_a_34_port, IN2(49) => n37, 
                           IN2(48) => n34, IN2(47) => negative_a_31_port, 
                           IN2(46) => negative_a_30_port, IN2(45) => 
                           negative_a_29_port, IN2(44) => negative_a_28_port, 
                           IN2(43) => negative_a_27_port, IN2(42) => 
                           negative_a_26_port, IN2(41) => negative_a_25_port, 
                           IN2(40) => negative_a_24_port, IN2(39) => 
                           negative_a_23_port, IN2(38) => negative_a_22_port, 
                           IN2(37) => negative_a_21_port, IN2(36) => 
                           negative_a_20_port, IN2(35) => negative_a_19_port, 
                           IN2(34) => negative_a_18_port, IN2(33) => 
                           negative_a_17_port, IN2(32) => negative_a_16_port, 
                           IN2(31) => negative_a_15_port, IN2(30) => 
                           negative_a_14_port, IN2(29) => negative_a_13_port, 
                           IN2(28) => negative_a_12_port, IN2(27) => 
                           negative_a_11_port, IN2(26) => negative_a_10_port, 
                           IN2(25) => negative_a_9_port, IN2(24) => 
                           negative_a_8_port, IN2(23) => negative_a_7_port, 
                           IN2(22) => negative_a_6_port, IN2(21) => 
                           negative_a_5_port, IN2(20) => negative_a_4_port, 
                           IN2(19) => negative_a_3_port, IN2(18) => 
                           negative_a_2_port, IN2(17) => negative_a_1_port, 
                           IN2(16) => negative_a_0_port, IN2(15) => 
                           X_Logic0_port, IN2(14) => X_Logic0_port, IN2(13) => 
                           X_Logic0_port, IN2(12) => X_Logic0_port, IN2(11) => 
                           X_Logic0_port, IN2(10) => X_Logic0_port, IN2(9) => 
                           X_Logic0_port, IN2(8) => X_Logic0_port, IN2(7) => 
                           X_Logic0_port, IN2(6) => X_Logic0_port, IN2(5) => 
                           X_Logic0_port, IN2(4) => X_Logic0_port, IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(63) => 
                           A(31), IN3(62) => A(31), IN3(61) => A(31), IN3(60) 
                           => A(31), IN3(59) => A(31), IN3(58) => A(31), 
                           IN3(57) => A(31), IN3(56) => A(31), IN3(55) => A(31)
                           , IN3(54) => A(31), IN3(53) => A(31), IN3(52) => 
                           A(31), IN3(51) => A(31), IN3(50) => A(31), IN3(49) 
                           => A(31), IN3(48) => A(31), IN3(47) => A(30), 
                           IN3(46) => A(29), IN3(45) => A(28), IN3(44) => A(27)
                           , IN3(43) => A(26), IN3(42) => A(25), IN3(41) => 
                           A(24), IN3(40) => A(23), IN3(39) => A(22), IN3(38) 
                           => A(21), IN3(37) => A(20), IN3(36) => A(19), 
                           IN3(35) => A(18), IN3(34) => A(17), IN3(33) => A(16)
                           , IN3(32) => A(15), IN3(31) => A(14), IN3(30) => 
                           A(13), IN3(29) => A(12), IN3(28) => A(11), IN3(27) 
                           => A(10), IN3(26) => A(9), IN3(25) => A(8), IN3(24) 
                           => A(7), IN3(23) => A(6), IN3(22) => A(5), IN3(21) 
                           => A(4), IN3(20) => A(3), IN3(19) => A(2), IN3(18) 
                           => A(1), IN3(17) => A(0), IN3(16) => X_Logic0_port, 
                           IN3(15) => X_Logic0_port, IN3(14) => X_Logic0_port, 
                           IN3(13) => X_Logic0_port, IN3(12) => X_Logic0_port, 
                           IN3(11) => X_Logic0_port, IN3(10) => X_Logic0_port, 
                           IN3(9) => X_Logic0_port, IN3(8) => X_Logic0_port, 
                           IN3(7) => X_Logic0_port, IN3(6) => X_Logic0_port, 
                           IN3(5) => X_Logic0_port, IN3(4) => X_Logic0_port, 
                           IN3(3) => X_Logic0_port, IN3(2) => X_Logic0_port, 
                           IN3(1) => X_Logic0_port, IN3(0) => X_Logic0_port, 
                           IN4(63) => negative_a_46_port, IN4(62) => 
                           negative_a_45_port, IN4(61) => negative_a_44_port, 
                           IN4(60) => negative_a_43_port, IN4(59) => 
                           negative_a_42_port, IN4(58) => negative_a_41_port, 
                           IN4(57) => negative_a_40_port, IN4(56) => 
                           negative_a_39_port, IN4(55) => negative_a_38_port, 
                           IN4(54) => negative_a_37_port, IN4(53) => 
                           negative_a_36_port, IN4(52) => negative_a_35_port, 
                           IN4(51) => negative_a_34_port, IN4(50) => n37, 
                           IN4(49) => n34, IN4(48) => negative_a_31_port, 
                           IN4(47) => negative_a_30_port, IN4(46) => 
                           negative_a_29_port, IN4(45) => negative_a_28_port, 
                           IN4(44) => negative_a_27_port, IN4(43) => 
                           negative_a_26_port, IN4(42) => negative_a_25_port, 
                           IN4(41) => negative_a_24_port, IN4(40) => 
                           negative_a_23_port, IN4(39) => negative_a_22_port, 
                           IN4(38) => negative_a_21_port, IN4(37) => 
                           negative_a_20_port, IN4(36) => negative_a_19_port, 
                           IN4(35) => negative_a_18_port, IN4(34) => 
                           negative_a_17_port, IN4(33) => negative_a_16_port, 
                           IN4(32) => negative_a_15_port, IN4(31) => 
                           negative_a_14_port, IN4(30) => negative_a_13_port, 
                           IN4(29) => negative_a_12_port, IN4(28) => 
                           negative_a_11_port, IN4(27) => negative_a_10_port, 
                           IN4(26) => negative_a_9_port, IN4(25) => 
                           negative_a_8_port, IN4(24) => negative_a_7_port, 
                           IN4(23) => negative_a_6_port, IN4(22) => 
                           negative_a_5_port, IN4(21) => negative_a_4_port, 
                           IN4(20) => negative_a_3_port, IN4(19) => 
                           negative_a_2_port, IN4(18) => negative_a_1_port, 
                           IN4(17) => negative_a_0_port, IN4(16) => 
                           X_Logic0_port, IN4(15) => X_Logic0_port, IN4(14) => 
                           X_Logic0_port, IN4(13) => X_Logic0_port, IN4(12) => 
                           X_Logic0_port, IN4(11) => X_Logic0_port, IN4(10) => 
                           X_Logic0_port, IN4(9) => X_Logic0_port, IN4(8) => 
                           X_Logic0_port, IN4(7) => X_Logic0_port, IN4(6) => 
                           X_Logic0_port, IN4(5) => X_Logic0_port, IN4(4) => 
                           X_Logic0_port, IN4(3) => X_Logic0_port, IN4(2) => 
                           X_Logic0_port, IN4(1) => X_Logic0_port, IN4(0) => 
                           X_Logic0_port, S(2) => muxs_encoded_signals_8_2_port
                           , S(1) => muxs_encoded_signals_8_1_port, S(0) => 
                           muxs_encoded_signals_8_0_port, O(63) => 
                           out_imux_8_63_port, O(62) => out_imux_8_62_port, 
                           O(61) => out_imux_8_61_port, O(60) => 
                           out_imux_8_60_port, O(59) => out_imux_8_59_port, 
                           O(58) => out_imux_8_58_port, O(57) => 
                           out_imux_8_57_port, O(56) => out_imux_8_56_port, 
                           O(55) => out_imux_8_55_port, O(54) => 
                           out_imux_8_54_port, O(53) => out_imux_8_53_port, 
                           O(52) => out_imux_8_52_port, O(51) => 
                           out_imux_8_51_port, O(50) => out_imux_8_50_port, 
                           O(49) => out_imux_8_49_port, O(48) => 
                           out_imux_8_48_port, O(47) => out_imux_8_47_port, 
                           O(46) => out_imux_8_46_port, O(45) => 
                           out_imux_8_45_port, O(44) => out_imux_8_44_port, 
                           O(43) => out_imux_8_43_port, O(42) => 
                           out_imux_8_42_port, O(41) => out_imux_8_41_port, 
                           O(40) => out_imux_8_40_port, O(39) => 
                           out_imux_8_39_port, O(38) => out_imux_8_38_port, 
                           O(37) => out_imux_8_37_port, O(36) => 
                           out_imux_8_36_port, O(35) => out_imux_8_35_port, 
                           O(34) => out_imux_8_34_port, O(33) => 
                           out_imux_8_33_port, O(32) => out_imux_8_32_port, 
                           O(31) => out_imux_8_31_port, O(30) => 
                           out_imux_8_30_port, O(29) => out_imux_8_29_port, 
                           O(28) => out_imux_8_28_port, O(27) => 
                           out_imux_8_27_port, O(26) => out_imux_8_26_port, 
                           O(25) => out_imux_8_25_port, O(24) => 
                           out_imux_8_24_port, O(23) => out_imux_8_23_port, 
                           O(22) => out_imux_8_22_port, O(21) => 
                           out_imux_8_21_port, O(20) => out_imux_8_20_port, 
                           O(19) => out_imux_8_19_port, O(18) => 
                           out_imux_8_18_port, O(17) => out_imux_8_17_port, 
                           O(16) => out_imux_8_16_port, O(15) => 
                           out_imux_8_15_port, O(14) => out_imux_8_14_port, 
                           O(13) => out_imux_8_13_port, O(12) => 
                           out_imux_8_12_port, O(11) => out_imux_8_11_port, 
                           O(10) => out_imux_8_10_port, O(9) => 
                           out_imux_8_9_port, O(8) => out_imux_8_8_port, O(7) 
                           => out_imux_8_7_port, O(6) => out_imux_8_6_port, 
                           O(5) => out_imux_8_5_port, O(4) => out_imux_8_4_port
                           , O(3) => out_imux_8_3_port, O(2) => 
                           out_imux_8_2_port, O(1) => out_imux_8_1_port, O(0) 
                           => out_imux_8_0_port);
   ADD64_i_8 : RCA_GENERIC_NBIT64_8 port map( A(63) => 
                           predigest_product_7_63_port, A(62) => 
                           predigest_product_7_62_port, A(61) => 
                           predigest_product_7_61_port, A(60) => 
                           predigest_product_7_60_port, A(59) => 
                           predigest_product_7_59_port, A(58) => 
                           predigest_product_7_58_port, A(57) => 
                           predigest_product_7_57_port, A(56) => 
                           predigest_product_7_56_port, A(55) => 
                           predigest_product_7_55_port, A(54) => 
                           predigest_product_7_54_port, A(53) => 
                           predigest_product_7_53_port, A(52) => 
                           predigest_product_7_52_port, A(51) => 
                           predigest_product_7_51_port, A(50) => 
                           predigest_product_7_50_port, A(49) => 
                           predigest_product_7_49_port, A(48) => 
                           predigest_product_7_48_port, A(47) => 
                           predigest_product_7_47_port, A(46) => 
                           predigest_product_7_46_port, A(45) => 
                           predigest_product_7_45_port, A(44) => 
                           predigest_product_7_44_port, A(43) => 
                           predigest_product_7_43_port, A(42) => 
                           predigest_product_7_42_port, A(41) => 
                           predigest_product_7_41_port, A(40) => 
                           predigest_product_7_40_port, A(39) => 
                           predigest_product_7_39_port, A(38) => 
                           predigest_product_7_38_port, A(37) => 
                           predigest_product_7_37_port, A(36) => 
                           predigest_product_7_36_port, A(35) => 
                           predigest_product_7_35_port, A(34) => 
                           predigest_product_7_34_port, A(33) => 
                           predigest_product_7_33_port, A(32) => 
                           predigest_product_7_32_port, A(31) => 
                           predigest_product_7_31_port, A(30) => 
                           predigest_product_7_30_port, A(29) => 
                           predigest_product_7_29_port, A(28) => 
                           predigest_product_7_28_port, A(27) => 
                           predigest_product_7_27_port, A(26) => 
                           predigest_product_7_26_port, A(25) => 
                           predigest_product_7_25_port, A(24) => 
                           predigest_product_7_24_port, A(23) => 
                           predigest_product_7_23_port, A(22) => 
                           predigest_product_7_22_port, A(21) => 
                           predigest_product_7_21_port, A(20) => 
                           predigest_product_7_20_port, A(19) => 
                           predigest_product_7_19_port, A(18) => 
                           predigest_product_7_18_port, A(17) => 
                           predigest_product_7_17_port, A(16) => 
                           predigest_product_7_16_port, A(15) => 
                           predigest_product_7_15_port, A(14) => 
                           predigest_product_7_14_port, A(13) => 
                           predigest_product_7_13_port, A(12) => 
                           predigest_product_7_12_port, A(11) => 
                           predigest_product_7_11_port, A(10) => 
                           predigest_product_7_10_port, A(9) => 
                           predigest_product_7_9_port, A(8) => 
                           predigest_product_7_8_port, A(7) => 
                           predigest_product_7_7_port, A(6) => 
                           predigest_product_7_6_port, A(5) => 
                           predigest_product_7_5_port, A(4) => 
                           predigest_product_7_4_port, A(3) => 
                           predigest_product_7_3_port, A(2) => 
                           predigest_product_7_2_port, A(1) => 
                           predigest_product_7_1_port, A(0) => 
                           predigest_product_7_0_port, B(63) => 
                           out_imux_8_63_port, B(62) => out_imux_8_62_port, 
                           B(61) => out_imux_8_61_port, B(60) => 
                           out_imux_8_60_port, B(59) => out_imux_8_59_port, 
                           B(58) => out_imux_8_58_port, B(57) => 
                           out_imux_8_57_port, B(56) => out_imux_8_56_port, 
                           B(55) => out_imux_8_55_port, B(54) => 
                           out_imux_8_54_port, B(53) => out_imux_8_53_port, 
                           B(52) => out_imux_8_52_port, B(51) => 
                           out_imux_8_51_port, B(50) => out_imux_8_50_port, 
                           B(49) => out_imux_8_49_port, B(48) => 
                           out_imux_8_48_port, B(47) => out_imux_8_47_port, 
                           B(46) => out_imux_8_46_port, B(45) => 
                           out_imux_8_45_port, B(44) => out_imux_8_44_port, 
                           B(43) => out_imux_8_43_port, B(42) => 
                           out_imux_8_42_port, B(41) => out_imux_8_41_port, 
                           B(40) => out_imux_8_40_port, B(39) => 
                           out_imux_8_39_port, B(38) => out_imux_8_38_port, 
                           B(37) => out_imux_8_37_port, B(36) => 
                           out_imux_8_36_port, B(35) => out_imux_8_35_port, 
                           B(34) => out_imux_8_34_port, B(33) => 
                           out_imux_8_33_port, B(32) => out_imux_8_32_port, 
                           B(31) => out_imux_8_31_port, B(30) => 
                           out_imux_8_30_port, B(29) => out_imux_8_29_port, 
                           B(28) => out_imux_8_28_port, B(27) => 
                           out_imux_8_27_port, B(26) => out_imux_8_26_port, 
                           B(25) => out_imux_8_25_port, B(24) => 
                           out_imux_8_24_port, B(23) => out_imux_8_23_port, 
                           B(22) => out_imux_8_22_port, B(21) => 
                           out_imux_8_21_port, B(20) => out_imux_8_20_port, 
                           B(19) => out_imux_8_19_port, B(18) => 
                           out_imux_8_18_port, B(17) => out_imux_8_17_port, 
                           B(16) => out_imux_8_16_port, B(15) => 
                           out_imux_8_15_port, B(14) => out_imux_8_14_port, 
                           B(13) => out_imux_8_13_port, B(12) => 
                           out_imux_8_12_port, B(11) => out_imux_8_11_port, 
                           B(10) => out_imux_8_10_port, B(9) => 
                           out_imux_8_9_port, B(8) => out_imux_8_8_port, B(7) 
                           => out_imux_8_7_port, B(6) => out_imux_8_6_port, 
                           B(5) => out_imux_8_5_port, B(4) => out_imux_8_4_port
                           , B(3) => out_imux_8_3_port, B(2) => 
                           out_imux_8_2_port, B(1) => out_imux_8_1_port, B(0) 
                           => out_imux_8_0_port, Ci => X_Logic0_port, S(63) => 
                           predigest_product_8_63_port, S(62) => 
                           predigest_product_8_62_port, S(61) => 
                           predigest_product_8_61_port, S(60) => 
                           predigest_product_8_60_port, S(59) => 
                           predigest_product_8_59_port, S(58) => 
                           predigest_product_8_58_port, S(57) => 
                           predigest_product_8_57_port, S(56) => 
                           predigest_product_8_56_port, S(55) => 
                           predigest_product_8_55_port, S(54) => 
                           predigest_product_8_54_port, S(53) => 
                           predigest_product_8_53_port, S(52) => 
                           predigest_product_8_52_port, S(51) => 
                           predigest_product_8_51_port, S(50) => 
                           predigest_product_8_50_port, S(49) => 
                           predigest_product_8_49_port, S(48) => 
                           predigest_product_8_48_port, S(47) => 
                           predigest_product_8_47_port, S(46) => 
                           predigest_product_8_46_port, S(45) => 
                           predigest_product_8_45_port, S(44) => 
                           predigest_product_8_44_port, S(43) => 
                           predigest_product_8_43_port, S(42) => 
                           predigest_product_8_42_port, S(41) => 
                           predigest_product_8_41_port, S(40) => 
                           predigest_product_8_40_port, S(39) => 
                           predigest_product_8_39_port, S(38) => 
                           predigest_product_8_38_port, S(37) => 
                           predigest_product_8_37_port, S(36) => 
                           predigest_product_8_36_port, S(35) => 
                           predigest_product_8_35_port, S(34) => 
                           predigest_product_8_34_port, S(33) => 
                           predigest_product_8_33_port, S(32) => 
                           predigest_product_8_32_port, S(31) => 
                           predigest_product_8_31_port, S(30) => 
                           predigest_product_8_30_port, S(29) => 
                           predigest_product_8_29_port, S(28) => 
                           predigest_product_8_28_port, S(27) => 
                           predigest_product_8_27_port, S(26) => 
                           predigest_product_8_26_port, S(25) => 
                           predigest_product_8_25_port, S(24) => 
                           predigest_product_8_24_port, S(23) => 
                           predigest_product_8_23_port, S(22) => 
                           predigest_product_8_22_port, S(21) => 
                           predigest_product_8_21_port, S(20) => 
                           predigest_product_8_20_port, S(19) => 
                           predigest_product_8_19_port, S(18) => 
                           predigest_product_8_18_port, S(17) => 
                           predigest_product_8_17_port, S(16) => 
                           predigest_product_8_16_port, S(15) => 
                           predigest_product_8_15_port, S(14) => 
                           predigest_product_8_14_port, S(13) => 
                           predigest_product_8_13_port, S(12) => 
                           predigest_product_8_12_port, S(11) => 
                           predigest_product_8_11_port, S(10) => 
                           predigest_product_8_10_port, S(9) => 
                           predigest_product_8_9_port, S(8) => 
                           predigest_product_8_8_port, S(7) => 
                           predigest_product_8_7_port, S(6) => 
                           predigest_product_8_6_port, S(5) => 
                           predigest_product_8_5_port, S(4) => 
                           predigest_product_8_4_port, S(3) => 
                           predigest_product_8_3_port, S(2) => 
                           predigest_product_8_2_port, S(1) => 
                           predigest_product_8_1_port, S(0) => 
                           predigest_product_8_0_port, Co => n_1099);
   ENC_i_9 : BOOTH_ENCODER_3BIT_11 port map( B(2) => B(19), B(1) => B(18), B(0)
                           => B(17), ENCODED(2) => 
                           muxs_encoded_signals_9_2_port, ENCODED(1) => 
                           muxs_encoded_signals_9_1_port, ENCODED(0) => 
                           muxs_encoded_signals_9_0_port);
   MUX_i_9 : MUX51_GENERIC_NBIT64_7 port map( IN0(63) => X_Logic0_port, IN0(62)
                           => X_Logic0_port, IN0(61) => X_Logic0_port, IN0(60) 
                           => X_Logic0_port, IN0(59) => X_Logic0_port, IN0(58) 
                           => X_Logic0_port, IN0(57) => X_Logic0_port, IN0(56) 
                           => X_Logic0_port, IN0(55) => X_Logic0_port, IN0(54) 
                           => X_Logic0_port, IN0(53) => X_Logic0_port, IN0(52) 
                           => X_Logic0_port, IN0(51) => X_Logic0_port, IN0(50) 
                           => X_Logic0_port, IN0(49) => X_Logic0_port, IN0(48) 
                           => X_Logic0_port, IN0(47) => X_Logic0_port, IN0(46) 
                           => X_Logic0_port, IN0(45) => X_Logic0_port, IN0(44) 
                           => X_Logic0_port, IN0(43) => X_Logic0_port, IN0(42) 
                           => X_Logic0_port, IN0(41) => X_Logic0_port, IN0(40) 
                           => X_Logic0_port, IN0(39) => X_Logic0_port, IN0(38) 
                           => X_Logic0_port, IN0(37) => X_Logic0_port, IN0(36) 
                           => X_Logic0_port, IN0(35) => X_Logic0_port, IN0(34) 
                           => X_Logic0_port, IN0(33) => X_Logic0_port, IN0(32) 
                           => X_Logic0_port, IN0(31) => X_Logic0_port, IN0(30) 
                           => X_Logic0_port, IN0(29) => X_Logic0_port, IN0(28) 
                           => X_Logic0_port, IN0(27) => X_Logic0_port, IN0(26) 
                           => X_Logic0_port, IN0(25) => X_Logic0_port, IN0(24) 
                           => X_Logic0_port, IN0(23) => X_Logic0_port, IN0(22) 
                           => X_Logic0_port, IN0(21) => X_Logic0_port, IN0(20) 
                           => X_Logic0_port, IN0(19) => X_Logic0_port, IN0(18) 
                           => X_Logic0_port, IN0(17) => X_Logic0_port, IN0(16) 
                           => X_Logic0_port, IN0(15) => X_Logic0_port, IN0(14) 
                           => X_Logic0_port, IN0(13) => X_Logic0_port, IN0(12) 
                           => X_Logic0_port, IN0(11) => X_Logic0_port, IN0(10) 
                           => X_Logic0_port, IN0(9) => X_Logic0_port, IN0(8) =>
                           X_Logic0_port, IN0(7) => X_Logic0_port, IN0(6) => 
                           X_Logic0_port, IN0(5) => X_Logic0_port, IN0(4) => 
                           X_Logic0_port, IN0(3) => X_Logic0_port, IN0(2) => 
                           X_Logic0_port, IN0(1) => X_Logic0_port, IN0(0) => 
                           X_Logic0_port, IN1(63) => A(31), IN1(62) => A(31), 
                           IN1(61) => A(31), IN1(60) => A(31), IN1(59) => A(31)
                           , IN1(58) => A(31), IN1(57) => A(31), IN1(56) => 
                           A(31), IN1(55) => A(31), IN1(54) => A(31), IN1(53) 
                           => A(31), IN1(52) => A(31), IN1(51) => A(31), 
                           IN1(50) => A(31), IN1(49) => A(31), IN1(48) => A(30)
                           , IN1(47) => A(29), IN1(46) => A(28), IN1(45) => 
                           A(27), IN1(44) => A(26), IN1(43) => A(25), IN1(42) 
                           => A(24), IN1(41) => A(23), IN1(40) => A(22), 
                           IN1(39) => A(21), IN1(38) => A(20), IN1(37) => A(19)
                           , IN1(36) => A(18), IN1(35) => A(17), IN1(34) => 
                           A(16), IN1(33) => A(15), IN1(32) => A(14), IN1(31) 
                           => A(13), IN1(30) => A(12), IN1(29) => A(11), 
                           IN1(28) => A(10), IN1(27) => A(9), IN1(26) => A(8), 
                           IN1(25) => A(7), IN1(24) => A(6), IN1(23) => A(5), 
                           IN1(22) => A(4), IN1(21) => A(3), IN1(20) => A(2), 
                           IN1(19) => A(1), IN1(18) => A(0), IN1(17) => 
                           X_Logic0_port, IN1(16) => X_Logic0_port, IN1(15) => 
                           X_Logic0_port, IN1(14) => X_Logic0_port, IN1(13) => 
                           X_Logic0_port, IN1(12) => X_Logic0_port, IN1(11) => 
                           X_Logic0_port, IN1(10) => X_Logic0_port, IN1(9) => 
                           X_Logic0_port, IN1(8) => X_Logic0_port, IN1(7) => 
                           X_Logic0_port, IN1(6) => X_Logic0_port, IN1(5) => 
                           X_Logic0_port, IN1(4) => X_Logic0_port, IN1(3) => 
                           X_Logic0_port, IN1(2) => X_Logic0_port, IN1(1) => 
                           X_Logic0_port, IN1(0) => X_Logic0_port, IN2(63) => 
                           negative_a_45_port, IN2(62) => negative_a_44_port, 
                           IN2(61) => negative_a_43_port, IN2(60) => 
                           negative_a_42_port, IN2(59) => negative_a_41_port, 
                           IN2(58) => negative_a_40_port, IN2(57) => 
                           negative_a_39_port, IN2(56) => negative_a_38_port, 
                           IN2(55) => negative_a_37_port, IN2(54) => 
                           negative_a_36_port, IN2(53) => negative_a_35_port, 
                           IN2(52) => negative_a_34_port, IN2(51) => n37, 
                           IN2(50) => n34, IN2(49) => negative_a_31_port, 
                           IN2(48) => negative_a_30_port, IN2(47) => 
                           negative_a_29_port, IN2(46) => negative_a_28_port, 
                           IN2(45) => negative_a_27_port, IN2(44) => 
                           negative_a_26_port, IN2(43) => negative_a_25_port, 
                           IN2(42) => negative_a_24_port, IN2(41) => 
                           negative_a_23_port, IN2(40) => negative_a_22_port, 
                           IN2(39) => negative_a_21_port, IN2(38) => 
                           negative_a_20_port, IN2(37) => negative_a_19_port, 
                           IN2(36) => negative_a_18_port, IN2(35) => 
                           negative_a_17_port, IN2(34) => negative_a_16_port, 
                           IN2(33) => negative_a_15_port, IN2(32) => 
                           negative_a_14_port, IN2(31) => negative_a_13_port, 
                           IN2(30) => negative_a_12_port, IN2(29) => 
                           negative_a_11_port, IN2(28) => negative_a_10_port, 
                           IN2(27) => negative_a_9_port, IN2(26) => 
                           negative_a_8_port, IN2(25) => negative_a_7_port, 
                           IN2(24) => negative_a_6_port, IN2(23) => 
                           negative_a_5_port, IN2(22) => negative_a_4_port, 
                           IN2(21) => negative_a_3_port, IN2(20) => 
                           negative_a_2_port, IN2(19) => negative_a_1_port, 
                           IN2(18) => negative_a_0_port, IN2(17) => 
                           X_Logic0_port, IN2(16) => X_Logic0_port, IN2(15) => 
                           X_Logic0_port, IN2(14) => X_Logic0_port, IN2(13) => 
                           X_Logic0_port, IN2(12) => X_Logic0_port, IN2(11) => 
                           X_Logic0_port, IN2(10) => X_Logic0_port, IN2(9) => 
                           X_Logic0_port, IN2(8) => X_Logic0_port, IN2(7) => 
                           X_Logic0_port, IN2(6) => X_Logic0_port, IN2(5) => 
                           X_Logic0_port, IN2(4) => X_Logic0_port, IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(63) => 
                           A(31), IN3(62) => A(31), IN3(61) => A(31), IN3(60) 
                           => A(31), IN3(59) => A(31), IN3(58) => A(31), 
                           IN3(57) => A(31), IN3(56) => A(31), IN3(55) => A(31)
                           , IN3(54) => A(31), IN3(53) => A(31), IN3(52) => 
                           A(31), IN3(51) => A(31), IN3(50) => A(31), IN3(49) 
                           => A(30), IN3(48) => A(29), IN3(47) => A(28), 
                           IN3(46) => A(27), IN3(45) => A(26), IN3(44) => A(25)
                           , IN3(43) => A(24), IN3(42) => A(23), IN3(41) => 
                           A(22), IN3(40) => A(21), IN3(39) => A(20), IN3(38) 
                           => A(19), IN3(37) => A(18), IN3(36) => A(17), 
                           IN3(35) => A(16), IN3(34) => A(15), IN3(33) => A(14)
                           , IN3(32) => A(13), IN3(31) => A(12), IN3(30) => 
                           A(11), IN3(29) => A(10), IN3(28) => A(9), IN3(27) =>
                           A(8), IN3(26) => A(7), IN3(25) => A(6), IN3(24) => 
                           A(5), IN3(23) => A(4), IN3(22) => A(3), IN3(21) => 
                           A(2), IN3(20) => A(1), IN3(19) => A(0), IN3(18) => 
                           X_Logic0_port, IN3(17) => X_Logic0_port, IN3(16) => 
                           X_Logic0_port, IN3(15) => X_Logic0_port, IN3(14) => 
                           X_Logic0_port, IN3(13) => X_Logic0_port, IN3(12) => 
                           X_Logic0_port, IN3(11) => X_Logic0_port, IN3(10) => 
                           X_Logic0_port, IN3(9) => X_Logic0_port, IN3(8) => 
                           X_Logic0_port, IN3(7) => X_Logic0_port, IN3(6) => 
                           X_Logic0_port, IN3(5) => X_Logic0_port, IN3(4) => 
                           X_Logic0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(63) => negative_a_44_port, 
                           IN4(62) => negative_a_43_port, IN4(61) => 
                           negative_a_42_port, IN4(60) => negative_a_41_port, 
                           IN4(59) => negative_a_40_port, IN4(58) => 
                           negative_a_39_port, IN4(57) => negative_a_38_port, 
                           IN4(56) => negative_a_37_port, IN4(55) => 
                           negative_a_36_port, IN4(54) => negative_a_35_port, 
                           IN4(53) => negative_a_34_port, IN4(52) => n37, 
                           IN4(51) => n34, IN4(50) => negative_a_31_port, 
                           IN4(49) => negative_a_30_port, IN4(48) => 
                           negative_a_29_port, IN4(47) => negative_a_28_port, 
                           IN4(46) => negative_a_27_port, IN4(45) => 
                           negative_a_26_port, IN4(44) => negative_a_25_port, 
                           IN4(43) => negative_a_24_port, IN4(42) => 
                           negative_a_23_port, IN4(41) => negative_a_22_port, 
                           IN4(40) => negative_a_21_port, IN4(39) => 
                           negative_a_20_port, IN4(38) => negative_a_19_port, 
                           IN4(37) => negative_a_18_port, IN4(36) => 
                           negative_a_17_port, IN4(35) => negative_a_16_port, 
                           IN4(34) => negative_a_15_port, IN4(33) => 
                           negative_a_14_port, IN4(32) => negative_a_13_port, 
                           IN4(31) => negative_a_12_port, IN4(30) => 
                           negative_a_11_port, IN4(29) => negative_a_10_port, 
                           IN4(28) => negative_a_9_port, IN4(27) => 
                           negative_a_8_port, IN4(26) => negative_a_7_port, 
                           IN4(25) => negative_a_6_port, IN4(24) => 
                           negative_a_5_port, IN4(23) => negative_a_4_port, 
                           IN4(22) => negative_a_3_port, IN4(21) => 
                           negative_a_2_port, IN4(20) => negative_a_1_port, 
                           IN4(19) => negative_a_0_port, IN4(18) => 
                           X_Logic0_port, IN4(17) => X_Logic0_port, IN4(16) => 
                           X_Logic0_port, IN4(15) => X_Logic0_port, IN4(14) => 
                           X_Logic0_port, IN4(13) => X_Logic0_port, IN4(12) => 
                           X_Logic0_port, IN4(11) => X_Logic0_port, IN4(10) => 
                           X_Logic0_port, IN4(9) => X_Logic0_port, IN4(8) => 
                           X_Logic0_port, IN4(7) => X_Logic0_port, IN4(6) => 
                           X_Logic0_port, IN4(5) => X_Logic0_port, IN4(4) => 
                           X_Logic0_port, IN4(3) => X_Logic0_port, IN4(2) => 
                           X_Logic0_port, IN4(1) => X_Logic0_port, IN4(0) => 
                           X_Logic0_port, S(2) => muxs_encoded_signals_9_2_port
                           , S(1) => muxs_encoded_signals_9_1_port, S(0) => 
                           muxs_encoded_signals_9_0_port, O(63) => 
                           out_imux_9_63_port, O(62) => out_imux_9_62_port, 
                           O(61) => out_imux_9_61_port, O(60) => 
                           out_imux_9_60_port, O(59) => out_imux_9_59_port, 
                           O(58) => out_imux_9_58_port, O(57) => 
                           out_imux_9_57_port, O(56) => out_imux_9_56_port, 
                           O(55) => out_imux_9_55_port, O(54) => 
                           out_imux_9_54_port, O(53) => out_imux_9_53_port, 
                           O(52) => out_imux_9_52_port, O(51) => 
                           out_imux_9_51_port, O(50) => out_imux_9_50_port, 
                           O(49) => out_imux_9_49_port, O(48) => 
                           out_imux_9_48_port, O(47) => out_imux_9_47_port, 
                           O(46) => out_imux_9_46_port, O(45) => 
                           out_imux_9_45_port, O(44) => out_imux_9_44_port, 
                           O(43) => out_imux_9_43_port, O(42) => 
                           out_imux_9_42_port, O(41) => out_imux_9_41_port, 
                           O(40) => out_imux_9_40_port, O(39) => 
                           out_imux_9_39_port, O(38) => out_imux_9_38_port, 
                           O(37) => out_imux_9_37_port, O(36) => 
                           out_imux_9_36_port, O(35) => out_imux_9_35_port, 
                           O(34) => out_imux_9_34_port, O(33) => 
                           out_imux_9_33_port, O(32) => out_imux_9_32_port, 
                           O(31) => out_imux_9_31_port, O(30) => 
                           out_imux_9_30_port, O(29) => out_imux_9_29_port, 
                           O(28) => out_imux_9_28_port, O(27) => 
                           out_imux_9_27_port, O(26) => out_imux_9_26_port, 
                           O(25) => out_imux_9_25_port, O(24) => 
                           out_imux_9_24_port, O(23) => out_imux_9_23_port, 
                           O(22) => out_imux_9_22_port, O(21) => 
                           out_imux_9_21_port, O(20) => out_imux_9_20_port, 
                           O(19) => out_imux_9_19_port, O(18) => 
                           out_imux_9_18_port, O(17) => out_imux_9_17_port, 
                           O(16) => out_imux_9_16_port, O(15) => 
                           out_imux_9_15_port, O(14) => out_imux_9_14_port, 
                           O(13) => out_imux_9_13_port, O(12) => 
                           out_imux_9_12_port, O(11) => out_imux_9_11_port, 
                           O(10) => out_imux_9_10_port, O(9) => 
                           out_imux_9_9_port, O(8) => out_imux_9_8_port, O(7) 
                           => out_imux_9_7_port, O(6) => out_imux_9_6_port, 
                           O(5) => out_imux_9_5_port, O(4) => out_imux_9_4_port
                           , O(3) => out_imux_9_3_port, O(2) => 
                           out_imux_9_2_port, O(1) => out_imux_9_1_port, O(0) 
                           => out_imux_9_0_port);
   ADD64_i_9 : RCA_GENERIC_NBIT64_7 port map( A(63) => 
                           predigest_product_8_63_port, A(62) => 
                           predigest_product_8_62_port, A(61) => 
                           predigest_product_8_61_port, A(60) => 
                           predigest_product_8_60_port, A(59) => 
                           predigest_product_8_59_port, A(58) => 
                           predigest_product_8_58_port, A(57) => 
                           predigest_product_8_57_port, A(56) => 
                           predigest_product_8_56_port, A(55) => 
                           predigest_product_8_55_port, A(54) => 
                           predigest_product_8_54_port, A(53) => 
                           predigest_product_8_53_port, A(52) => 
                           predigest_product_8_52_port, A(51) => 
                           predigest_product_8_51_port, A(50) => 
                           predigest_product_8_50_port, A(49) => 
                           predigest_product_8_49_port, A(48) => 
                           predigest_product_8_48_port, A(47) => 
                           predigest_product_8_47_port, A(46) => 
                           predigest_product_8_46_port, A(45) => 
                           predigest_product_8_45_port, A(44) => 
                           predigest_product_8_44_port, A(43) => 
                           predigest_product_8_43_port, A(42) => 
                           predigest_product_8_42_port, A(41) => 
                           predigest_product_8_41_port, A(40) => 
                           predigest_product_8_40_port, A(39) => 
                           predigest_product_8_39_port, A(38) => 
                           predigest_product_8_38_port, A(37) => 
                           predigest_product_8_37_port, A(36) => 
                           predigest_product_8_36_port, A(35) => 
                           predigest_product_8_35_port, A(34) => 
                           predigest_product_8_34_port, A(33) => 
                           predigest_product_8_33_port, A(32) => 
                           predigest_product_8_32_port, A(31) => 
                           predigest_product_8_31_port, A(30) => 
                           predigest_product_8_30_port, A(29) => 
                           predigest_product_8_29_port, A(28) => 
                           predigest_product_8_28_port, A(27) => 
                           predigest_product_8_27_port, A(26) => 
                           predigest_product_8_26_port, A(25) => 
                           predigest_product_8_25_port, A(24) => 
                           predigest_product_8_24_port, A(23) => 
                           predigest_product_8_23_port, A(22) => 
                           predigest_product_8_22_port, A(21) => 
                           predigest_product_8_21_port, A(20) => 
                           predigest_product_8_20_port, A(19) => 
                           predigest_product_8_19_port, A(18) => 
                           predigest_product_8_18_port, A(17) => 
                           predigest_product_8_17_port, A(16) => 
                           predigest_product_8_16_port, A(15) => 
                           predigest_product_8_15_port, A(14) => 
                           predigest_product_8_14_port, A(13) => 
                           predigest_product_8_13_port, A(12) => 
                           predigest_product_8_12_port, A(11) => 
                           predigest_product_8_11_port, A(10) => 
                           predigest_product_8_10_port, A(9) => 
                           predigest_product_8_9_port, A(8) => 
                           predigest_product_8_8_port, A(7) => 
                           predigest_product_8_7_port, A(6) => 
                           predigest_product_8_6_port, A(5) => 
                           predigest_product_8_5_port, A(4) => 
                           predigest_product_8_4_port, A(3) => 
                           predigest_product_8_3_port, A(2) => 
                           predigest_product_8_2_port, A(1) => 
                           predigest_product_8_1_port, A(0) => 
                           predigest_product_8_0_port, B(63) => 
                           out_imux_9_63_port, B(62) => out_imux_9_62_port, 
                           B(61) => out_imux_9_61_port, B(60) => 
                           out_imux_9_60_port, B(59) => out_imux_9_59_port, 
                           B(58) => out_imux_9_58_port, B(57) => 
                           out_imux_9_57_port, B(56) => out_imux_9_56_port, 
                           B(55) => out_imux_9_55_port, B(54) => 
                           out_imux_9_54_port, B(53) => out_imux_9_53_port, 
                           B(52) => out_imux_9_52_port, B(51) => 
                           out_imux_9_51_port, B(50) => out_imux_9_50_port, 
                           B(49) => out_imux_9_49_port, B(48) => 
                           out_imux_9_48_port, B(47) => out_imux_9_47_port, 
                           B(46) => out_imux_9_46_port, B(45) => 
                           out_imux_9_45_port, B(44) => out_imux_9_44_port, 
                           B(43) => out_imux_9_43_port, B(42) => 
                           out_imux_9_42_port, B(41) => out_imux_9_41_port, 
                           B(40) => out_imux_9_40_port, B(39) => 
                           out_imux_9_39_port, B(38) => out_imux_9_38_port, 
                           B(37) => out_imux_9_37_port, B(36) => 
                           out_imux_9_36_port, B(35) => out_imux_9_35_port, 
                           B(34) => out_imux_9_34_port, B(33) => 
                           out_imux_9_33_port, B(32) => out_imux_9_32_port, 
                           B(31) => out_imux_9_31_port, B(30) => 
                           out_imux_9_30_port, B(29) => out_imux_9_29_port, 
                           B(28) => out_imux_9_28_port, B(27) => 
                           out_imux_9_27_port, B(26) => out_imux_9_26_port, 
                           B(25) => out_imux_9_25_port, B(24) => 
                           out_imux_9_24_port, B(23) => out_imux_9_23_port, 
                           B(22) => out_imux_9_22_port, B(21) => 
                           out_imux_9_21_port, B(20) => out_imux_9_20_port, 
                           B(19) => out_imux_9_19_port, B(18) => 
                           out_imux_9_18_port, B(17) => out_imux_9_17_port, 
                           B(16) => out_imux_9_16_port, B(15) => 
                           out_imux_9_15_port, B(14) => out_imux_9_14_port, 
                           B(13) => out_imux_9_13_port, B(12) => 
                           out_imux_9_12_port, B(11) => out_imux_9_11_port, 
                           B(10) => out_imux_9_10_port, B(9) => 
                           out_imux_9_9_port, B(8) => out_imux_9_8_port, B(7) 
                           => out_imux_9_7_port, B(6) => out_imux_9_6_port, 
                           B(5) => out_imux_9_5_port, B(4) => out_imux_9_4_port
                           , B(3) => out_imux_9_3_port, B(2) => 
                           out_imux_9_2_port, B(1) => out_imux_9_1_port, B(0) 
                           => out_imux_9_0_port, Ci => X_Logic0_port, S(63) => 
                           predigest_product_9_63_port, S(62) => 
                           predigest_product_9_62_port, S(61) => 
                           predigest_product_9_61_port, S(60) => 
                           predigest_product_9_60_port, S(59) => 
                           predigest_product_9_59_port, S(58) => 
                           predigest_product_9_58_port, S(57) => 
                           predigest_product_9_57_port, S(56) => 
                           predigest_product_9_56_port, S(55) => 
                           predigest_product_9_55_port, S(54) => 
                           predigest_product_9_54_port, S(53) => 
                           predigest_product_9_53_port, S(52) => 
                           predigest_product_9_52_port, S(51) => 
                           predigest_product_9_51_port, S(50) => 
                           predigest_product_9_50_port, S(49) => 
                           predigest_product_9_49_port, S(48) => 
                           predigest_product_9_48_port, S(47) => 
                           predigest_product_9_47_port, S(46) => 
                           predigest_product_9_46_port, S(45) => 
                           predigest_product_9_45_port, S(44) => 
                           predigest_product_9_44_port, S(43) => 
                           predigest_product_9_43_port, S(42) => 
                           predigest_product_9_42_port, S(41) => 
                           predigest_product_9_41_port, S(40) => 
                           predigest_product_9_40_port, S(39) => 
                           predigest_product_9_39_port, S(38) => 
                           predigest_product_9_38_port, S(37) => 
                           predigest_product_9_37_port, S(36) => 
                           predigest_product_9_36_port, S(35) => 
                           predigest_product_9_35_port, S(34) => 
                           predigest_product_9_34_port, S(33) => 
                           predigest_product_9_33_port, S(32) => 
                           predigest_product_9_32_port, S(31) => 
                           predigest_product_9_31_port, S(30) => 
                           predigest_product_9_30_port, S(29) => 
                           predigest_product_9_29_port, S(28) => 
                           predigest_product_9_28_port, S(27) => 
                           predigest_product_9_27_port, S(26) => 
                           predigest_product_9_26_port, S(25) => 
                           predigest_product_9_25_port, S(24) => 
                           predigest_product_9_24_port, S(23) => 
                           predigest_product_9_23_port, S(22) => 
                           predigest_product_9_22_port, S(21) => 
                           predigest_product_9_21_port, S(20) => 
                           predigest_product_9_20_port, S(19) => 
                           predigest_product_9_19_port, S(18) => 
                           predigest_product_9_18_port, S(17) => 
                           predigest_product_9_17_port, S(16) => 
                           predigest_product_9_16_port, S(15) => 
                           predigest_product_9_15_port, S(14) => 
                           predigest_product_9_14_port, S(13) => 
                           predigest_product_9_13_port, S(12) => 
                           predigest_product_9_12_port, S(11) => 
                           predigest_product_9_11_port, S(10) => 
                           predigest_product_9_10_port, S(9) => 
                           predigest_product_9_9_port, S(8) => 
                           predigest_product_9_8_port, S(7) => 
                           predigest_product_9_7_port, S(6) => 
                           predigest_product_9_6_port, S(5) => 
                           predigest_product_9_5_port, S(4) => 
                           predigest_product_9_4_port, S(3) => 
                           predigest_product_9_3_port, S(2) => 
                           predigest_product_9_2_port, S(1) => 
                           predigest_product_9_1_port, S(0) => 
                           predigest_product_9_0_port, Co => n_1100);
   ENC_i_10 : BOOTH_ENCODER_3BIT_10 port map( B(2) => B(21), B(1) => B(20), 
                           B(0) => B(19), ENCODED(2) => 
                           muxs_encoded_signals_10_2_port, ENCODED(1) => 
                           muxs_encoded_signals_10_1_port, ENCODED(0) => 
                           muxs_encoded_signals_10_0_port);
   MUX_i_10 : MUX51_GENERIC_NBIT64_6 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(31), IN1(51) 
                           => A(31), IN1(50) => A(30), IN1(49) => A(29), 
                           IN1(48) => A(28), IN1(47) => A(27), IN1(46) => A(26)
                           , IN1(45) => A(25), IN1(44) => A(24), IN1(43) => 
                           A(23), IN1(42) => A(22), IN1(41) => A(21), IN1(40) 
                           => A(20), IN1(39) => A(19), IN1(38) => A(18), 
                           IN1(37) => A(17), IN1(36) => A(16), IN1(35) => A(15)
                           , IN1(34) => A(14), IN1(33) => A(13), IN1(32) => 
                           A(12), IN1(31) => A(11), IN1(30) => A(10), IN1(29) 
                           => A(9), IN1(28) => A(8), IN1(27) => A(7), IN1(26) 
                           => A(6), IN1(25) => A(5), IN1(24) => A(4), IN1(23) 
                           => A(3), IN1(22) => A(2), IN1(21) => A(1), IN1(20) 
                           => A(0), IN1(19) => X_Logic0_port, IN1(18) => 
                           X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) => 
                           X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) => 
                           X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) => 
                           X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) => 
                           X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) => 
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(63) => negative_a_43_port, 
                           IN2(62) => negative_a_42_port, IN2(61) => 
                           negative_a_41_port, IN2(60) => negative_a_40_port, 
                           IN2(59) => negative_a_39_port, IN2(58) => 
                           negative_a_38_port, IN2(57) => negative_a_37_port, 
                           IN2(56) => negative_a_36_port, IN2(55) => 
                           negative_a_35_port, IN2(54) => negative_a_34_port, 
                           IN2(53) => n37, IN2(52) => n34, IN2(51) => 
                           negative_a_31_port, IN2(50) => negative_a_30_port, 
                           IN2(49) => negative_a_29_port, IN2(48) => 
                           negative_a_28_port, IN2(47) => negative_a_27_port, 
                           IN2(46) => negative_a_26_port, IN2(45) => 
                           negative_a_25_port, IN2(44) => negative_a_24_port, 
                           IN2(43) => negative_a_23_port, IN2(42) => 
                           negative_a_22_port, IN2(41) => negative_a_21_port, 
                           IN2(40) => negative_a_20_port, IN2(39) => 
                           negative_a_19_port, IN2(38) => negative_a_18_port, 
                           IN2(37) => negative_a_17_port, IN2(36) => 
                           negative_a_16_port, IN2(35) => negative_a_15_port, 
                           IN2(34) => negative_a_14_port, IN2(33) => 
                           negative_a_13_port, IN2(32) => negative_a_12_port, 
                           IN2(31) => negative_a_11_port, IN2(30) => 
                           negative_a_10_port, IN2(29) => negative_a_9_port, 
                           IN2(28) => negative_a_8_port, IN2(27) => 
                           negative_a_7_port, IN2(26) => negative_a_6_port, 
                           IN2(25) => negative_a_5_port, IN2(24) => 
                           negative_a_4_port, IN2(23) => negative_a_3_port, 
                           IN2(22) => negative_a_2_port, IN2(21) => 
                           negative_a_1_port, IN2(20) => negative_a_0_port, 
                           IN2(19) => X_Logic0_port, IN2(18) => X_Logic0_port, 
                           IN2(17) => X_Logic0_port, IN2(16) => X_Logic0_port, 
                           IN2(15) => X_Logic0_port, IN2(14) => X_Logic0_port, 
                           IN2(13) => X_Logic0_port, IN2(12) => X_Logic0_port, 
                           IN2(11) => X_Logic0_port, IN2(10) => X_Logic0_port, 
                           IN2(9) => X_Logic0_port, IN2(8) => X_Logic0_port, 
                           IN2(7) => X_Logic0_port, IN2(6) => X_Logic0_port, 
                           IN2(5) => X_Logic0_port, IN2(4) => X_Logic0_port, 
                           IN2(3) => X_Logic0_port, IN2(2) => X_Logic0_port, 
                           IN2(1) => X_Logic0_port, IN2(0) => X_Logic0_port, 
                           IN3(63) => A(31), IN3(62) => A(31), IN3(61) => A(31)
                           , IN3(60) => A(31), IN3(59) => A(31), IN3(58) => 
                           A(31), IN3(57) => A(31), IN3(56) => A(31), IN3(55) 
                           => A(31), IN3(54) => A(31), IN3(53) => A(31), 
                           IN3(52) => A(31), IN3(51) => A(30), IN3(50) => A(29)
                           , IN3(49) => A(28), IN3(48) => A(27), IN3(47) => 
                           A(26), IN3(46) => A(25), IN3(45) => A(24), IN3(44) 
                           => A(23), IN3(43) => A(22), IN3(42) => A(21), 
                           IN3(41) => A(20), IN3(40) => A(19), IN3(39) => A(18)
                           , IN3(38) => A(17), IN3(37) => A(16), IN3(36) => 
                           A(15), IN3(35) => A(14), IN3(34) => A(13), IN3(33) 
                           => A(12), IN3(32) => A(11), IN3(31) => A(10), 
                           IN3(30) => A(9), IN3(29) => A(8), IN3(28) => A(7), 
                           IN3(27) => A(6), IN3(26) => A(5), IN3(25) => A(4), 
                           IN3(24) => A(3), IN3(23) => A(2), IN3(22) => A(1), 
                           IN3(21) => A(0), IN3(20) => X_Logic0_port, IN3(19) 
                           => X_Logic0_port, IN3(18) => X_Logic0_port, IN3(17) 
                           => X_Logic0_port, IN3(16) => X_Logic0_port, IN3(15) 
                           => X_Logic0_port, IN3(14) => X_Logic0_port, IN3(13) 
                           => X_Logic0_port, IN3(12) => X_Logic0_port, IN3(11) 
                           => X_Logic0_port, IN3(10) => X_Logic0_port, IN3(9) 
                           => X_Logic0_port, IN3(8) => X_Logic0_port, IN3(7) =>
                           X_Logic0_port, IN3(6) => X_Logic0_port, IN3(5) => 
                           X_Logic0_port, IN3(4) => X_Logic0_port, IN3(3) => 
                           X_Logic0_port, IN3(2) => X_Logic0_port, IN3(1) => 
                           X_Logic0_port, IN3(0) => X_Logic0_port, IN4(63) => 
                           negative_a_42_port, IN4(62) => negative_a_41_port, 
                           IN4(61) => negative_a_40_port, IN4(60) => 
                           negative_a_39_port, IN4(59) => negative_a_38_port, 
                           IN4(58) => negative_a_37_port, IN4(57) => 
                           negative_a_36_port, IN4(56) => negative_a_35_port, 
                           IN4(55) => negative_a_34_port, IN4(54) => n37, 
                           IN4(53) => n34, IN4(52) => negative_a_31_port, 
                           IN4(51) => negative_a_30_port, IN4(50) => 
                           negative_a_29_port, IN4(49) => negative_a_28_port, 
                           IN4(48) => negative_a_27_port, IN4(47) => 
                           negative_a_26_port, IN4(46) => negative_a_25_port, 
                           IN4(45) => negative_a_24_port, IN4(44) => 
                           negative_a_23_port, IN4(43) => negative_a_22_port, 
                           IN4(42) => negative_a_21_port, IN4(41) => 
                           negative_a_20_port, IN4(40) => negative_a_19_port, 
                           IN4(39) => negative_a_18_port, IN4(38) => 
                           negative_a_17_port, IN4(37) => negative_a_16_port, 
                           IN4(36) => negative_a_15_port, IN4(35) => 
                           negative_a_14_port, IN4(34) => negative_a_13_port, 
                           IN4(33) => negative_a_12_port, IN4(32) => 
                           negative_a_11_port, IN4(31) => negative_a_10_port, 
                           IN4(30) => negative_a_9_port, IN4(29) => 
                           negative_a_8_port, IN4(28) => negative_a_7_port, 
                           IN4(27) => negative_a_6_port, IN4(26) => 
                           negative_a_5_port, IN4(25) => negative_a_4_port, 
                           IN4(24) => negative_a_3_port, IN4(23) => 
                           negative_a_2_port, IN4(22) => negative_a_1_port, 
                           IN4(21) => negative_a_0_port, IN4(20) => 
                           X_Logic0_port, IN4(19) => X_Logic0_port, IN4(18) => 
                           X_Logic0_port, IN4(17) => X_Logic0_port, IN4(16) => 
                           X_Logic0_port, IN4(15) => X_Logic0_port, IN4(14) => 
                           X_Logic0_port, IN4(13) => X_Logic0_port, IN4(12) => 
                           X_Logic0_port, IN4(11) => X_Logic0_port, IN4(10) => 
                           X_Logic0_port, IN4(9) => X_Logic0_port, IN4(8) => 
                           X_Logic0_port, IN4(7) => X_Logic0_port, IN4(6) => 
                           X_Logic0_port, IN4(5) => X_Logic0_port, IN4(4) => 
                           X_Logic0_port, IN4(3) => X_Logic0_port, IN4(2) => 
                           X_Logic0_port, IN4(1) => X_Logic0_port, IN4(0) => 
                           X_Logic0_port, S(2) => 
                           muxs_encoded_signals_10_2_port, S(1) => 
                           muxs_encoded_signals_10_1_port, S(0) => 
                           muxs_encoded_signals_10_0_port, O(63) => 
                           out_imux_10_63_port, O(62) => out_imux_10_62_port, 
                           O(61) => out_imux_10_61_port, O(60) => 
                           out_imux_10_60_port, O(59) => out_imux_10_59_port, 
                           O(58) => out_imux_10_58_port, O(57) => 
                           out_imux_10_57_port, O(56) => out_imux_10_56_port, 
                           O(55) => out_imux_10_55_port, O(54) => 
                           out_imux_10_54_port, O(53) => out_imux_10_53_port, 
                           O(52) => out_imux_10_52_port, O(51) => 
                           out_imux_10_51_port, O(50) => out_imux_10_50_port, 
                           O(49) => out_imux_10_49_port, O(48) => 
                           out_imux_10_48_port, O(47) => out_imux_10_47_port, 
                           O(46) => out_imux_10_46_port, O(45) => 
                           out_imux_10_45_port, O(44) => out_imux_10_44_port, 
                           O(43) => out_imux_10_43_port, O(42) => 
                           out_imux_10_42_port, O(41) => out_imux_10_41_port, 
                           O(40) => out_imux_10_40_port, O(39) => 
                           out_imux_10_39_port, O(38) => out_imux_10_38_port, 
                           O(37) => out_imux_10_37_port, O(36) => 
                           out_imux_10_36_port, O(35) => out_imux_10_35_port, 
                           O(34) => out_imux_10_34_port, O(33) => 
                           out_imux_10_33_port, O(32) => out_imux_10_32_port, 
                           O(31) => out_imux_10_31_port, O(30) => 
                           out_imux_10_30_port, O(29) => out_imux_10_29_port, 
                           O(28) => out_imux_10_28_port, O(27) => 
                           out_imux_10_27_port, O(26) => out_imux_10_26_port, 
                           O(25) => out_imux_10_25_port, O(24) => 
                           out_imux_10_24_port, O(23) => out_imux_10_23_port, 
                           O(22) => out_imux_10_22_port, O(21) => 
                           out_imux_10_21_port, O(20) => out_imux_10_20_port, 
                           O(19) => out_imux_10_19_port, O(18) => 
                           out_imux_10_18_port, O(17) => out_imux_10_17_port, 
                           O(16) => out_imux_10_16_port, O(15) => 
                           out_imux_10_15_port, O(14) => out_imux_10_14_port, 
                           O(13) => out_imux_10_13_port, O(12) => 
                           out_imux_10_12_port, O(11) => out_imux_10_11_port, 
                           O(10) => out_imux_10_10_port, O(9) => 
                           out_imux_10_9_port, O(8) => out_imux_10_8_port, O(7)
                           => out_imux_10_7_port, O(6) => out_imux_10_6_port, 
                           O(5) => out_imux_10_5_port, O(4) => 
                           out_imux_10_4_port, O(3) => out_imux_10_3_port, O(2)
                           => out_imux_10_2_port, O(1) => out_imux_10_1_port, 
                           O(0) => out_imux_10_0_port);
   ADD64_i_10 : RCA_GENERIC_NBIT64_6 port map( A(63) => 
                           predigest_product_9_63_port, A(62) => 
                           predigest_product_9_62_port, A(61) => 
                           predigest_product_9_61_port, A(60) => 
                           predigest_product_9_60_port, A(59) => 
                           predigest_product_9_59_port, A(58) => 
                           predigest_product_9_58_port, A(57) => 
                           predigest_product_9_57_port, A(56) => 
                           predigest_product_9_56_port, A(55) => 
                           predigest_product_9_55_port, A(54) => 
                           predigest_product_9_54_port, A(53) => 
                           predigest_product_9_53_port, A(52) => 
                           predigest_product_9_52_port, A(51) => 
                           predigest_product_9_51_port, A(50) => 
                           predigest_product_9_50_port, A(49) => 
                           predigest_product_9_49_port, A(48) => 
                           predigest_product_9_48_port, A(47) => 
                           predigest_product_9_47_port, A(46) => 
                           predigest_product_9_46_port, A(45) => 
                           predigest_product_9_45_port, A(44) => 
                           predigest_product_9_44_port, A(43) => 
                           predigest_product_9_43_port, A(42) => 
                           predigest_product_9_42_port, A(41) => 
                           predigest_product_9_41_port, A(40) => 
                           predigest_product_9_40_port, A(39) => 
                           predigest_product_9_39_port, A(38) => 
                           predigest_product_9_38_port, A(37) => 
                           predigest_product_9_37_port, A(36) => 
                           predigest_product_9_36_port, A(35) => 
                           predigest_product_9_35_port, A(34) => 
                           predigest_product_9_34_port, A(33) => 
                           predigest_product_9_33_port, A(32) => 
                           predigest_product_9_32_port, A(31) => 
                           predigest_product_9_31_port, A(30) => 
                           predigest_product_9_30_port, A(29) => 
                           predigest_product_9_29_port, A(28) => 
                           predigest_product_9_28_port, A(27) => 
                           predigest_product_9_27_port, A(26) => 
                           predigest_product_9_26_port, A(25) => 
                           predigest_product_9_25_port, A(24) => 
                           predigest_product_9_24_port, A(23) => 
                           predigest_product_9_23_port, A(22) => 
                           predigest_product_9_22_port, A(21) => 
                           predigest_product_9_21_port, A(20) => 
                           predigest_product_9_20_port, A(19) => 
                           predigest_product_9_19_port, A(18) => 
                           predigest_product_9_18_port, A(17) => 
                           predigest_product_9_17_port, A(16) => 
                           predigest_product_9_16_port, A(15) => 
                           predigest_product_9_15_port, A(14) => 
                           predigest_product_9_14_port, A(13) => 
                           predigest_product_9_13_port, A(12) => 
                           predigest_product_9_12_port, A(11) => 
                           predigest_product_9_11_port, A(10) => 
                           predigest_product_9_10_port, A(9) => 
                           predigest_product_9_9_port, A(8) => 
                           predigest_product_9_8_port, A(7) => 
                           predigest_product_9_7_port, A(6) => 
                           predigest_product_9_6_port, A(5) => 
                           predigest_product_9_5_port, A(4) => 
                           predigest_product_9_4_port, A(3) => 
                           predigest_product_9_3_port, A(2) => 
                           predigest_product_9_2_port, A(1) => 
                           predigest_product_9_1_port, A(0) => 
                           predigest_product_9_0_port, B(63) => 
                           out_imux_10_63_port, B(62) => out_imux_10_62_port, 
                           B(61) => out_imux_10_61_port, B(60) => 
                           out_imux_10_60_port, B(59) => out_imux_10_59_port, 
                           B(58) => out_imux_10_58_port, B(57) => 
                           out_imux_10_57_port, B(56) => out_imux_10_56_port, 
                           B(55) => out_imux_10_55_port, B(54) => 
                           out_imux_10_54_port, B(53) => out_imux_10_53_port, 
                           B(52) => out_imux_10_52_port, B(51) => 
                           out_imux_10_51_port, B(50) => out_imux_10_50_port, 
                           B(49) => out_imux_10_49_port, B(48) => 
                           out_imux_10_48_port, B(47) => out_imux_10_47_port, 
                           B(46) => out_imux_10_46_port, B(45) => 
                           out_imux_10_45_port, B(44) => out_imux_10_44_port, 
                           B(43) => out_imux_10_43_port, B(42) => 
                           out_imux_10_42_port, B(41) => out_imux_10_41_port, 
                           B(40) => out_imux_10_40_port, B(39) => 
                           out_imux_10_39_port, B(38) => out_imux_10_38_port, 
                           B(37) => out_imux_10_37_port, B(36) => 
                           out_imux_10_36_port, B(35) => out_imux_10_35_port, 
                           B(34) => out_imux_10_34_port, B(33) => 
                           out_imux_10_33_port, B(32) => out_imux_10_32_port, 
                           B(31) => out_imux_10_31_port, B(30) => 
                           out_imux_10_30_port, B(29) => out_imux_10_29_port, 
                           B(28) => out_imux_10_28_port, B(27) => 
                           out_imux_10_27_port, B(26) => out_imux_10_26_port, 
                           B(25) => out_imux_10_25_port, B(24) => 
                           out_imux_10_24_port, B(23) => out_imux_10_23_port, 
                           B(22) => out_imux_10_22_port, B(21) => 
                           out_imux_10_21_port, B(20) => out_imux_10_20_port, 
                           B(19) => out_imux_10_19_port, B(18) => 
                           out_imux_10_18_port, B(17) => out_imux_10_17_port, 
                           B(16) => out_imux_10_16_port, B(15) => 
                           out_imux_10_15_port, B(14) => out_imux_10_14_port, 
                           B(13) => out_imux_10_13_port, B(12) => 
                           out_imux_10_12_port, B(11) => out_imux_10_11_port, 
                           B(10) => out_imux_10_10_port, B(9) => 
                           out_imux_10_9_port, B(8) => out_imux_10_8_port, B(7)
                           => out_imux_10_7_port, B(6) => out_imux_10_6_port, 
                           B(5) => out_imux_10_5_port, B(4) => 
                           out_imux_10_4_port, B(3) => out_imux_10_3_port, B(2)
                           => out_imux_10_2_port, B(1) => out_imux_10_1_port, 
                           B(0) => out_imux_10_0_port, Ci => X_Logic0_port, 
                           S(63) => predigest_product_10_63_port, S(62) => 
                           predigest_product_10_62_port, S(61) => 
                           predigest_product_10_61_port, S(60) => 
                           predigest_product_10_60_port, S(59) => 
                           predigest_product_10_59_port, S(58) => 
                           predigest_product_10_58_port, S(57) => 
                           predigest_product_10_57_port, S(56) => 
                           predigest_product_10_56_port, S(55) => 
                           predigest_product_10_55_port, S(54) => 
                           predigest_product_10_54_port, S(53) => 
                           predigest_product_10_53_port, S(52) => 
                           predigest_product_10_52_port, S(51) => 
                           predigest_product_10_51_port, S(50) => 
                           predigest_product_10_50_port, S(49) => 
                           predigest_product_10_49_port, S(48) => 
                           predigest_product_10_48_port, S(47) => 
                           predigest_product_10_47_port, S(46) => 
                           predigest_product_10_46_port, S(45) => 
                           predigest_product_10_45_port, S(44) => 
                           predigest_product_10_44_port, S(43) => 
                           predigest_product_10_43_port, S(42) => 
                           predigest_product_10_42_port, S(41) => 
                           predigest_product_10_41_port, S(40) => 
                           predigest_product_10_40_port, S(39) => 
                           predigest_product_10_39_port, S(38) => 
                           predigest_product_10_38_port, S(37) => 
                           predigest_product_10_37_port, S(36) => 
                           predigest_product_10_36_port, S(35) => 
                           predigest_product_10_35_port, S(34) => 
                           predigest_product_10_34_port, S(33) => 
                           predigest_product_10_33_port, S(32) => 
                           predigest_product_10_32_port, S(31) => 
                           predigest_product_10_31_port, S(30) => 
                           predigest_product_10_30_port, S(29) => 
                           predigest_product_10_29_port, S(28) => 
                           predigest_product_10_28_port, S(27) => 
                           predigest_product_10_27_port, S(26) => 
                           predigest_product_10_26_port, S(25) => 
                           predigest_product_10_25_port, S(24) => 
                           predigest_product_10_24_port, S(23) => 
                           predigest_product_10_23_port, S(22) => 
                           predigest_product_10_22_port, S(21) => 
                           predigest_product_10_21_port, S(20) => 
                           predigest_product_10_20_port, S(19) => 
                           predigest_product_10_19_port, S(18) => 
                           predigest_product_10_18_port, S(17) => 
                           predigest_product_10_17_port, S(16) => 
                           predigest_product_10_16_port, S(15) => 
                           predigest_product_10_15_port, S(14) => 
                           predigest_product_10_14_port, S(13) => 
                           predigest_product_10_13_port, S(12) => 
                           predigest_product_10_12_port, S(11) => 
                           predigest_product_10_11_port, S(10) => 
                           predigest_product_10_10_port, S(9) => 
                           predigest_product_10_9_port, S(8) => 
                           predigest_product_10_8_port, S(7) => 
                           predigest_product_10_7_port, S(6) => 
                           predigest_product_10_6_port, S(5) => 
                           predigest_product_10_5_port, S(4) => 
                           predigest_product_10_4_port, S(3) => 
                           predigest_product_10_3_port, S(2) => 
                           predigest_product_10_2_port, S(1) => 
                           predigest_product_10_1_port, S(0) => 
                           predigest_product_10_0_port, Co => n_1101);
   ENC_i_11 : BOOTH_ENCODER_3BIT_9 port map( B(2) => B(23), B(1) => B(22), B(0)
                           => B(21), ENCODED(2) => 
                           muxs_encoded_signals_11_2_port, ENCODED(1) => 
                           muxs_encoded_signals_11_1_port, ENCODED(0) => 
                           muxs_encoded_signals_11_0_port);
   MUX_i_11 : MUX51_GENERIC_NBIT64_5 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(31), IN1(53) => A(31), IN1(52) => A(30), IN1(51) 
                           => A(29), IN1(50) => A(28), IN1(49) => A(27), 
                           IN1(48) => A(26), IN1(47) => A(25), IN1(46) => A(24)
                           , IN1(45) => A(23), IN1(44) => A(22), IN1(43) => 
                           A(21), IN1(42) => A(20), IN1(41) => A(19), IN1(40) 
                           => A(18), IN1(39) => A(17), IN1(38) => A(16), 
                           IN1(37) => A(15), IN1(36) => A(14), IN1(35) => A(13)
                           , IN1(34) => A(12), IN1(33) => A(11), IN1(32) => 
                           A(10), IN1(31) => A(9), IN1(30) => A(8), IN1(29) => 
                           A(7), IN1(28) => A(6), IN1(27) => A(5), IN1(26) => 
                           A(4), IN1(25) => A(3), IN1(24) => A(2), IN1(23) => 
                           A(1), IN1(22) => A(0), IN1(21) => X_Logic0_port, 
                           IN1(20) => X_Logic0_port, IN1(19) => X_Logic0_port, 
                           IN1(18) => X_Logic0_port, IN1(17) => X_Logic0_port, 
                           IN1(16) => X_Logic0_port, IN1(15) => X_Logic0_port, 
                           IN1(14) => X_Logic0_port, IN1(13) => X_Logic0_port, 
                           IN1(12) => X_Logic0_port, IN1(11) => X_Logic0_port, 
                           IN1(10) => X_Logic0_port, IN1(9) => X_Logic0_port, 
                           IN1(8) => X_Logic0_port, IN1(7) => X_Logic0_port, 
                           IN1(6) => X_Logic0_port, IN1(5) => X_Logic0_port, 
                           IN1(4) => X_Logic0_port, IN1(3) => X_Logic0_port, 
                           IN1(2) => X_Logic0_port, IN1(1) => X_Logic0_port, 
                           IN1(0) => X_Logic0_port, IN2(63) => 
                           negative_a_41_port, IN2(62) => negative_a_40_port, 
                           IN2(61) => negative_a_39_port, IN2(60) => 
                           negative_a_38_port, IN2(59) => negative_a_37_port, 
                           IN2(58) => negative_a_36_port, IN2(57) => 
                           negative_a_35_port, IN2(56) => negative_a_34_port, 
                           IN2(55) => n37, IN2(54) => n34, IN2(53) => 
                           negative_a_31_port, IN2(52) => negative_a_30_port, 
                           IN2(51) => negative_a_29_port, IN2(50) => 
                           negative_a_28_port, IN2(49) => negative_a_27_port, 
                           IN2(48) => negative_a_26_port, IN2(47) => 
                           negative_a_25_port, IN2(46) => negative_a_24_port, 
                           IN2(45) => negative_a_23_port, IN2(44) => 
                           negative_a_22_port, IN2(43) => negative_a_21_port, 
                           IN2(42) => negative_a_20_port, IN2(41) => 
                           negative_a_19_port, IN2(40) => negative_a_18_port, 
                           IN2(39) => negative_a_17_port, IN2(38) => 
                           negative_a_16_port, IN2(37) => negative_a_15_port, 
                           IN2(36) => negative_a_14_port, IN2(35) => 
                           negative_a_13_port, IN2(34) => negative_a_12_port, 
                           IN2(33) => negative_a_11_port, IN2(32) => 
                           negative_a_10_port, IN2(31) => negative_a_9_port, 
                           IN2(30) => negative_a_8_port, IN2(29) => 
                           negative_a_7_port, IN2(28) => negative_a_6_port, 
                           IN2(27) => negative_a_5_port, IN2(26) => 
                           negative_a_4_port, IN2(25) => negative_a_3_port, 
                           IN2(24) => negative_a_2_port, IN2(23) => 
                           negative_a_1_port, IN2(22) => negative_a_0_port, 
                           IN2(21) => X_Logic0_port, IN2(20) => X_Logic0_port, 
                           IN2(19) => X_Logic0_port, IN2(18) => X_Logic0_port, 
                           IN2(17) => X_Logic0_port, IN2(16) => X_Logic0_port, 
                           IN2(15) => X_Logic0_port, IN2(14) => X_Logic0_port, 
                           IN2(13) => X_Logic0_port, IN2(12) => X_Logic0_port, 
                           IN2(11) => X_Logic0_port, IN2(10) => X_Logic0_port, 
                           IN2(9) => X_Logic0_port, IN2(8) => X_Logic0_port, 
                           IN2(7) => X_Logic0_port, IN2(6) => X_Logic0_port, 
                           IN2(5) => X_Logic0_port, IN2(4) => X_Logic0_port, 
                           IN2(3) => X_Logic0_port, IN2(2) => X_Logic0_port, 
                           IN2(1) => X_Logic0_port, IN2(0) => X_Logic0_port, 
                           IN3(63) => A(31), IN3(62) => A(31), IN3(61) => A(31)
                           , IN3(60) => A(31), IN3(59) => A(31), IN3(58) => 
                           A(31), IN3(57) => A(31), IN3(56) => A(31), IN3(55) 
                           => A(31), IN3(54) => A(31), IN3(53) => A(30), 
                           IN3(52) => A(29), IN3(51) => A(28), IN3(50) => A(27)
                           , IN3(49) => A(26), IN3(48) => A(25), IN3(47) => 
                           A(24), IN3(46) => A(23), IN3(45) => A(22), IN3(44) 
                           => A(21), IN3(43) => A(20), IN3(42) => A(19), 
                           IN3(41) => A(18), IN3(40) => A(17), IN3(39) => A(16)
                           , IN3(38) => A(15), IN3(37) => A(14), IN3(36) => 
                           A(13), IN3(35) => A(12), IN3(34) => A(11), IN3(33) 
                           => A(10), IN3(32) => A(9), IN3(31) => A(8), IN3(30) 
                           => A(7), IN3(29) => A(6), IN3(28) => A(5), IN3(27) 
                           => A(4), IN3(26) => A(3), IN3(25) => A(2), IN3(24) 
                           => A(1), IN3(23) => A(0), IN3(22) => X_Logic0_port, 
                           IN3(21) => X_Logic0_port, IN3(20) => X_Logic0_port, 
                           IN3(19) => X_Logic0_port, IN3(18) => X_Logic0_port, 
                           IN3(17) => X_Logic0_port, IN3(16) => X_Logic0_port, 
                           IN3(15) => X_Logic0_port, IN3(14) => X_Logic0_port, 
                           IN3(13) => X_Logic0_port, IN3(12) => X_Logic0_port, 
                           IN3(11) => X_Logic0_port, IN3(10) => X_Logic0_port, 
                           IN3(9) => X_Logic0_port, IN3(8) => X_Logic0_port, 
                           IN3(7) => X_Logic0_port, IN3(6) => X_Logic0_port, 
                           IN3(5) => X_Logic0_port, IN3(4) => X_Logic0_port, 
                           IN3(3) => X_Logic0_port, IN3(2) => X_Logic0_port, 
                           IN3(1) => X_Logic0_port, IN3(0) => X_Logic0_port, 
                           IN4(63) => negative_a_40_port, IN4(62) => 
                           negative_a_39_port, IN4(61) => negative_a_38_port, 
                           IN4(60) => negative_a_37_port, IN4(59) => 
                           negative_a_36_port, IN4(58) => negative_a_35_port, 
                           IN4(57) => negative_a_34_port, IN4(56) => n37, 
                           IN4(55) => n34, IN4(54) => negative_a_31_port, 
                           IN4(53) => negative_a_30_port, IN4(52) => 
                           negative_a_29_port, IN4(51) => negative_a_28_port, 
                           IN4(50) => negative_a_27_port, IN4(49) => 
                           negative_a_26_port, IN4(48) => negative_a_25_port, 
                           IN4(47) => negative_a_24_port, IN4(46) => 
                           negative_a_23_port, IN4(45) => negative_a_22_port, 
                           IN4(44) => negative_a_21_port, IN4(43) => 
                           negative_a_20_port, IN4(42) => negative_a_19_port, 
                           IN4(41) => negative_a_18_port, IN4(40) => 
                           negative_a_17_port, IN4(39) => negative_a_16_port, 
                           IN4(38) => negative_a_15_port, IN4(37) => 
                           negative_a_14_port, IN4(36) => negative_a_13_port, 
                           IN4(35) => negative_a_12_port, IN4(34) => 
                           negative_a_11_port, IN4(33) => negative_a_10_port, 
                           IN4(32) => negative_a_9_port, IN4(31) => 
                           negative_a_8_port, IN4(30) => negative_a_7_port, 
                           IN4(29) => negative_a_6_port, IN4(28) => 
                           negative_a_5_port, IN4(27) => negative_a_4_port, 
                           IN4(26) => negative_a_3_port, IN4(25) => 
                           negative_a_2_port, IN4(24) => negative_a_1_port, 
                           IN4(23) => negative_a_0_port, IN4(22) => 
                           X_Logic0_port, IN4(21) => X_Logic0_port, IN4(20) => 
                           X_Logic0_port, IN4(19) => X_Logic0_port, IN4(18) => 
                           X_Logic0_port, IN4(17) => X_Logic0_port, IN4(16) => 
                           X_Logic0_port, IN4(15) => X_Logic0_port, IN4(14) => 
                           X_Logic0_port, IN4(13) => X_Logic0_port, IN4(12) => 
                           X_Logic0_port, IN4(11) => X_Logic0_port, IN4(10) => 
                           X_Logic0_port, IN4(9) => X_Logic0_port, IN4(8) => 
                           X_Logic0_port, IN4(7) => X_Logic0_port, IN4(6) => 
                           X_Logic0_port, IN4(5) => X_Logic0_port, IN4(4) => 
                           X_Logic0_port, IN4(3) => X_Logic0_port, IN4(2) => 
                           X_Logic0_port, IN4(1) => X_Logic0_port, IN4(0) => 
                           X_Logic0_port, S(2) => 
                           muxs_encoded_signals_11_2_port, S(1) => 
                           muxs_encoded_signals_11_1_port, S(0) => 
                           muxs_encoded_signals_11_0_port, O(63) => 
                           out_imux_11_63_port, O(62) => out_imux_11_62_port, 
                           O(61) => out_imux_11_61_port, O(60) => 
                           out_imux_11_60_port, O(59) => out_imux_11_59_port, 
                           O(58) => out_imux_11_58_port, O(57) => 
                           out_imux_11_57_port, O(56) => out_imux_11_56_port, 
                           O(55) => out_imux_11_55_port, O(54) => 
                           out_imux_11_54_port, O(53) => out_imux_11_53_port, 
                           O(52) => out_imux_11_52_port, O(51) => 
                           out_imux_11_51_port, O(50) => out_imux_11_50_port, 
                           O(49) => out_imux_11_49_port, O(48) => 
                           out_imux_11_48_port, O(47) => out_imux_11_47_port, 
                           O(46) => out_imux_11_46_port, O(45) => 
                           out_imux_11_45_port, O(44) => out_imux_11_44_port, 
                           O(43) => out_imux_11_43_port, O(42) => 
                           out_imux_11_42_port, O(41) => out_imux_11_41_port, 
                           O(40) => out_imux_11_40_port, O(39) => 
                           out_imux_11_39_port, O(38) => out_imux_11_38_port, 
                           O(37) => out_imux_11_37_port, O(36) => 
                           out_imux_11_36_port, O(35) => out_imux_11_35_port, 
                           O(34) => out_imux_11_34_port, O(33) => 
                           out_imux_11_33_port, O(32) => out_imux_11_32_port, 
                           O(31) => out_imux_11_31_port, O(30) => 
                           out_imux_11_30_port, O(29) => out_imux_11_29_port, 
                           O(28) => out_imux_11_28_port, O(27) => 
                           out_imux_11_27_port, O(26) => out_imux_11_26_port, 
                           O(25) => out_imux_11_25_port, O(24) => 
                           out_imux_11_24_port, O(23) => out_imux_11_23_port, 
                           O(22) => out_imux_11_22_port, O(21) => 
                           out_imux_11_21_port, O(20) => out_imux_11_20_port, 
                           O(19) => out_imux_11_19_port, O(18) => 
                           out_imux_11_18_port, O(17) => out_imux_11_17_port, 
                           O(16) => out_imux_11_16_port, O(15) => 
                           out_imux_11_15_port, O(14) => out_imux_11_14_port, 
                           O(13) => out_imux_11_13_port, O(12) => 
                           out_imux_11_12_port, O(11) => out_imux_11_11_port, 
                           O(10) => out_imux_11_10_port, O(9) => 
                           out_imux_11_9_port, O(8) => out_imux_11_8_port, O(7)
                           => out_imux_11_7_port, O(6) => out_imux_11_6_port, 
                           O(5) => out_imux_11_5_port, O(4) => 
                           out_imux_11_4_port, O(3) => out_imux_11_3_port, O(2)
                           => out_imux_11_2_port, O(1) => out_imux_11_1_port, 
                           O(0) => out_imux_11_0_port);
   ADD64_i_11 : RCA_GENERIC_NBIT64_5 port map( A(63) => 
                           predigest_product_10_63_port, A(62) => 
                           predigest_product_10_62_port, A(61) => 
                           predigest_product_10_61_port, A(60) => 
                           predigest_product_10_60_port, A(59) => 
                           predigest_product_10_59_port, A(58) => 
                           predigest_product_10_58_port, A(57) => 
                           predigest_product_10_57_port, A(56) => 
                           predigest_product_10_56_port, A(55) => 
                           predigest_product_10_55_port, A(54) => 
                           predigest_product_10_54_port, A(53) => 
                           predigest_product_10_53_port, A(52) => 
                           predigest_product_10_52_port, A(51) => 
                           predigest_product_10_51_port, A(50) => 
                           predigest_product_10_50_port, A(49) => 
                           predigest_product_10_49_port, A(48) => 
                           predigest_product_10_48_port, A(47) => 
                           predigest_product_10_47_port, A(46) => 
                           predigest_product_10_46_port, A(45) => 
                           predigest_product_10_45_port, A(44) => 
                           predigest_product_10_44_port, A(43) => 
                           predigest_product_10_43_port, A(42) => 
                           predigest_product_10_42_port, A(41) => 
                           predigest_product_10_41_port, A(40) => 
                           predigest_product_10_40_port, A(39) => 
                           predigest_product_10_39_port, A(38) => 
                           predigest_product_10_38_port, A(37) => 
                           predigest_product_10_37_port, A(36) => 
                           predigest_product_10_36_port, A(35) => 
                           predigest_product_10_35_port, A(34) => 
                           predigest_product_10_34_port, A(33) => 
                           predigest_product_10_33_port, A(32) => 
                           predigest_product_10_32_port, A(31) => 
                           predigest_product_10_31_port, A(30) => 
                           predigest_product_10_30_port, A(29) => 
                           predigest_product_10_29_port, A(28) => 
                           predigest_product_10_28_port, A(27) => 
                           predigest_product_10_27_port, A(26) => 
                           predigest_product_10_26_port, A(25) => 
                           predigest_product_10_25_port, A(24) => 
                           predigest_product_10_24_port, A(23) => 
                           predigest_product_10_23_port, A(22) => 
                           predigest_product_10_22_port, A(21) => 
                           predigest_product_10_21_port, A(20) => 
                           predigest_product_10_20_port, A(19) => 
                           predigest_product_10_19_port, A(18) => 
                           predigest_product_10_18_port, A(17) => 
                           predigest_product_10_17_port, A(16) => 
                           predigest_product_10_16_port, A(15) => 
                           predigest_product_10_15_port, A(14) => 
                           predigest_product_10_14_port, A(13) => 
                           predigest_product_10_13_port, A(12) => 
                           predigest_product_10_12_port, A(11) => 
                           predigest_product_10_11_port, A(10) => 
                           predigest_product_10_10_port, A(9) => 
                           predigest_product_10_9_port, A(8) => 
                           predigest_product_10_8_port, A(7) => 
                           predigest_product_10_7_port, A(6) => 
                           predigest_product_10_6_port, A(5) => 
                           predigest_product_10_5_port, A(4) => 
                           predigest_product_10_4_port, A(3) => 
                           predigest_product_10_3_port, A(2) => 
                           predigest_product_10_2_port, A(1) => 
                           predigest_product_10_1_port, A(0) => 
                           predigest_product_10_0_port, B(63) => 
                           out_imux_11_63_port, B(62) => out_imux_11_62_port, 
                           B(61) => out_imux_11_61_port, B(60) => 
                           out_imux_11_60_port, B(59) => out_imux_11_59_port, 
                           B(58) => out_imux_11_58_port, B(57) => 
                           out_imux_11_57_port, B(56) => out_imux_11_56_port, 
                           B(55) => out_imux_11_55_port, B(54) => 
                           out_imux_11_54_port, B(53) => out_imux_11_53_port, 
                           B(52) => out_imux_11_52_port, B(51) => 
                           out_imux_11_51_port, B(50) => out_imux_11_50_port, 
                           B(49) => out_imux_11_49_port, B(48) => 
                           out_imux_11_48_port, B(47) => out_imux_11_47_port, 
                           B(46) => out_imux_11_46_port, B(45) => 
                           out_imux_11_45_port, B(44) => out_imux_11_44_port, 
                           B(43) => out_imux_11_43_port, B(42) => 
                           out_imux_11_42_port, B(41) => out_imux_11_41_port, 
                           B(40) => out_imux_11_40_port, B(39) => 
                           out_imux_11_39_port, B(38) => out_imux_11_38_port, 
                           B(37) => out_imux_11_37_port, B(36) => 
                           out_imux_11_36_port, B(35) => out_imux_11_35_port, 
                           B(34) => out_imux_11_34_port, B(33) => 
                           out_imux_11_33_port, B(32) => out_imux_11_32_port, 
                           B(31) => out_imux_11_31_port, B(30) => 
                           out_imux_11_30_port, B(29) => out_imux_11_29_port, 
                           B(28) => out_imux_11_28_port, B(27) => 
                           out_imux_11_27_port, B(26) => out_imux_11_26_port, 
                           B(25) => out_imux_11_25_port, B(24) => 
                           out_imux_11_24_port, B(23) => out_imux_11_23_port, 
                           B(22) => out_imux_11_22_port, B(21) => 
                           out_imux_11_21_port, B(20) => out_imux_11_20_port, 
                           B(19) => out_imux_11_19_port, B(18) => 
                           out_imux_11_18_port, B(17) => out_imux_11_17_port, 
                           B(16) => out_imux_11_16_port, B(15) => 
                           out_imux_11_15_port, B(14) => out_imux_11_14_port, 
                           B(13) => out_imux_11_13_port, B(12) => 
                           out_imux_11_12_port, B(11) => out_imux_11_11_port, 
                           B(10) => out_imux_11_10_port, B(9) => 
                           out_imux_11_9_port, B(8) => out_imux_11_8_port, B(7)
                           => out_imux_11_7_port, B(6) => out_imux_11_6_port, 
                           B(5) => out_imux_11_5_port, B(4) => 
                           out_imux_11_4_port, B(3) => out_imux_11_3_port, B(2)
                           => out_imux_11_2_port, B(1) => out_imux_11_1_port, 
                           B(0) => out_imux_11_0_port, Ci => X_Logic0_port, 
                           S(63) => predigest_product_11_63_port, S(62) => 
                           predigest_product_11_62_port, S(61) => 
                           predigest_product_11_61_port, S(60) => 
                           predigest_product_11_60_port, S(59) => 
                           predigest_product_11_59_port, S(58) => 
                           predigest_product_11_58_port, S(57) => 
                           predigest_product_11_57_port, S(56) => 
                           predigest_product_11_56_port, S(55) => 
                           predigest_product_11_55_port, S(54) => 
                           predigest_product_11_54_port, S(53) => 
                           predigest_product_11_53_port, S(52) => 
                           predigest_product_11_52_port, S(51) => 
                           predigest_product_11_51_port, S(50) => 
                           predigest_product_11_50_port, S(49) => 
                           predigest_product_11_49_port, S(48) => 
                           predigest_product_11_48_port, S(47) => 
                           predigest_product_11_47_port, S(46) => 
                           predigest_product_11_46_port, S(45) => 
                           predigest_product_11_45_port, S(44) => 
                           predigest_product_11_44_port, S(43) => 
                           predigest_product_11_43_port, S(42) => 
                           predigest_product_11_42_port, S(41) => 
                           predigest_product_11_41_port, S(40) => 
                           predigest_product_11_40_port, S(39) => 
                           predigest_product_11_39_port, S(38) => 
                           predigest_product_11_38_port, S(37) => 
                           predigest_product_11_37_port, S(36) => 
                           predigest_product_11_36_port, S(35) => 
                           predigest_product_11_35_port, S(34) => 
                           predigest_product_11_34_port, S(33) => 
                           predigest_product_11_33_port, S(32) => 
                           predigest_product_11_32_port, S(31) => 
                           predigest_product_11_31_port, S(30) => 
                           predigest_product_11_30_port, S(29) => 
                           predigest_product_11_29_port, S(28) => 
                           predigest_product_11_28_port, S(27) => 
                           predigest_product_11_27_port, S(26) => 
                           predigest_product_11_26_port, S(25) => 
                           predigest_product_11_25_port, S(24) => 
                           predigest_product_11_24_port, S(23) => 
                           predigest_product_11_23_port, S(22) => 
                           predigest_product_11_22_port, S(21) => 
                           predigest_product_11_21_port, S(20) => 
                           predigest_product_11_20_port, S(19) => 
                           predigest_product_11_19_port, S(18) => 
                           predigest_product_11_18_port, S(17) => 
                           predigest_product_11_17_port, S(16) => 
                           predigest_product_11_16_port, S(15) => 
                           predigest_product_11_15_port, S(14) => 
                           predigest_product_11_14_port, S(13) => 
                           predigest_product_11_13_port, S(12) => 
                           predigest_product_11_12_port, S(11) => 
                           predigest_product_11_11_port, S(10) => 
                           predigest_product_11_10_port, S(9) => 
                           predigest_product_11_9_port, S(8) => 
                           predigest_product_11_8_port, S(7) => 
                           predigest_product_11_7_port, S(6) => 
                           predigest_product_11_6_port, S(5) => 
                           predigest_product_11_5_port, S(4) => 
                           predigest_product_11_4_port, S(3) => 
                           predigest_product_11_3_port, S(2) => 
                           predigest_product_11_2_port, S(1) => 
                           predigest_product_11_1_port, S(0) => 
                           predigest_product_11_0_port, Co => n_1102);
   ENC_i_12 : BOOTH_ENCODER_3BIT_8 port map( B(2) => B(25), B(1) => B(24), B(0)
                           => B(23), ENCODED(2) => 
                           muxs_encoded_signals_12_2_port, ENCODED(1) => 
                           muxs_encoded_signals_12_1_port, ENCODED(0) => 
                           muxs_encoded_signals_12_0_port);
   MUX_i_12 : MUX51_GENERIC_NBIT64_4 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(31), IN1(55) => A(31), IN1(54) => 
                           A(30), IN1(53) => A(29), IN1(52) => A(28), IN1(51) 
                           => A(27), IN1(50) => A(26), IN1(49) => A(25), 
                           IN1(48) => A(24), IN1(47) => A(23), IN1(46) => A(22)
                           , IN1(45) => A(21), IN1(44) => A(20), IN1(43) => 
                           A(19), IN1(42) => A(18), IN1(41) => A(17), IN1(40) 
                           => A(16), IN1(39) => A(15), IN1(38) => A(14), 
                           IN1(37) => A(13), IN1(36) => A(12), IN1(35) => A(11)
                           , IN1(34) => A(10), IN1(33) => A(9), IN1(32) => A(8)
                           , IN1(31) => A(7), IN1(30) => A(6), IN1(29) => A(5),
                           IN1(28) => A(4), IN1(27) => A(3), IN1(26) => A(2), 
                           IN1(25) => A(1), IN1(24) => A(0), IN1(23) => 
                           X_Logic0_port, IN1(22) => X_Logic0_port, IN1(21) => 
                           X_Logic0_port, IN1(20) => X_Logic0_port, IN1(19) => 
                           X_Logic0_port, IN1(18) => X_Logic0_port, IN1(17) => 
                           X_Logic0_port, IN1(16) => X_Logic0_port, IN1(15) => 
                           X_Logic0_port, IN1(14) => X_Logic0_port, IN1(13) => 
                           X_Logic0_port, IN1(12) => X_Logic0_port, IN1(11) => 
                           X_Logic0_port, IN1(10) => X_Logic0_port, IN1(9) => 
                           X_Logic0_port, IN1(8) => X_Logic0_port, IN1(7) => 
                           X_Logic0_port, IN1(6) => X_Logic0_port, IN1(5) => 
                           X_Logic0_port, IN1(4) => X_Logic0_port, IN1(3) => 
                           X_Logic0_port, IN1(2) => X_Logic0_port, IN1(1) => 
                           X_Logic0_port, IN1(0) => X_Logic0_port, IN2(63) => 
                           negative_a_39_port, IN2(62) => negative_a_38_port, 
                           IN2(61) => negative_a_37_port, IN2(60) => 
                           negative_a_36_port, IN2(59) => negative_a_35_port, 
                           IN2(58) => negative_a_34_port, IN2(57) => n38, 
                           IN2(56) => n35, IN2(55) => negative_a_31_port, 
                           IN2(54) => negative_a_30_port, IN2(53) => 
                           negative_a_29_port, IN2(52) => negative_a_28_port, 
                           IN2(51) => negative_a_27_port, IN2(50) => 
                           negative_a_26_port, IN2(49) => negative_a_25_port, 
                           IN2(48) => negative_a_24_port, IN2(47) => 
                           negative_a_23_port, IN2(46) => negative_a_22_port, 
                           IN2(45) => negative_a_21_port, IN2(44) => 
                           negative_a_20_port, IN2(43) => negative_a_19_port, 
                           IN2(42) => negative_a_18_port, IN2(41) => 
                           negative_a_17_port, IN2(40) => negative_a_16_port, 
                           IN2(39) => negative_a_15_port, IN2(38) => 
                           negative_a_14_port, IN2(37) => negative_a_13_port, 
                           IN2(36) => negative_a_12_port, IN2(35) => 
                           negative_a_11_port, IN2(34) => negative_a_10_port, 
                           IN2(33) => negative_a_9_port, IN2(32) => 
                           negative_a_8_port, IN2(31) => negative_a_7_port, 
                           IN2(30) => negative_a_6_port, IN2(29) => 
                           negative_a_5_port, IN2(28) => negative_a_4_port, 
                           IN2(27) => negative_a_3_port, IN2(26) => 
                           negative_a_2_port, IN2(25) => negative_a_1_port, 
                           IN2(24) => negative_a_0_port, IN2(23) => 
                           X_Logic0_port, IN2(22) => X_Logic0_port, IN2(21) => 
                           X_Logic0_port, IN2(20) => X_Logic0_port, IN2(19) => 
                           X_Logic0_port, IN2(18) => X_Logic0_port, IN2(17) => 
                           X_Logic0_port, IN2(16) => X_Logic0_port, IN2(15) => 
                           X_Logic0_port, IN2(14) => X_Logic0_port, IN2(13) => 
                           X_Logic0_port, IN2(12) => X_Logic0_port, IN2(11) => 
                           X_Logic0_port, IN2(10) => X_Logic0_port, IN2(9) => 
                           X_Logic0_port, IN2(8) => X_Logic0_port, IN2(7) => 
                           X_Logic0_port, IN2(6) => X_Logic0_port, IN2(5) => 
                           X_Logic0_port, IN2(4) => X_Logic0_port, IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(63) => 
                           A(31), IN3(62) => A(31), IN3(61) => A(31), IN3(60) 
                           => A(31), IN3(59) => A(31), IN3(58) => A(31), 
                           IN3(57) => A(31), IN3(56) => A(31), IN3(55) => A(30)
                           , IN3(54) => A(29), IN3(53) => A(28), IN3(52) => 
                           A(27), IN3(51) => A(26), IN3(50) => A(25), IN3(49) 
                           => A(24), IN3(48) => A(23), IN3(47) => A(22), 
                           IN3(46) => A(21), IN3(45) => A(20), IN3(44) => A(19)
                           , IN3(43) => A(18), IN3(42) => A(17), IN3(41) => 
                           A(16), IN3(40) => A(15), IN3(39) => A(14), IN3(38) 
                           => A(13), IN3(37) => A(12), IN3(36) => A(11), 
                           IN3(35) => A(10), IN3(34) => A(9), IN3(33) => A(8), 
                           IN3(32) => A(7), IN3(31) => A(6), IN3(30) => A(5), 
                           IN3(29) => A(4), IN3(28) => A(3), IN3(27) => A(2), 
                           IN3(26) => A(1), IN3(25) => A(0), IN3(24) => 
                           X_Logic0_port, IN3(23) => X_Logic0_port, IN3(22) => 
                           X_Logic0_port, IN3(21) => X_Logic0_port, IN3(20) => 
                           X_Logic0_port, IN3(19) => X_Logic0_port, IN3(18) => 
                           X_Logic0_port, IN3(17) => X_Logic0_port, IN3(16) => 
                           X_Logic0_port, IN3(15) => X_Logic0_port, IN3(14) => 
                           X_Logic0_port, IN3(13) => X_Logic0_port, IN3(12) => 
                           X_Logic0_port, IN3(11) => X_Logic0_port, IN3(10) => 
                           X_Logic0_port, IN3(9) => X_Logic0_port, IN3(8) => 
                           X_Logic0_port, IN3(7) => X_Logic0_port, IN3(6) => 
                           X_Logic0_port, IN3(5) => X_Logic0_port, IN3(4) => 
                           X_Logic0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(63) => negative_a_38_port, 
                           IN4(62) => negative_a_37_port, IN4(61) => 
                           negative_a_36_port, IN4(60) => negative_a_35_port, 
                           IN4(59) => negative_a_34_port, IN4(58) => n38, 
                           IN4(57) => n35, IN4(56) => negative_a_31_port, 
                           IN4(55) => negative_a_30_port, IN4(54) => 
                           negative_a_29_port, IN4(53) => negative_a_28_port, 
                           IN4(52) => negative_a_27_port, IN4(51) => 
                           negative_a_26_port, IN4(50) => negative_a_25_port, 
                           IN4(49) => negative_a_24_port, IN4(48) => 
                           negative_a_23_port, IN4(47) => negative_a_22_port, 
                           IN4(46) => negative_a_21_port, IN4(45) => 
                           negative_a_20_port, IN4(44) => negative_a_19_port, 
                           IN4(43) => negative_a_18_port, IN4(42) => 
                           negative_a_17_port, IN4(41) => negative_a_16_port, 
                           IN4(40) => negative_a_15_port, IN4(39) => 
                           negative_a_14_port, IN4(38) => negative_a_13_port, 
                           IN4(37) => negative_a_12_port, IN4(36) => 
                           negative_a_11_port, IN4(35) => negative_a_10_port, 
                           IN4(34) => negative_a_9_port, IN4(33) => 
                           negative_a_8_port, IN4(32) => negative_a_7_port, 
                           IN4(31) => negative_a_6_port, IN4(30) => 
                           negative_a_5_port, IN4(29) => negative_a_4_port, 
                           IN4(28) => negative_a_3_port, IN4(27) => 
                           negative_a_2_port, IN4(26) => negative_a_1_port, 
                           IN4(25) => negative_a_0_port, IN4(24) => 
                           X_Logic0_port, IN4(23) => X_Logic0_port, IN4(22) => 
                           X_Logic0_port, IN4(21) => X_Logic0_port, IN4(20) => 
                           X_Logic0_port, IN4(19) => X_Logic0_port, IN4(18) => 
                           X_Logic0_port, IN4(17) => X_Logic0_port, IN4(16) => 
                           X_Logic0_port, IN4(15) => X_Logic0_port, IN4(14) => 
                           X_Logic0_port, IN4(13) => X_Logic0_port, IN4(12) => 
                           X_Logic0_port, IN4(11) => X_Logic0_port, IN4(10) => 
                           X_Logic0_port, IN4(9) => X_Logic0_port, IN4(8) => 
                           X_Logic0_port, IN4(7) => X_Logic0_port, IN4(6) => 
                           X_Logic0_port, IN4(5) => X_Logic0_port, IN4(4) => 
                           X_Logic0_port, IN4(3) => X_Logic0_port, IN4(2) => 
                           X_Logic0_port, IN4(1) => X_Logic0_port, IN4(0) => 
                           X_Logic0_port, S(2) => 
                           muxs_encoded_signals_12_2_port, S(1) => 
                           muxs_encoded_signals_12_1_port, S(0) => 
                           muxs_encoded_signals_12_0_port, O(63) => 
                           out_imux_12_63_port, O(62) => out_imux_12_62_port, 
                           O(61) => out_imux_12_61_port, O(60) => 
                           out_imux_12_60_port, O(59) => out_imux_12_59_port, 
                           O(58) => out_imux_12_58_port, O(57) => 
                           out_imux_12_57_port, O(56) => out_imux_12_56_port, 
                           O(55) => out_imux_12_55_port, O(54) => 
                           out_imux_12_54_port, O(53) => out_imux_12_53_port, 
                           O(52) => out_imux_12_52_port, O(51) => 
                           out_imux_12_51_port, O(50) => out_imux_12_50_port, 
                           O(49) => out_imux_12_49_port, O(48) => 
                           out_imux_12_48_port, O(47) => out_imux_12_47_port, 
                           O(46) => out_imux_12_46_port, O(45) => 
                           out_imux_12_45_port, O(44) => out_imux_12_44_port, 
                           O(43) => out_imux_12_43_port, O(42) => 
                           out_imux_12_42_port, O(41) => out_imux_12_41_port, 
                           O(40) => out_imux_12_40_port, O(39) => 
                           out_imux_12_39_port, O(38) => out_imux_12_38_port, 
                           O(37) => out_imux_12_37_port, O(36) => 
                           out_imux_12_36_port, O(35) => out_imux_12_35_port, 
                           O(34) => out_imux_12_34_port, O(33) => 
                           out_imux_12_33_port, O(32) => out_imux_12_32_port, 
                           O(31) => out_imux_12_31_port, O(30) => 
                           out_imux_12_30_port, O(29) => out_imux_12_29_port, 
                           O(28) => out_imux_12_28_port, O(27) => 
                           out_imux_12_27_port, O(26) => out_imux_12_26_port, 
                           O(25) => out_imux_12_25_port, O(24) => 
                           out_imux_12_24_port, O(23) => out_imux_12_23_port, 
                           O(22) => out_imux_12_22_port, O(21) => 
                           out_imux_12_21_port, O(20) => out_imux_12_20_port, 
                           O(19) => out_imux_12_19_port, O(18) => 
                           out_imux_12_18_port, O(17) => out_imux_12_17_port, 
                           O(16) => out_imux_12_16_port, O(15) => 
                           out_imux_12_15_port, O(14) => out_imux_12_14_port, 
                           O(13) => out_imux_12_13_port, O(12) => 
                           out_imux_12_12_port, O(11) => out_imux_12_11_port, 
                           O(10) => out_imux_12_10_port, O(9) => 
                           out_imux_12_9_port, O(8) => out_imux_12_8_port, O(7)
                           => out_imux_12_7_port, O(6) => out_imux_12_6_port, 
                           O(5) => out_imux_12_5_port, O(4) => 
                           out_imux_12_4_port, O(3) => out_imux_12_3_port, O(2)
                           => out_imux_12_2_port, O(1) => out_imux_12_1_port, 
                           O(0) => out_imux_12_0_port);
   ADD64_i_12 : RCA_GENERIC_NBIT64_4 port map( A(63) => 
                           predigest_product_11_63_port, A(62) => 
                           predigest_product_11_62_port, A(61) => 
                           predigest_product_11_61_port, A(60) => 
                           predigest_product_11_60_port, A(59) => 
                           predigest_product_11_59_port, A(58) => 
                           predigest_product_11_58_port, A(57) => 
                           predigest_product_11_57_port, A(56) => 
                           predigest_product_11_56_port, A(55) => 
                           predigest_product_11_55_port, A(54) => 
                           predigest_product_11_54_port, A(53) => 
                           predigest_product_11_53_port, A(52) => 
                           predigest_product_11_52_port, A(51) => 
                           predigest_product_11_51_port, A(50) => 
                           predigest_product_11_50_port, A(49) => 
                           predigest_product_11_49_port, A(48) => 
                           predigest_product_11_48_port, A(47) => 
                           predigest_product_11_47_port, A(46) => 
                           predigest_product_11_46_port, A(45) => 
                           predigest_product_11_45_port, A(44) => 
                           predigest_product_11_44_port, A(43) => 
                           predigest_product_11_43_port, A(42) => 
                           predigest_product_11_42_port, A(41) => 
                           predigest_product_11_41_port, A(40) => 
                           predigest_product_11_40_port, A(39) => 
                           predigest_product_11_39_port, A(38) => 
                           predigest_product_11_38_port, A(37) => 
                           predigest_product_11_37_port, A(36) => 
                           predigest_product_11_36_port, A(35) => 
                           predigest_product_11_35_port, A(34) => 
                           predigest_product_11_34_port, A(33) => 
                           predigest_product_11_33_port, A(32) => 
                           predigest_product_11_32_port, A(31) => 
                           predigest_product_11_31_port, A(30) => 
                           predigest_product_11_30_port, A(29) => 
                           predigest_product_11_29_port, A(28) => 
                           predigest_product_11_28_port, A(27) => 
                           predigest_product_11_27_port, A(26) => 
                           predigest_product_11_26_port, A(25) => 
                           predigest_product_11_25_port, A(24) => 
                           predigest_product_11_24_port, A(23) => 
                           predigest_product_11_23_port, A(22) => 
                           predigest_product_11_22_port, A(21) => 
                           predigest_product_11_21_port, A(20) => 
                           predigest_product_11_20_port, A(19) => 
                           predigest_product_11_19_port, A(18) => 
                           predigest_product_11_18_port, A(17) => 
                           predigest_product_11_17_port, A(16) => 
                           predigest_product_11_16_port, A(15) => 
                           predigest_product_11_15_port, A(14) => 
                           predigest_product_11_14_port, A(13) => 
                           predigest_product_11_13_port, A(12) => 
                           predigest_product_11_12_port, A(11) => 
                           predigest_product_11_11_port, A(10) => 
                           predigest_product_11_10_port, A(9) => 
                           predigest_product_11_9_port, A(8) => 
                           predigest_product_11_8_port, A(7) => 
                           predigest_product_11_7_port, A(6) => 
                           predigest_product_11_6_port, A(5) => 
                           predigest_product_11_5_port, A(4) => 
                           predigest_product_11_4_port, A(3) => 
                           predigest_product_11_3_port, A(2) => 
                           predigest_product_11_2_port, A(1) => 
                           predigest_product_11_1_port, A(0) => 
                           predigest_product_11_0_port, B(63) => 
                           out_imux_12_63_port, B(62) => out_imux_12_62_port, 
                           B(61) => out_imux_12_61_port, B(60) => 
                           out_imux_12_60_port, B(59) => out_imux_12_59_port, 
                           B(58) => out_imux_12_58_port, B(57) => 
                           out_imux_12_57_port, B(56) => out_imux_12_56_port, 
                           B(55) => out_imux_12_55_port, B(54) => 
                           out_imux_12_54_port, B(53) => out_imux_12_53_port, 
                           B(52) => out_imux_12_52_port, B(51) => 
                           out_imux_12_51_port, B(50) => out_imux_12_50_port, 
                           B(49) => out_imux_12_49_port, B(48) => 
                           out_imux_12_48_port, B(47) => out_imux_12_47_port, 
                           B(46) => out_imux_12_46_port, B(45) => 
                           out_imux_12_45_port, B(44) => out_imux_12_44_port, 
                           B(43) => out_imux_12_43_port, B(42) => 
                           out_imux_12_42_port, B(41) => out_imux_12_41_port, 
                           B(40) => out_imux_12_40_port, B(39) => 
                           out_imux_12_39_port, B(38) => out_imux_12_38_port, 
                           B(37) => out_imux_12_37_port, B(36) => 
                           out_imux_12_36_port, B(35) => out_imux_12_35_port, 
                           B(34) => out_imux_12_34_port, B(33) => 
                           out_imux_12_33_port, B(32) => out_imux_12_32_port, 
                           B(31) => out_imux_12_31_port, B(30) => 
                           out_imux_12_30_port, B(29) => out_imux_12_29_port, 
                           B(28) => out_imux_12_28_port, B(27) => 
                           out_imux_12_27_port, B(26) => out_imux_12_26_port, 
                           B(25) => out_imux_12_25_port, B(24) => 
                           out_imux_12_24_port, B(23) => out_imux_12_23_port, 
                           B(22) => out_imux_12_22_port, B(21) => 
                           out_imux_12_21_port, B(20) => out_imux_12_20_port, 
                           B(19) => out_imux_12_19_port, B(18) => 
                           out_imux_12_18_port, B(17) => out_imux_12_17_port, 
                           B(16) => out_imux_12_16_port, B(15) => 
                           out_imux_12_15_port, B(14) => out_imux_12_14_port, 
                           B(13) => out_imux_12_13_port, B(12) => 
                           out_imux_12_12_port, B(11) => out_imux_12_11_port, 
                           B(10) => out_imux_12_10_port, B(9) => 
                           out_imux_12_9_port, B(8) => out_imux_12_8_port, B(7)
                           => out_imux_12_7_port, B(6) => out_imux_12_6_port, 
                           B(5) => out_imux_12_5_port, B(4) => 
                           out_imux_12_4_port, B(3) => out_imux_12_3_port, B(2)
                           => out_imux_12_2_port, B(1) => out_imux_12_1_port, 
                           B(0) => out_imux_12_0_port, Ci => X_Logic0_port, 
                           S(63) => predigest_product_12_63_port, S(62) => 
                           predigest_product_12_62_port, S(61) => 
                           predigest_product_12_61_port, S(60) => 
                           predigest_product_12_60_port, S(59) => 
                           predigest_product_12_59_port, S(58) => 
                           predigest_product_12_58_port, S(57) => 
                           predigest_product_12_57_port, S(56) => 
                           predigest_product_12_56_port, S(55) => 
                           predigest_product_12_55_port, S(54) => 
                           predigest_product_12_54_port, S(53) => 
                           predigest_product_12_53_port, S(52) => 
                           predigest_product_12_52_port, S(51) => 
                           predigest_product_12_51_port, S(50) => 
                           predigest_product_12_50_port, S(49) => 
                           predigest_product_12_49_port, S(48) => 
                           predigest_product_12_48_port, S(47) => 
                           predigest_product_12_47_port, S(46) => 
                           predigest_product_12_46_port, S(45) => 
                           predigest_product_12_45_port, S(44) => 
                           predigest_product_12_44_port, S(43) => 
                           predigest_product_12_43_port, S(42) => 
                           predigest_product_12_42_port, S(41) => 
                           predigest_product_12_41_port, S(40) => 
                           predigest_product_12_40_port, S(39) => 
                           predigest_product_12_39_port, S(38) => 
                           predigest_product_12_38_port, S(37) => 
                           predigest_product_12_37_port, S(36) => 
                           predigest_product_12_36_port, S(35) => 
                           predigest_product_12_35_port, S(34) => 
                           predigest_product_12_34_port, S(33) => 
                           predigest_product_12_33_port, S(32) => 
                           predigest_product_12_32_port, S(31) => 
                           predigest_product_12_31_port, S(30) => 
                           predigest_product_12_30_port, S(29) => 
                           predigest_product_12_29_port, S(28) => 
                           predigest_product_12_28_port, S(27) => 
                           predigest_product_12_27_port, S(26) => 
                           predigest_product_12_26_port, S(25) => 
                           predigest_product_12_25_port, S(24) => 
                           predigest_product_12_24_port, S(23) => 
                           predigest_product_12_23_port, S(22) => 
                           predigest_product_12_22_port, S(21) => 
                           predigest_product_12_21_port, S(20) => 
                           predigest_product_12_20_port, S(19) => 
                           predigest_product_12_19_port, S(18) => 
                           predigest_product_12_18_port, S(17) => 
                           predigest_product_12_17_port, S(16) => 
                           predigest_product_12_16_port, S(15) => 
                           predigest_product_12_15_port, S(14) => 
                           predigest_product_12_14_port, S(13) => 
                           predigest_product_12_13_port, S(12) => 
                           predigest_product_12_12_port, S(11) => 
                           predigest_product_12_11_port, S(10) => 
                           predigest_product_12_10_port, S(9) => 
                           predigest_product_12_9_port, S(8) => 
                           predigest_product_12_8_port, S(7) => 
                           predigest_product_12_7_port, S(6) => 
                           predigest_product_12_6_port, S(5) => 
                           predigest_product_12_5_port, S(4) => 
                           predigest_product_12_4_port, S(3) => 
                           predigest_product_12_3_port, S(2) => 
                           predigest_product_12_2_port, S(1) => 
                           predigest_product_12_1_port, S(0) => 
                           predigest_product_12_0_port, Co => n_1103);
   ENC_i_13 : BOOTH_ENCODER_3BIT_7 port map( B(2) => B(27), B(1) => B(26), B(0)
                           => B(25), ENCODED(2) => 
                           muxs_encoded_signals_13_2_port, ENCODED(1) => 
                           muxs_encoded_signals_13_1_port, ENCODED(0) => 
                           muxs_encoded_signals_13_0_port);
   MUX_i_13 : MUX51_GENERIC_NBIT64_3 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(31), IN1(57) => A(31)
                           , IN1(56) => A(30), IN1(55) => A(29), IN1(54) => 
                           A(28), IN1(53) => A(27), IN1(52) => A(26), IN1(51) 
                           => A(25), IN1(50) => A(24), IN1(49) => A(23), 
                           IN1(48) => A(22), IN1(47) => A(21), IN1(46) => A(20)
                           , IN1(45) => A(19), IN1(44) => A(18), IN1(43) => 
                           A(17), IN1(42) => A(16), IN1(41) => A(15), IN1(40) 
                           => A(14), IN1(39) => A(13), IN1(38) => A(12), 
                           IN1(37) => A(11), IN1(36) => A(10), IN1(35) => A(9),
                           IN1(34) => A(8), IN1(33) => A(7), IN1(32) => A(6), 
                           IN1(31) => A(5), IN1(30) => A(4), IN1(29) => A(3), 
                           IN1(28) => A(2), IN1(27) => A(1), IN1(26) => A(0), 
                           IN1(25) => X_Logic0_port, IN1(24) => X_Logic0_port, 
                           IN1(23) => X_Logic0_port, IN1(22) => X_Logic0_port, 
                           IN1(21) => X_Logic0_port, IN1(20) => X_Logic0_port, 
                           IN1(19) => X_Logic0_port, IN1(18) => X_Logic0_port, 
                           IN1(17) => X_Logic0_port, IN1(16) => X_Logic0_port, 
                           IN1(15) => X_Logic0_port, IN1(14) => X_Logic0_port, 
                           IN1(13) => X_Logic0_port, IN1(12) => X_Logic0_port, 
                           IN1(11) => X_Logic0_port, IN1(10) => X_Logic0_port, 
                           IN1(9) => X_Logic0_port, IN1(8) => X_Logic0_port, 
                           IN1(7) => X_Logic0_port, IN1(6) => X_Logic0_port, 
                           IN1(5) => X_Logic0_port, IN1(4) => X_Logic0_port, 
                           IN1(3) => X_Logic0_port, IN1(2) => X_Logic0_port, 
                           IN1(1) => X_Logic0_port, IN1(0) => X_Logic0_port, 
                           IN2(63) => negative_a_37_port, IN2(62) => 
                           negative_a_36_port, IN2(61) => negative_a_35_port, 
                           IN2(60) => negative_a_34_port, IN2(59) => n38, 
                           IN2(58) => n35, IN2(57) => negative_a_31_port, 
                           IN2(56) => negative_a_30_port, IN2(55) => 
                           negative_a_29_port, IN2(54) => negative_a_28_port, 
                           IN2(53) => negative_a_27_port, IN2(52) => 
                           negative_a_26_port, IN2(51) => negative_a_25_port, 
                           IN2(50) => negative_a_24_port, IN2(49) => 
                           negative_a_23_port, IN2(48) => negative_a_22_port, 
                           IN2(47) => negative_a_21_port, IN2(46) => 
                           negative_a_20_port, IN2(45) => negative_a_19_port, 
                           IN2(44) => negative_a_18_port, IN2(43) => 
                           negative_a_17_port, IN2(42) => negative_a_16_port, 
                           IN2(41) => negative_a_15_port, IN2(40) => 
                           negative_a_14_port, IN2(39) => negative_a_13_port, 
                           IN2(38) => negative_a_12_port, IN2(37) => 
                           negative_a_11_port, IN2(36) => negative_a_10_port, 
                           IN2(35) => negative_a_9_port, IN2(34) => 
                           negative_a_8_port, IN2(33) => negative_a_7_port, 
                           IN2(32) => negative_a_6_port, IN2(31) => 
                           negative_a_5_port, IN2(30) => negative_a_4_port, 
                           IN2(29) => negative_a_3_port, IN2(28) => 
                           negative_a_2_port, IN2(27) => negative_a_1_port, 
                           IN2(26) => negative_a_0_port, IN2(25) => 
                           X_Logic0_port, IN2(24) => X_Logic0_port, IN2(23) => 
                           X_Logic0_port, IN2(22) => X_Logic0_port, IN2(21) => 
                           X_Logic0_port, IN2(20) => X_Logic0_port, IN2(19) => 
                           X_Logic0_port, IN2(18) => X_Logic0_port, IN2(17) => 
                           X_Logic0_port, IN2(16) => X_Logic0_port, IN2(15) => 
                           X_Logic0_port, IN2(14) => X_Logic0_port, IN2(13) => 
                           X_Logic0_port, IN2(12) => X_Logic0_port, IN2(11) => 
                           X_Logic0_port, IN2(10) => X_Logic0_port, IN2(9) => 
                           X_Logic0_port, IN2(8) => X_Logic0_port, IN2(7) => 
                           X_Logic0_port, IN2(6) => X_Logic0_port, IN2(5) => 
                           X_Logic0_port, IN2(4) => X_Logic0_port, IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(63) => 
                           A(31), IN3(62) => A(31), IN3(61) => A(31), IN3(60) 
                           => A(31), IN3(59) => A(31), IN3(58) => A(31), 
                           IN3(57) => A(30), IN3(56) => A(29), IN3(55) => A(28)
                           , IN3(54) => A(27), IN3(53) => A(26), IN3(52) => 
                           A(25), IN3(51) => A(24), IN3(50) => A(23), IN3(49) 
                           => A(22), IN3(48) => A(21), IN3(47) => A(20), 
                           IN3(46) => A(19), IN3(45) => A(18), IN3(44) => A(17)
                           , IN3(43) => A(16), IN3(42) => A(15), IN3(41) => 
                           A(14), IN3(40) => A(13), IN3(39) => A(12), IN3(38) 
                           => A(11), IN3(37) => A(10), IN3(36) => A(9), IN3(35)
                           => A(8), IN3(34) => A(7), IN3(33) => A(6), IN3(32) 
                           => A(5), IN3(31) => A(4), IN3(30) => A(3), IN3(29) 
                           => A(2), IN3(28) => A(1), IN3(27) => A(0), IN3(26) 
                           => X_Logic0_port, IN3(25) => X_Logic0_port, IN3(24) 
                           => X_Logic0_port, IN3(23) => X_Logic0_port, IN3(22) 
                           => X_Logic0_port, IN3(21) => X_Logic0_port, IN3(20) 
                           => X_Logic0_port, IN3(19) => X_Logic0_port, IN3(18) 
                           => X_Logic0_port, IN3(17) => X_Logic0_port, IN3(16) 
                           => X_Logic0_port, IN3(15) => X_Logic0_port, IN3(14) 
                           => X_Logic0_port, IN3(13) => X_Logic0_port, IN3(12) 
                           => X_Logic0_port, IN3(11) => X_Logic0_port, IN3(10) 
                           => X_Logic0_port, IN3(9) => X_Logic0_port, IN3(8) =>
                           X_Logic0_port, IN3(7) => X_Logic0_port, IN3(6) => 
                           X_Logic0_port, IN3(5) => X_Logic0_port, IN3(4) => 
                           X_Logic0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(63) => negative_a_36_port, 
                           IN4(62) => negative_a_35_port, IN4(61) => 
                           negative_a_34_port, IN4(60) => n38, IN4(59) => n35, 
                           IN4(58) => negative_a_31_port, IN4(57) => 
                           negative_a_30_port, IN4(56) => negative_a_29_port, 
                           IN4(55) => negative_a_28_port, IN4(54) => 
                           negative_a_27_port, IN4(53) => negative_a_26_port, 
                           IN4(52) => negative_a_25_port, IN4(51) => 
                           negative_a_24_port, IN4(50) => negative_a_23_port, 
                           IN4(49) => negative_a_22_port, IN4(48) => 
                           negative_a_21_port, IN4(47) => negative_a_20_port, 
                           IN4(46) => negative_a_19_port, IN4(45) => 
                           negative_a_18_port, IN4(44) => negative_a_17_port, 
                           IN4(43) => negative_a_16_port, IN4(42) => 
                           negative_a_15_port, IN4(41) => negative_a_14_port, 
                           IN4(40) => negative_a_13_port, IN4(39) => 
                           negative_a_12_port, IN4(38) => negative_a_11_port, 
                           IN4(37) => negative_a_10_port, IN4(36) => 
                           negative_a_9_port, IN4(35) => negative_a_8_port, 
                           IN4(34) => negative_a_7_port, IN4(33) => 
                           negative_a_6_port, IN4(32) => negative_a_5_port, 
                           IN4(31) => negative_a_4_port, IN4(30) => 
                           negative_a_3_port, IN4(29) => negative_a_2_port, 
                           IN4(28) => negative_a_1_port, IN4(27) => 
                           negative_a_0_port, IN4(26) => X_Logic0_port, IN4(25)
                           => X_Logic0_port, IN4(24) => X_Logic0_port, IN4(23) 
                           => X_Logic0_port, IN4(22) => X_Logic0_port, IN4(21) 
                           => X_Logic0_port, IN4(20) => X_Logic0_port, IN4(19) 
                           => X_Logic0_port, IN4(18) => X_Logic0_port, IN4(17) 
                           => X_Logic0_port, IN4(16) => X_Logic0_port, IN4(15) 
                           => X_Logic0_port, IN4(14) => X_Logic0_port, IN4(13) 
                           => X_Logic0_port, IN4(12) => X_Logic0_port, IN4(11) 
                           => X_Logic0_port, IN4(10) => X_Logic0_port, IN4(9) 
                           => X_Logic0_port, IN4(8) => X_Logic0_port, IN4(7) =>
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_13_2_port, S(1) => 
                           muxs_encoded_signals_13_1_port, S(0) => 
                           muxs_encoded_signals_13_0_port, O(63) => 
                           out_imux_13_63_port, O(62) => out_imux_13_62_port, 
                           O(61) => out_imux_13_61_port, O(60) => 
                           out_imux_13_60_port, O(59) => out_imux_13_59_port, 
                           O(58) => out_imux_13_58_port, O(57) => 
                           out_imux_13_57_port, O(56) => out_imux_13_56_port, 
                           O(55) => out_imux_13_55_port, O(54) => 
                           out_imux_13_54_port, O(53) => out_imux_13_53_port, 
                           O(52) => out_imux_13_52_port, O(51) => 
                           out_imux_13_51_port, O(50) => out_imux_13_50_port, 
                           O(49) => out_imux_13_49_port, O(48) => 
                           out_imux_13_48_port, O(47) => out_imux_13_47_port, 
                           O(46) => out_imux_13_46_port, O(45) => 
                           out_imux_13_45_port, O(44) => out_imux_13_44_port, 
                           O(43) => out_imux_13_43_port, O(42) => 
                           out_imux_13_42_port, O(41) => out_imux_13_41_port, 
                           O(40) => out_imux_13_40_port, O(39) => 
                           out_imux_13_39_port, O(38) => out_imux_13_38_port, 
                           O(37) => out_imux_13_37_port, O(36) => 
                           out_imux_13_36_port, O(35) => out_imux_13_35_port, 
                           O(34) => out_imux_13_34_port, O(33) => 
                           out_imux_13_33_port, O(32) => out_imux_13_32_port, 
                           O(31) => out_imux_13_31_port, O(30) => 
                           out_imux_13_30_port, O(29) => out_imux_13_29_port, 
                           O(28) => out_imux_13_28_port, O(27) => 
                           out_imux_13_27_port, O(26) => out_imux_13_26_port, 
                           O(25) => out_imux_13_25_port, O(24) => 
                           out_imux_13_24_port, O(23) => out_imux_13_23_port, 
                           O(22) => out_imux_13_22_port, O(21) => 
                           out_imux_13_21_port, O(20) => out_imux_13_20_port, 
                           O(19) => out_imux_13_19_port, O(18) => 
                           out_imux_13_18_port, O(17) => out_imux_13_17_port, 
                           O(16) => out_imux_13_16_port, O(15) => 
                           out_imux_13_15_port, O(14) => out_imux_13_14_port, 
                           O(13) => out_imux_13_13_port, O(12) => 
                           out_imux_13_12_port, O(11) => out_imux_13_11_port, 
                           O(10) => out_imux_13_10_port, O(9) => 
                           out_imux_13_9_port, O(8) => out_imux_13_8_port, O(7)
                           => out_imux_13_7_port, O(6) => out_imux_13_6_port, 
                           O(5) => out_imux_13_5_port, O(4) => 
                           out_imux_13_4_port, O(3) => out_imux_13_3_port, O(2)
                           => out_imux_13_2_port, O(1) => out_imux_13_1_port, 
                           O(0) => out_imux_13_0_port);
   ADD64_i_13 : RCA_GENERIC_NBIT64_3 port map( A(63) => 
                           predigest_product_12_63_port, A(62) => 
                           predigest_product_12_62_port, A(61) => 
                           predigest_product_12_61_port, A(60) => 
                           predigest_product_12_60_port, A(59) => 
                           predigest_product_12_59_port, A(58) => 
                           predigest_product_12_58_port, A(57) => 
                           predigest_product_12_57_port, A(56) => 
                           predigest_product_12_56_port, A(55) => 
                           predigest_product_12_55_port, A(54) => 
                           predigest_product_12_54_port, A(53) => 
                           predigest_product_12_53_port, A(52) => 
                           predigest_product_12_52_port, A(51) => 
                           predigest_product_12_51_port, A(50) => 
                           predigest_product_12_50_port, A(49) => 
                           predigest_product_12_49_port, A(48) => 
                           predigest_product_12_48_port, A(47) => 
                           predigest_product_12_47_port, A(46) => 
                           predigest_product_12_46_port, A(45) => 
                           predigest_product_12_45_port, A(44) => 
                           predigest_product_12_44_port, A(43) => 
                           predigest_product_12_43_port, A(42) => 
                           predigest_product_12_42_port, A(41) => 
                           predigest_product_12_41_port, A(40) => 
                           predigest_product_12_40_port, A(39) => 
                           predigest_product_12_39_port, A(38) => 
                           predigest_product_12_38_port, A(37) => 
                           predigest_product_12_37_port, A(36) => 
                           predigest_product_12_36_port, A(35) => 
                           predigest_product_12_35_port, A(34) => 
                           predigest_product_12_34_port, A(33) => 
                           predigest_product_12_33_port, A(32) => 
                           predigest_product_12_32_port, A(31) => 
                           predigest_product_12_31_port, A(30) => 
                           predigest_product_12_30_port, A(29) => 
                           predigest_product_12_29_port, A(28) => 
                           predigest_product_12_28_port, A(27) => 
                           predigest_product_12_27_port, A(26) => 
                           predigest_product_12_26_port, A(25) => 
                           predigest_product_12_25_port, A(24) => 
                           predigest_product_12_24_port, A(23) => 
                           predigest_product_12_23_port, A(22) => 
                           predigest_product_12_22_port, A(21) => 
                           predigest_product_12_21_port, A(20) => 
                           predigest_product_12_20_port, A(19) => 
                           predigest_product_12_19_port, A(18) => 
                           predigest_product_12_18_port, A(17) => 
                           predigest_product_12_17_port, A(16) => 
                           predigest_product_12_16_port, A(15) => 
                           predigest_product_12_15_port, A(14) => 
                           predigest_product_12_14_port, A(13) => 
                           predigest_product_12_13_port, A(12) => 
                           predigest_product_12_12_port, A(11) => 
                           predigest_product_12_11_port, A(10) => 
                           predigest_product_12_10_port, A(9) => 
                           predigest_product_12_9_port, A(8) => 
                           predigest_product_12_8_port, A(7) => 
                           predigest_product_12_7_port, A(6) => 
                           predigest_product_12_6_port, A(5) => 
                           predigest_product_12_5_port, A(4) => 
                           predigest_product_12_4_port, A(3) => 
                           predigest_product_12_3_port, A(2) => 
                           predigest_product_12_2_port, A(1) => 
                           predigest_product_12_1_port, A(0) => 
                           predigest_product_12_0_port, B(63) => 
                           out_imux_13_63_port, B(62) => out_imux_13_62_port, 
                           B(61) => out_imux_13_61_port, B(60) => 
                           out_imux_13_60_port, B(59) => out_imux_13_59_port, 
                           B(58) => out_imux_13_58_port, B(57) => 
                           out_imux_13_57_port, B(56) => out_imux_13_56_port, 
                           B(55) => out_imux_13_55_port, B(54) => 
                           out_imux_13_54_port, B(53) => out_imux_13_53_port, 
                           B(52) => out_imux_13_52_port, B(51) => 
                           out_imux_13_51_port, B(50) => out_imux_13_50_port, 
                           B(49) => out_imux_13_49_port, B(48) => 
                           out_imux_13_48_port, B(47) => out_imux_13_47_port, 
                           B(46) => out_imux_13_46_port, B(45) => 
                           out_imux_13_45_port, B(44) => out_imux_13_44_port, 
                           B(43) => out_imux_13_43_port, B(42) => 
                           out_imux_13_42_port, B(41) => out_imux_13_41_port, 
                           B(40) => out_imux_13_40_port, B(39) => 
                           out_imux_13_39_port, B(38) => out_imux_13_38_port, 
                           B(37) => out_imux_13_37_port, B(36) => 
                           out_imux_13_36_port, B(35) => out_imux_13_35_port, 
                           B(34) => out_imux_13_34_port, B(33) => 
                           out_imux_13_33_port, B(32) => out_imux_13_32_port, 
                           B(31) => out_imux_13_31_port, B(30) => 
                           out_imux_13_30_port, B(29) => out_imux_13_29_port, 
                           B(28) => out_imux_13_28_port, B(27) => 
                           out_imux_13_27_port, B(26) => out_imux_13_26_port, 
                           B(25) => out_imux_13_25_port, B(24) => 
                           out_imux_13_24_port, B(23) => out_imux_13_23_port, 
                           B(22) => out_imux_13_22_port, B(21) => 
                           out_imux_13_21_port, B(20) => out_imux_13_20_port, 
                           B(19) => out_imux_13_19_port, B(18) => 
                           out_imux_13_18_port, B(17) => out_imux_13_17_port, 
                           B(16) => out_imux_13_16_port, B(15) => 
                           out_imux_13_15_port, B(14) => out_imux_13_14_port, 
                           B(13) => out_imux_13_13_port, B(12) => 
                           out_imux_13_12_port, B(11) => out_imux_13_11_port, 
                           B(10) => out_imux_13_10_port, B(9) => 
                           out_imux_13_9_port, B(8) => out_imux_13_8_port, B(7)
                           => out_imux_13_7_port, B(6) => out_imux_13_6_port, 
                           B(5) => out_imux_13_5_port, B(4) => 
                           out_imux_13_4_port, B(3) => out_imux_13_3_port, B(2)
                           => out_imux_13_2_port, B(1) => out_imux_13_1_port, 
                           B(0) => out_imux_13_0_port, Ci => X_Logic0_port, 
                           S(63) => predigest_product_13_63_port, S(62) => 
                           predigest_product_13_62_port, S(61) => 
                           predigest_product_13_61_port, S(60) => 
                           predigest_product_13_60_port, S(59) => 
                           predigest_product_13_59_port, S(58) => 
                           predigest_product_13_58_port, S(57) => 
                           predigest_product_13_57_port, S(56) => 
                           predigest_product_13_56_port, S(55) => 
                           predigest_product_13_55_port, S(54) => 
                           predigest_product_13_54_port, S(53) => 
                           predigest_product_13_53_port, S(52) => 
                           predigest_product_13_52_port, S(51) => 
                           predigest_product_13_51_port, S(50) => 
                           predigest_product_13_50_port, S(49) => 
                           predigest_product_13_49_port, S(48) => 
                           predigest_product_13_48_port, S(47) => 
                           predigest_product_13_47_port, S(46) => 
                           predigest_product_13_46_port, S(45) => 
                           predigest_product_13_45_port, S(44) => 
                           predigest_product_13_44_port, S(43) => 
                           predigest_product_13_43_port, S(42) => 
                           predigest_product_13_42_port, S(41) => 
                           predigest_product_13_41_port, S(40) => 
                           predigest_product_13_40_port, S(39) => 
                           predigest_product_13_39_port, S(38) => 
                           predigest_product_13_38_port, S(37) => 
                           predigest_product_13_37_port, S(36) => 
                           predigest_product_13_36_port, S(35) => 
                           predigest_product_13_35_port, S(34) => 
                           predigest_product_13_34_port, S(33) => 
                           predigest_product_13_33_port, S(32) => 
                           predigest_product_13_32_port, S(31) => 
                           predigest_product_13_31_port, S(30) => 
                           predigest_product_13_30_port, S(29) => 
                           predigest_product_13_29_port, S(28) => 
                           predigest_product_13_28_port, S(27) => 
                           predigest_product_13_27_port, S(26) => 
                           predigest_product_13_26_port, S(25) => 
                           predigest_product_13_25_port, S(24) => 
                           predigest_product_13_24_port, S(23) => 
                           predigest_product_13_23_port, S(22) => 
                           predigest_product_13_22_port, S(21) => 
                           predigest_product_13_21_port, S(20) => 
                           predigest_product_13_20_port, S(19) => 
                           predigest_product_13_19_port, S(18) => 
                           predigest_product_13_18_port, S(17) => 
                           predigest_product_13_17_port, S(16) => 
                           predigest_product_13_16_port, S(15) => 
                           predigest_product_13_15_port, S(14) => 
                           predigest_product_13_14_port, S(13) => 
                           predigest_product_13_13_port, S(12) => 
                           predigest_product_13_12_port, S(11) => 
                           predigest_product_13_11_port, S(10) => 
                           predigest_product_13_10_port, S(9) => 
                           predigest_product_13_9_port, S(8) => 
                           predigest_product_13_8_port, S(7) => 
                           predigest_product_13_7_port, S(6) => 
                           predigest_product_13_6_port, S(5) => 
                           predigest_product_13_5_port, S(4) => 
                           predigest_product_13_4_port, S(3) => 
                           predigest_product_13_3_port, S(2) => 
                           predigest_product_13_2_port, S(1) => 
                           predigest_product_13_1_port, S(0) => 
                           predigest_product_13_0_port, Co => n_1104);
   ENC_i_14 : BOOTH_ENCODER_3BIT_6 port map( B(2) => B(29), B(1) => B(28), B(0)
                           => B(27), ENCODED(2) => 
                           muxs_encoded_signals_14_2_port, ENCODED(1) => 
                           muxs_encoded_signals_14_1_port, ENCODED(0) => 
                           muxs_encoded_signals_14_0_port);
   MUX_i_14 : MUX51_GENERIC_NBIT64_2 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(31), 
                           IN1(59) => A(31), IN1(58) => A(30), IN1(57) => A(29)
                           , IN1(56) => A(28), IN1(55) => A(27), IN1(54) => 
                           A(26), IN1(53) => A(25), IN1(52) => A(24), IN1(51) 
                           => A(23), IN1(50) => A(22), IN1(49) => A(21), 
                           IN1(48) => A(20), IN1(47) => A(19), IN1(46) => A(18)
                           , IN1(45) => A(17), IN1(44) => A(16), IN1(43) => 
                           A(15), IN1(42) => A(14), IN1(41) => A(13), IN1(40) 
                           => A(12), IN1(39) => A(11), IN1(38) => A(10), 
                           IN1(37) => A(9), IN1(36) => A(8), IN1(35) => A(7), 
                           IN1(34) => A(6), IN1(33) => A(5), IN1(32) => A(4), 
                           IN1(31) => A(3), IN1(30) => A(2), IN1(29) => A(1), 
                           IN1(28) => A(0), IN1(27) => X_Logic0_port, IN1(26) 
                           => X_Logic0_port, IN1(25) => X_Logic0_port, IN1(24) 
                           => X_Logic0_port, IN1(23) => X_Logic0_port, IN1(22) 
                           => X_Logic0_port, IN1(21) => X_Logic0_port, IN1(20) 
                           => X_Logic0_port, IN1(19) => X_Logic0_port, IN1(18) 
                           => X_Logic0_port, IN1(17) => X_Logic0_port, IN1(16) 
                           => X_Logic0_port, IN1(15) => X_Logic0_port, IN1(14) 
                           => X_Logic0_port, IN1(13) => X_Logic0_port, IN1(12) 
                           => X_Logic0_port, IN1(11) => X_Logic0_port, IN1(10) 
                           => X_Logic0_port, IN1(9) => X_Logic0_port, IN1(8) =>
                           X_Logic0_port, IN1(7) => X_Logic0_port, IN1(6) => 
                           X_Logic0_port, IN1(5) => X_Logic0_port, IN1(4) => 
                           X_Logic0_port, IN1(3) => X_Logic0_port, IN1(2) => 
                           X_Logic0_port, IN1(1) => X_Logic0_port, IN1(0) => 
                           X_Logic0_port, IN2(63) => negative_a_35_port, 
                           IN2(62) => negative_a_34_port, IN2(61) => n38, 
                           IN2(60) => n35, IN2(59) => negative_a_31_port, 
                           IN2(58) => negative_a_30_port, IN2(57) => 
                           negative_a_29_port, IN2(56) => negative_a_28_port, 
                           IN2(55) => negative_a_27_port, IN2(54) => 
                           negative_a_26_port, IN2(53) => negative_a_25_port, 
                           IN2(52) => negative_a_24_port, IN2(51) => 
                           negative_a_23_port, IN2(50) => negative_a_22_port, 
                           IN2(49) => negative_a_21_port, IN2(48) => 
                           negative_a_20_port, IN2(47) => negative_a_19_port, 
                           IN2(46) => negative_a_18_port, IN2(45) => 
                           negative_a_17_port, IN2(44) => negative_a_16_port, 
                           IN2(43) => negative_a_15_port, IN2(42) => 
                           negative_a_14_port, IN2(41) => negative_a_13_port, 
                           IN2(40) => negative_a_12_port, IN2(39) => 
                           negative_a_11_port, IN2(38) => negative_a_10_port, 
                           IN2(37) => negative_a_9_port, IN2(36) => 
                           negative_a_8_port, IN2(35) => negative_a_7_port, 
                           IN2(34) => negative_a_6_port, IN2(33) => 
                           negative_a_5_port, IN2(32) => negative_a_4_port, 
                           IN2(31) => negative_a_3_port, IN2(30) => 
                           negative_a_2_port, IN2(29) => negative_a_1_port, 
                           IN2(28) => negative_a_0_port, IN2(27) => 
                           X_Logic0_port, IN2(26) => X_Logic0_port, IN2(25) => 
                           X_Logic0_port, IN2(24) => X_Logic0_port, IN2(23) => 
                           X_Logic0_port, IN2(22) => X_Logic0_port, IN2(21) => 
                           X_Logic0_port, IN2(20) => X_Logic0_port, IN2(19) => 
                           X_Logic0_port, IN2(18) => X_Logic0_port, IN2(17) => 
                           X_Logic0_port, IN2(16) => X_Logic0_port, IN2(15) => 
                           X_Logic0_port, IN2(14) => X_Logic0_port, IN2(13) => 
                           X_Logic0_port, IN2(12) => X_Logic0_port, IN2(11) => 
                           X_Logic0_port, IN2(10) => X_Logic0_port, IN2(9) => 
                           X_Logic0_port, IN2(8) => X_Logic0_port, IN2(7) => 
                           X_Logic0_port, IN2(6) => X_Logic0_port, IN2(5) => 
                           X_Logic0_port, IN2(4) => X_Logic0_port, IN2(3) => 
                           X_Logic0_port, IN2(2) => X_Logic0_port, IN2(1) => 
                           X_Logic0_port, IN2(0) => X_Logic0_port, IN3(63) => 
                           A(31), IN3(62) => A(31), IN3(61) => A(31), IN3(60) 
                           => A(31), IN3(59) => A(30), IN3(58) => A(29), 
                           IN3(57) => A(28), IN3(56) => A(27), IN3(55) => A(26)
                           , IN3(54) => A(25), IN3(53) => A(24), IN3(52) => 
                           A(23), IN3(51) => A(22), IN3(50) => A(21), IN3(49) 
                           => A(20), IN3(48) => A(19), IN3(47) => A(18), 
                           IN3(46) => A(17), IN3(45) => A(16), IN3(44) => A(15)
                           , IN3(43) => A(14), IN3(42) => A(13), IN3(41) => 
                           A(12), IN3(40) => A(11), IN3(39) => A(10), IN3(38) 
                           => A(9), IN3(37) => A(8), IN3(36) => A(7), IN3(35) 
                           => A(6), IN3(34) => A(5), IN3(33) => A(4), IN3(32) 
                           => A(3), IN3(31) => A(2), IN3(30) => A(1), IN3(29) 
                           => A(0), IN3(28) => X_Logic0_port, IN3(27) => 
                           X_Logic0_port, IN3(26) => X_Logic0_port, IN3(25) => 
                           X_Logic0_port, IN3(24) => X_Logic0_port, IN3(23) => 
                           X_Logic0_port, IN3(22) => X_Logic0_port, IN3(21) => 
                           X_Logic0_port, IN3(20) => X_Logic0_port, IN3(19) => 
                           X_Logic0_port, IN3(18) => X_Logic0_port, IN3(17) => 
                           X_Logic0_port, IN3(16) => X_Logic0_port, IN3(15) => 
                           X_Logic0_port, IN3(14) => X_Logic0_port, IN3(13) => 
                           X_Logic0_port, IN3(12) => X_Logic0_port, IN3(11) => 
                           X_Logic0_port, IN3(10) => X_Logic0_port, IN3(9) => 
                           X_Logic0_port, IN3(8) => X_Logic0_port, IN3(7) => 
                           X_Logic0_port, IN3(6) => X_Logic0_port, IN3(5) => 
                           X_Logic0_port, IN3(4) => X_Logic0_port, IN3(3) => 
                           X_Logic0_port, IN3(2) => X_Logic0_port, IN3(1) => 
                           X_Logic0_port, IN3(0) => X_Logic0_port, IN4(63) => 
                           negative_a_34_port, IN4(62) => n38, IN4(61) => n35, 
                           IN4(60) => negative_a_31_port, IN4(59) => 
                           negative_a_30_port, IN4(58) => negative_a_29_port, 
                           IN4(57) => negative_a_28_port, IN4(56) => 
                           negative_a_27_port, IN4(55) => negative_a_26_port, 
                           IN4(54) => negative_a_25_port, IN4(53) => 
                           negative_a_24_port, IN4(52) => negative_a_23_port, 
                           IN4(51) => negative_a_22_port, IN4(50) => 
                           negative_a_21_port, IN4(49) => negative_a_20_port, 
                           IN4(48) => negative_a_19_port, IN4(47) => 
                           negative_a_18_port, IN4(46) => negative_a_17_port, 
                           IN4(45) => negative_a_16_port, IN4(44) => 
                           negative_a_15_port, IN4(43) => negative_a_14_port, 
                           IN4(42) => negative_a_13_port, IN4(41) => 
                           negative_a_12_port, IN4(40) => negative_a_11_port, 
                           IN4(39) => negative_a_10_port, IN4(38) => 
                           negative_a_9_port, IN4(37) => negative_a_8_port, 
                           IN4(36) => negative_a_7_port, IN4(35) => 
                           negative_a_6_port, IN4(34) => negative_a_5_port, 
                           IN4(33) => negative_a_4_port, IN4(32) => 
                           negative_a_3_port, IN4(31) => negative_a_2_port, 
                           IN4(30) => negative_a_1_port, IN4(29) => 
                           negative_a_0_port, IN4(28) => X_Logic0_port, IN4(27)
                           => X_Logic0_port, IN4(26) => X_Logic0_port, IN4(25) 
                           => X_Logic0_port, IN4(24) => X_Logic0_port, IN4(23) 
                           => X_Logic0_port, IN4(22) => X_Logic0_port, IN4(21) 
                           => X_Logic0_port, IN4(20) => X_Logic0_port, IN4(19) 
                           => X_Logic0_port, IN4(18) => X_Logic0_port, IN4(17) 
                           => X_Logic0_port, IN4(16) => X_Logic0_port, IN4(15) 
                           => X_Logic0_port, IN4(14) => X_Logic0_port, IN4(13) 
                           => X_Logic0_port, IN4(12) => X_Logic0_port, IN4(11) 
                           => X_Logic0_port, IN4(10) => X_Logic0_port, IN4(9) 
                           => X_Logic0_port, IN4(8) => X_Logic0_port, IN4(7) =>
                           X_Logic0_port, IN4(6) => X_Logic0_port, IN4(5) => 
                           X_Logic0_port, IN4(4) => X_Logic0_port, IN4(3) => 
                           X_Logic0_port, IN4(2) => X_Logic0_port, IN4(1) => 
                           X_Logic0_port, IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_14_2_port, S(1) => 
                           muxs_encoded_signals_14_1_port, S(0) => 
                           muxs_encoded_signals_14_0_port, O(63) => 
                           out_imux_14_63_port, O(62) => out_imux_14_62_port, 
                           O(61) => out_imux_14_61_port, O(60) => 
                           out_imux_14_60_port, O(59) => out_imux_14_59_port, 
                           O(58) => out_imux_14_58_port, O(57) => 
                           out_imux_14_57_port, O(56) => out_imux_14_56_port, 
                           O(55) => out_imux_14_55_port, O(54) => 
                           out_imux_14_54_port, O(53) => out_imux_14_53_port, 
                           O(52) => out_imux_14_52_port, O(51) => 
                           out_imux_14_51_port, O(50) => out_imux_14_50_port, 
                           O(49) => out_imux_14_49_port, O(48) => 
                           out_imux_14_48_port, O(47) => out_imux_14_47_port, 
                           O(46) => out_imux_14_46_port, O(45) => 
                           out_imux_14_45_port, O(44) => out_imux_14_44_port, 
                           O(43) => out_imux_14_43_port, O(42) => 
                           out_imux_14_42_port, O(41) => out_imux_14_41_port, 
                           O(40) => out_imux_14_40_port, O(39) => 
                           out_imux_14_39_port, O(38) => out_imux_14_38_port, 
                           O(37) => out_imux_14_37_port, O(36) => 
                           out_imux_14_36_port, O(35) => out_imux_14_35_port, 
                           O(34) => out_imux_14_34_port, O(33) => 
                           out_imux_14_33_port, O(32) => out_imux_14_32_port, 
                           O(31) => out_imux_14_31_port, O(30) => 
                           out_imux_14_30_port, O(29) => out_imux_14_29_port, 
                           O(28) => out_imux_14_28_port, O(27) => 
                           out_imux_14_27_port, O(26) => out_imux_14_26_port, 
                           O(25) => out_imux_14_25_port, O(24) => 
                           out_imux_14_24_port, O(23) => out_imux_14_23_port, 
                           O(22) => out_imux_14_22_port, O(21) => 
                           out_imux_14_21_port, O(20) => out_imux_14_20_port, 
                           O(19) => out_imux_14_19_port, O(18) => 
                           out_imux_14_18_port, O(17) => out_imux_14_17_port, 
                           O(16) => out_imux_14_16_port, O(15) => 
                           out_imux_14_15_port, O(14) => out_imux_14_14_port, 
                           O(13) => out_imux_14_13_port, O(12) => 
                           out_imux_14_12_port, O(11) => out_imux_14_11_port, 
                           O(10) => out_imux_14_10_port, O(9) => 
                           out_imux_14_9_port, O(8) => out_imux_14_8_port, O(7)
                           => out_imux_14_7_port, O(6) => out_imux_14_6_port, 
                           O(5) => out_imux_14_5_port, O(4) => 
                           out_imux_14_4_port, O(3) => out_imux_14_3_port, O(2)
                           => out_imux_14_2_port, O(1) => out_imux_14_1_port, 
                           O(0) => out_imux_14_0_port);
   ADD64_i_14 : RCA_GENERIC_NBIT64_2 port map( A(63) => 
                           predigest_product_13_63_port, A(62) => 
                           predigest_product_13_62_port, A(61) => 
                           predigest_product_13_61_port, A(60) => 
                           predigest_product_13_60_port, A(59) => 
                           predigest_product_13_59_port, A(58) => 
                           predigest_product_13_58_port, A(57) => 
                           predigest_product_13_57_port, A(56) => 
                           predigest_product_13_56_port, A(55) => 
                           predigest_product_13_55_port, A(54) => 
                           predigest_product_13_54_port, A(53) => 
                           predigest_product_13_53_port, A(52) => 
                           predigest_product_13_52_port, A(51) => 
                           predigest_product_13_51_port, A(50) => 
                           predigest_product_13_50_port, A(49) => 
                           predigest_product_13_49_port, A(48) => 
                           predigest_product_13_48_port, A(47) => 
                           predigest_product_13_47_port, A(46) => 
                           predigest_product_13_46_port, A(45) => 
                           predigest_product_13_45_port, A(44) => 
                           predigest_product_13_44_port, A(43) => 
                           predigest_product_13_43_port, A(42) => 
                           predigest_product_13_42_port, A(41) => 
                           predigest_product_13_41_port, A(40) => 
                           predigest_product_13_40_port, A(39) => 
                           predigest_product_13_39_port, A(38) => 
                           predigest_product_13_38_port, A(37) => 
                           predigest_product_13_37_port, A(36) => 
                           predigest_product_13_36_port, A(35) => 
                           predigest_product_13_35_port, A(34) => 
                           predigest_product_13_34_port, A(33) => 
                           predigest_product_13_33_port, A(32) => 
                           predigest_product_13_32_port, A(31) => 
                           predigest_product_13_31_port, A(30) => 
                           predigest_product_13_30_port, A(29) => 
                           predigest_product_13_29_port, A(28) => 
                           predigest_product_13_28_port, A(27) => 
                           predigest_product_13_27_port, A(26) => 
                           predigest_product_13_26_port, A(25) => 
                           predigest_product_13_25_port, A(24) => 
                           predigest_product_13_24_port, A(23) => 
                           predigest_product_13_23_port, A(22) => 
                           predigest_product_13_22_port, A(21) => 
                           predigest_product_13_21_port, A(20) => 
                           predigest_product_13_20_port, A(19) => 
                           predigest_product_13_19_port, A(18) => 
                           predigest_product_13_18_port, A(17) => 
                           predigest_product_13_17_port, A(16) => 
                           predigest_product_13_16_port, A(15) => 
                           predigest_product_13_15_port, A(14) => 
                           predigest_product_13_14_port, A(13) => 
                           predigest_product_13_13_port, A(12) => 
                           predigest_product_13_12_port, A(11) => 
                           predigest_product_13_11_port, A(10) => 
                           predigest_product_13_10_port, A(9) => 
                           predigest_product_13_9_port, A(8) => 
                           predigest_product_13_8_port, A(7) => 
                           predigest_product_13_7_port, A(6) => 
                           predigest_product_13_6_port, A(5) => 
                           predigest_product_13_5_port, A(4) => 
                           predigest_product_13_4_port, A(3) => 
                           predigest_product_13_3_port, A(2) => 
                           predigest_product_13_2_port, A(1) => 
                           predigest_product_13_1_port, A(0) => 
                           predigest_product_13_0_port, B(63) => 
                           out_imux_14_63_port, B(62) => out_imux_14_62_port, 
                           B(61) => out_imux_14_61_port, B(60) => 
                           out_imux_14_60_port, B(59) => out_imux_14_59_port, 
                           B(58) => out_imux_14_58_port, B(57) => 
                           out_imux_14_57_port, B(56) => out_imux_14_56_port, 
                           B(55) => out_imux_14_55_port, B(54) => 
                           out_imux_14_54_port, B(53) => out_imux_14_53_port, 
                           B(52) => out_imux_14_52_port, B(51) => 
                           out_imux_14_51_port, B(50) => out_imux_14_50_port, 
                           B(49) => out_imux_14_49_port, B(48) => 
                           out_imux_14_48_port, B(47) => out_imux_14_47_port, 
                           B(46) => out_imux_14_46_port, B(45) => 
                           out_imux_14_45_port, B(44) => out_imux_14_44_port, 
                           B(43) => out_imux_14_43_port, B(42) => 
                           out_imux_14_42_port, B(41) => out_imux_14_41_port, 
                           B(40) => out_imux_14_40_port, B(39) => 
                           out_imux_14_39_port, B(38) => out_imux_14_38_port, 
                           B(37) => out_imux_14_37_port, B(36) => 
                           out_imux_14_36_port, B(35) => out_imux_14_35_port, 
                           B(34) => out_imux_14_34_port, B(33) => 
                           out_imux_14_33_port, B(32) => out_imux_14_32_port, 
                           B(31) => out_imux_14_31_port, B(30) => 
                           out_imux_14_30_port, B(29) => out_imux_14_29_port, 
                           B(28) => out_imux_14_28_port, B(27) => 
                           out_imux_14_27_port, B(26) => out_imux_14_26_port, 
                           B(25) => out_imux_14_25_port, B(24) => 
                           out_imux_14_24_port, B(23) => out_imux_14_23_port, 
                           B(22) => out_imux_14_22_port, B(21) => 
                           out_imux_14_21_port, B(20) => out_imux_14_20_port, 
                           B(19) => out_imux_14_19_port, B(18) => 
                           out_imux_14_18_port, B(17) => out_imux_14_17_port, 
                           B(16) => out_imux_14_16_port, B(15) => 
                           out_imux_14_15_port, B(14) => out_imux_14_14_port, 
                           B(13) => out_imux_14_13_port, B(12) => 
                           out_imux_14_12_port, B(11) => out_imux_14_11_port, 
                           B(10) => out_imux_14_10_port, B(9) => 
                           out_imux_14_9_port, B(8) => out_imux_14_8_port, B(7)
                           => out_imux_14_7_port, B(6) => out_imux_14_6_port, 
                           B(5) => out_imux_14_5_port, B(4) => 
                           out_imux_14_4_port, B(3) => out_imux_14_3_port, B(2)
                           => out_imux_14_2_port, B(1) => out_imux_14_1_port, 
                           B(0) => out_imux_14_0_port, Ci => X_Logic0_port, 
                           S(63) => predigest_product_14_63_port, S(62) => 
                           predigest_product_14_62_port, S(61) => 
                           predigest_product_14_61_port, S(60) => 
                           predigest_product_14_60_port, S(59) => 
                           predigest_product_14_59_port, S(58) => 
                           predigest_product_14_58_port, S(57) => 
                           predigest_product_14_57_port, S(56) => 
                           predigest_product_14_56_port, S(55) => 
                           predigest_product_14_55_port, S(54) => 
                           predigest_product_14_54_port, S(53) => 
                           predigest_product_14_53_port, S(52) => 
                           predigest_product_14_52_port, S(51) => 
                           predigest_product_14_51_port, S(50) => 
                           predigest_product_14_50_port, S(49) => 
                           predigest_product_14_49_port, S(48) => 
                           predigest_product_14_48_port, S(47) => 
                           predigest_product_14_47_port, S(46) => 
                           predigest_product_14_46_port, S(45) => 
                           predigest_product_14_45_port, S(44) => 
                           predigest_product_14_44_port, S(43) => 
                           predigest_product_14_43_port, S(42) => 
                           predigest_product_14_42_port, S(41) => 
                           predigest_product_14_41_port, S(40) => 
                           predigest_product_14_40_port, S(39) => 
                           predigest_product_14_39_port, S(38) => 
                           predigest_product_14_38_port, S(37) => 
                           predigest_product_14_37_port, S(36) => 
                           predigest_product_14_36_port, S(35) => 
                           predigest_product_14_35_port, S(34) => 
                           predigest_product_14_34_port, S(33) => 
                           predigest_product_14_33_port, S(32) => 
                           predigest_product_14_32_port, S(31) => 
                           predigest_product_14_31_port, S(30) => 
                           predigest_product_14_30_port, S(29) => 
                           predigest_product_14_29_port, S(28) => 
                           predigest_product_14_28_port, S(27) => 
                           predigest_product_14_27_port, S(26) => 
                           predigest_product_14_26_port, S(25) => 
                           predigest_product_14_25_port, S(24) => 
                           predigest_product_14_24_port, S(23) => 
                           predigest_product_14_23_port, S(22) => 
                           predigest_product_14_22_port, S(21) => 
                           predigest_product_14_21_port, S(20) => 
                           predigest_product_14_20_port, S(19) => 
                           predigest_product_14_19_port, S(18) => 
                           predigest_product_14_18_port, S(17) => 
                           predigest_product_14_17_port, S(16) => 
                           predigest_product_14_16_port, S(15) => 
                           predigest_product_14_15_port, S(14) => 
                           predigest_product_14_14_port, S(13) => 
                           predigest_product_14_13_port, S(12) => 
                           predigest_product_14_12_port, S(11) => 
                           predigest_product_14_11_port, S(10) => 
                           predigest_product_14_10_port, S(9) => 
                           predigest_product_14_9_port, S(8) => 
                           predigest_product_14_8_port, S(7) => 
                           predigest_product_14_7_port, S(6) => 
                           predigest_product_14_6_port, S(5) => 
                           predigest_product_14_5_port, S(4) => 
                           predigest_product_14_4_port, S(3) => 
                           predigest_product_14_3_port, S(2) => 
                           predigest_product_14_2_port, S(1) => 
                           predigest_product_14_1_port, S(0) => 
                           predigest_product_14_0_port, Co => n_1105);
   ENC_i_15 : BOOTH_ENCODER_3BIT_5 port map( B(2) => B(31), B(1) => B(30), B(0)
                           => B(29), ENCODED(2) => 
                           muxs_encoded_signals_15_2_port, ENCODED(1) => 
                           muxs_encoded_signals_15_1_port, ENCODED(0) => 
                           muxs_encoded_signals_15_0_port);
   MUX_i_15 : MUX51_GENERIC_NBIT64_1 port map( IN0(63) => X_Logic0_port, 
                           IN0(62) => X_Logic0_port, IN0(61) => X_Logic0_port, 
                           IN0(60) => X_Logic0_port, IN0(59) => X_Logic0_port, 
                           IN0(58) => X_Logic0_port, IN0(57) => X_Logic0_port, 
                           IN0(56) => X_Logic0_port, IN0(55) => X_Logic0_port, 
                           IN0(54) => X_Logic0_port, IN0(53) => X_Logic0_port, 
                           IN0(52) => X_Logic0_port, IN0(51) => X_Logic0_port, 
                           IN0(50) => X_Logic0_port, IN0(49) => X_Logic0_port, 
                           IN0(48) => X_Logic0_port, IN0(47) => X_Logic0_port, 
                           IN0(46) => X_Logic0_port, IN0(45) => X_Logic0_port, 
                           IN0(44) => X_Logic0_port, IN0(43) => X_Logic0_port, 
                           IN0(42) => X_Logic0_port, IN0(41) => X_Logic0_port, 
                           IN0(40) => X_Logic0_port, IN0(39) => X_Logic0_port, 
                           IN0(38) => X_Logic0_port, IN0(37) => X_Logic0_port, 
                           IN0(36) => X_Logic0_port, IN0(35) => X_Logic0_port, 
                           IN0(34) => X_Logic0_port, IN0(33) => X_Logic0_port, 
                           IN0(32) => X_Logic0_port, IN0(31) => X_Logic0_port, 
                           IN0(30) => X_Logic0_port, IN0(29) => X_Logic0_port, 
                           IN0(28) => X_Logic0_port, IN0(27) => X_Logic0_port, 
                           IN0(26) => X_Logic0_port, IN0(25) => X_Logic0_port, 
                           IN0(24) => X_Logic0_port, IN0(23) => X_Logic0_port, 
                           IN0(22) => X_Logic0_port, IN0(21) => X_Logic0_port, 
                           IN0(20) => X_Logic0_port, IN0(19) => X_Logic0_port, 
                           IN0(18) => X_Logic0_port, IN0(17) => X_Logic0_port, 
                           IN0(16) => X_Logic0_port, IN0(15) => X_Logic0_port, 
                           IN0(14) => X_Logic0_port, IN0(13) => X_Logic0_port, 
                           IN0(12) => X_Logic0_port, IN0(11) => X_Logic0_port, 
                           IN0(10) => X_Logic0_port, IN0(9) => X_Logic0_port, 
                           IN0(8) => X_Logic0_port, IN0(7) => X_Logic0_port, 
                           IN0(6) => X_Logic0_port, IN0(5) => X_Logic0_port, 
                           IN0(4) => X_Logic0_port, IN0(3) => X_Logic0_port, 
                           IN0(2) => X_Logic0_port, IN0(1) => X_Logic0_port, 
                           IN0(0) => X_Logic0_port, IN1(63) => A(31), IN1(62) 
                           => A(31), IN1(61) => A(31), IN1(60) => A(30), 
                           IN1(59) => A(29), IN1(58) => A(28), IN1(57) => A(27)
                           , IN1(56) => A(26), IN1(55) => A(25), IN1(54) => 
                           A(24), IN1(53) => A(23), IN1(52) => A(22), IN1(51) 
                           => A(21), IN1(50) => A(20), IN1(49) => A(19), 
                           IN1(48) => A(18), IN1(47) => A(17), IN1(46) => A(16)
                           , IN1(45) => A(15), IN1(44) => A(14), IN1(43) => 
                           A(13), IN1(42) => A(12), IN1(41) => A(11), IN1(40) 
                           => A(10), IN1(39) => A(9), IN1(38) => A(8), IN1(37) 
                           => A(7), IN1(36) => A(6), IN1(35) => A(5), IN1(34) 
                           => A(4), IN1(33) => A(3), IN1(32) => A(2), IN1(31) 
                           => A(1), IN1(30) => A(0), IN1(29) => X_Logic0_port, 
                           IN1(28) => X_Logic0_port, IN1(27) => X_Logic0_port, 
                           IN1(26) => X_Logic0_port, IN1(25) => X_Logic0_port, 
                           IN1(24) => X_Logic0_port, IN1(23) => X_Logic0_port, 
                           IN1(22) => X_Logic0_port, IN1(21) => X_Logic0_port, 
                           IN1(20) => X_Logic0_port, IN1(19) => X_Logic0_port, 
                           IN1(18) => X_Logic0_port, IN1(17) => X_Logic0_port, 
                           IN1(16) => X_Logic0_port, IN1(15) => X_Logic0_port, 
                           IN1(14) => X_Logic0_port, IN1(13) => X_Logic0_port, 
                           IN1(12) => X_Logic0_port, IN1(11) => X_Logic0_port, 
                           IN1(10) => X_Logic0_port, IN1(9) => X_Logic0_port, 
                           IN1(8) => X_Logic0_port, IN1(7) => X_Logic0_port, 
                           IN1(6) => X_Logic0_port, IN1(5) => X_Logic0_port, 
                           IN1(4) => X_Logic0_port, IN1(3) => X_Logic0_port, 
                           IN1(2) => X_Logic0_port, IN1(1) => X_Logic0_port, 
                           IN1(0) => X_Logic0_port, IN2(63) => n38, IN2(62) => 
                           n35, IN2(61) => negative_a_31_port, IN2(60) => 
                           negative_a_30_port, IN2(59) => negative_a_29_port, 
                           IN2(58) => negative_a_28_port, IN2(57) => 
                           negative_a_27_port, IN2(56) => negative_a_26_port, 
                           IN2(55) => negative_a_25_port, IN2(54) => 
                           negative_a_24_port, IN2(53) => negative_a_23_port, 
                           IN2(52) => negative_a_22_port, IN2(51) => 
                           negative_a_21_port, IN2(50) => negative_a_20_port, 
                           IN2(49) => negative_a_19_port, IN2(48) => 
                           negative_a_18_port, IN2(47) => negative_a_17_port, 
                           IN2(46) => negative_a_16_port, IN2(45) => 
                           negative_a_15_port, IN2(44) => negative_a_14_port, 
                           IN2(43) => negative_a_13_port, IN2(42) => 
                           negative_a_12_port, IN2(41) => negative_a_11_port, 
                           IN2(40) => negative_a_10_port, IN2(39) => 
                           negative_a_9_port, IN2(38) => negative_a_8_port, 
                           IN2(37) => negative_a_7_port, IN2(36) => 
                           negative_a_6_port, IN2(35) => negative_a_5_port, 
                           IN2(34) => negative_a_4_port, IN2(33) => 
                           negative_a_3_port, IN2(32) => negative_a_2_port, 
                           IN2(31) => negative_a_1_port, IN2(30) => 
                           negative_a_0_port, IN2(29) => X_Logic0_port, IN2(28)
                           => X_Logic0_port, IN2(27) => X_Logic0_port, IN2(26) 
                           => X_Logic0_port, IN2(25) => X_Logic0_port, IN2(24) 
                           => X_Logic0_port, IN2(23) => X_Logic0_port, IN2(22) 
                           => X_Logic0_port, IN2(21) => X_Logic0_port, IN2(20) 
                           => X_Logic0_port, IN2(19) => X_Logic0_port, IN2(18) 
                           => X_Logic0_port, IN2(17) => X_Logic0_port, IN2(16) 
                           => X_Logic0_port, IN2(15) => X_Logic0_port, IN2(14) 
                           => X_Logic0_port, IN2(13) => X_Logic0_port, IN2(12) 
                           => X_Logic0_port, IN2(11) => X_Logic0_port, IN2(10) 
                           => X_Logic0_port, IN2(9) => X_Logic0_port, IN2(8) =>
                           X_Logic0_port, IN2(7) => X_Logic0_port, IN2(6) => 
                           X_Logic0_port, IN2(5) => X_Logic0_port, IN2(4) => 
                           X_Logic0_port, IN2(3) => X_Logic0_port, IN2(2) => 
                           X_Logic0_port, IN2(1) => X_Logic0_port, IN2(0) => 
                           X_Logic0_port, IN3(63) => A(31), IN3(62) => A(31), 
                           IN3(61) => A(30), IN3(60) => A(29), IN3(59) => A(28)
                           , IN3(58) => A(27), IN3(57) => A(26), IN3(56) => 
                           A(25), IN3(55) => A(24), IN3(54) => A(23), IN3(53) 
                           => A(22), IN3(52) => A(21), IN3(51) => A(20), 
                           IN3(50) => A(19), IN3(49) => A(18), IN3(48) => A(17)
                           , IN3(47) => A(16), IN3(46) => A(15), IN3(45) => 
                           A(14), IN3(44) => A(13), IN3(43) => A(12), IN3(42) 
                           => A(11), IN3(41) => A(10), IN3(40) => A(9), IN3(39)
                           => A(8), IN3(38) => A(7), IN3(37) => A(6), IN3(36) 
                           => A(5), IN3(35) => A(4), IN3(34) => A(3), IN3(33) 
                           => A(2), IN3(32) => A(1), IN3(31) => A(0), IN3(30) 
                           => X_Logic0_port, IN3(29) => X_Logic0_port, IN3(28) 
                           => X_Logic0_port, IN3(27) => X_Logic0_port, IN3(26) 
                           => X_Logic0_port, IN3(25) => X_Logic0_port, IN3(24) 
                           => X_Logic0_port, IN3(23) => X_Logic0_port, IN3(22) 
                           => X_Logic0_port, IN3(21) => X_Logic0_port, IN3(20) 
                           => X_Logic0_port, IN3(19) => X_Logic0_port, IN3(18) 
                           => X_Logic0_port, IN3(17) => X_Logic0_port, IN3(16) 
                           => X_Logic0_port, IN3(15) => X_Logic0_port, IN3(14) 
                           => X_Logic0_port, IN3(13) => X_Logic0_port, IN3(12) 
                           => X_Logic0_port, IN3(11) => X_Logic0_port, IN3(10) 
                           => X_Logic0_port, IN3(9) => X_Logic0_port, IN3(8) =>
                           X_Logic0_port, IN3(7) => X_Logic0_port, IN3(6) => 
                           X_Logic0_port, IN3(5) => X_Logic0_port, IN3(4) => 
                           X_Logic0_port, IN3(3) => X_Logic0_port, IN3(2) => 
                           X_Logic0_port, IN3(1) => X_Logic0_port, IN3(0) => 
                           X_Logic0_port, IN4(63) => n35, IN4(62) => 
                           negative_a_31_port, IN4(61) => negative_a_30_port, 
                           IN4(60) => negative_a_29_port, IN4(59) => 
                           negative_a_28_port, IN4(58) => negative_a_27_port, 
                           IN4(57) => negative_a_26_port, IN4(56) => 
                           negative_a_25_port, IN4(55) => negative_a_24_port, 
                           IN4(54) => negative_a_23_port, IN4(53) => 
                           negative_a_22_port, IN4(52) => negative_a_21_port, 
                           IN4(51) => negative_a_20_port, IN4(50) => 
                           negative_a_19_port, IN4(49) => negative_a_18_port, 
                           IN4(48) => negative_a_17_port, IN4(47) => 
                           negative_a_16_port, IN4(46) => negative_a_15_port, 
                           IN4(45) => negative_a_14_port, IN4(44) => 
                           negative_a_13_port, IN4(43) => negative_a_12_port, 
                           IN4(42) => negative_a_11_port, IN4(41) => 
                           negative_a_10_port, IN4(40) => negative_a_9_port, 
                           IN4(39) => negative_a_8_port, IN4(38) => 
                           negative_a_7_port, IN4(37) => negative_a_6_port, 
                           IN4(36) => negative_a_5_port, IN4(35) => 
                           negative_a_4_port, IN4(34) => negative_a_3_port, 
                           IN4(33) => negative_a_2_port, IN4(32) => 
                           negative_a_1_port, IN4(31) => negative_a_0_port, 
                           IN4(30) => X_Logic0_port, IN4(29) => X_Logic0_port, 
                           IN4(28) => X_Logic0_port, IN4(27) => X_Logic0_port, 
                           IN4(26) => X_Logic0_port, IN4(25) => X_Logic0_port, 
                           IN4(24) => X_Logic0_port, IN4(23) => X_Logic0_port, 
                           IN4(22) => X_Logic0_port, IN4(21) => X_Logic0_port, 
                           IN4(20) => X_Logic0_port, IN4(19) => X_Logic0_port, 
                           IN4(18) => X_Logic0_port, IN4(17) => X_Logic0_port, 
                           IN4(16) => X_Logic0_port, IN4(15) => X_Logic0_port, 
                           IN4(14) => X_Logic0_port, IN4(13) => X_Logic0_port, 
                           IN4(12) => X_Logic0_port, IN4(11) => X_Logic0_port, 
                           IN4(10) => X_Logic0_port, IN4(9) => X_Logic0_port, 
                           IN4(8) => X_Logic0_port, IN4(7) => X_Logic0_port, 
                           IN4(6) => X_Logic0_port, IN4(5) => X_Logic0_port, 
                           IN4(4) => X_Logic0_port, IN4(3) => X_Logic0_port, 
                           IN4(2) => X_Logic0_port, IN4(1) => X_Logic0_port, 
                           IN4(0) => X_Logic0_port, S(2) => 
                           muxs_encoded_signals_15_2_port, S(1) => 
                           muxs_encoded_signals_15_1_port, S(0) => 
                           muxs_encoded_signals_15_0_port, O(63) => 
                           out_imux_15_63_port, O(62) => out_imux_15_62_port, 
                           O(61) => out_imux_15_61_port, O(60) => 
                           out_imux_15_60_port, O(59) => out_imux_15_59_port, 
                           O(58) => out_imux_15_58_port, O(57) => 
                           out_imux_15_57_port, O(56) => out_imux_15_56_port, 
                           O(55) => out_imux_15_55_port, O(54) => 
                           out_imux_15_54_port, O(53) => out_imux_15_53_port, 
                           O(52) => out_imux_15_52_port, O(51) => 
                           out_imux_15_51_port, O(50) => out_imux_15_50_port, 
                           O(49) => out_imux_15_49_port, O(48) => 
                           out_imux_15_48_port, O(47) => out_imux_15_47_port, 
                           O(46) => out_imux_15_46_port, O(45) => 
                           out_imux_15_45_port, O(44) => out_imux_15_44_port, 
                           O(43) => out_imux_15_43_port, O(42) => 
                           out_imux_15_42_port, O(41) => out_imux_15_41_port, 
                           O(40) => out_imux_15_40_port, O(39) => 
                           out_imux_15_39_port, O(38) => out_imux_15_38_port, 
                           O(37) => out_imux_15_37_port, O(36) => 
                           out_imux_15_36_port, O(35) => out_imux_15_35_port, 
                           O(34) => out_imux_15_34_port, O(33) => 
                           out_imux_15_33_port, O(32) => out_imux_15_32_port, 
                           O(31) => out_imux_15_31_port, O(30) => 
                           out_imux_15_30_port, O(29) => out_imux_15_29_port, 
                           O(28) => out_imux_15_28_port, O(27) => 
                           out_imux_15_27_port, O(26) => out_imux_15_26_port, 
                           O(25) => out_imux_15_25_port, O(24) => 
                           out_imux_15_24_port, O(23) => out_imux_15_23_port, 
                           O(22) => out_imux_15_22_port, O(21) => 
                           out_imux_15_21_port, O(20) => out_imux_15_20_port, 
                           O(19) => out_imux_15_19_port, O(18) => 
                           out_imux_15_18_port, O(17) => out_imux_15_17_port, 
                           O(16) => out_imux_15_16_port, O(15) => 
                           out_imux_15_15_port, O(14) => out_imux_15_14_port, 
                           O(13) => out_imux_15_13_port, O(12) => 
                           out_imux_15_12_port, O(11) => out_imux_15_11_port, 
                           O(10) => out_imux_15_10_port, O(9) => 
                           out_imux_15_9_port, O(8) => out_imux_15_8_port, O(7)
                           => out_imux_15_7_port, O(6) => out_imux_15_6_port, 
                           O(5) => out_imux_15_5_port, O(4) => 
                           out_imux_15_4_port, O(3) => out_imux_15_3_port, O(2)
                           => out_imux_15_2_port, O(1) => out_imux_15_1_port, 
                           O(0) => out_imux_15_0_port);
   ADD64_i_15 : RCA_GENERIC_NBIT64_1 port map( A(63) => 
                           predigest_product_14_63_port, A(62) => 
                           predigest_product_14_62_port, A(61) => 
                           predigest_product_14_61_port, A(60) => 
                           predigest_product_14_60_port, A(59) => 
                           predigest_product_14_59_port, A(58) => 
                           predigest_product_14_58_port, A(57) => 
                           predigest_product_14_57_port, A(56) => 
                           predigest_product_14_56_port, A(55) => 
                           predigest_product_14_55_port, A(54) => 
                           predigest_product_14_54_port, A(53) => 
                           predigest_product_14_53_port, A(52) => 
                           predigest_product_14_52_port, A(51) => 
                           predigest_product_14_51_port, A(50) => 
                           predigest_product_14_50_port, A(49) => 
                           predigest_product_14_49_port, A(48) => 
                           predigest_product_14_48_port, A(47) => 
                           predigest_product_14_47_port, A(46) => 
                           predigest_product_14_46_port, A(45) => 
                           predigest_product_14_45_port, A(44) => 
                           predigest_product_14_44_port, A(43) => 
                           predigest_product_14_43_port, A(42) => 
                           predigest_product_14_42_port, A(41) => 
                           predigest_product_14_41_port, A(40) => 
                           predigest_product_14_40_port, A(39) => 
                           predigest_product_14_39_port, A(38) => 
                           predigest_product_14_38_port, A(37) => 
                           predigest_product_14_37_port, A(36) => 
                           predigest_product_14_36_port, A(35) => 
                           predigest_product_14_35_port, A(34) => 
                           predigest_product_14_34_port, A(33) => 
                           predigest_product_14_33_port, A(32) => 
                           predigest_product_14_32_port, A(31) => 
                           predigest_product_14_31_port, A(30) => 
                           predigest_product_14_30_port, A(29) => 
                           predigest_product_14_29_port, A(28) => 
                           predigest_product_14_28_port, A(27) => 
                           predigest_product_14_27_port, A(26) => 
                           predigest_product_14_26_port, A(25) => 
                           predigest_product_14_25_port, A(24) => 
                           predigest_product_14_24_port, A(23) => 
                           predigest_product_14_23_port, A(22) => 
                           predigest_product_14_22_port, A(21) => 
                           predigest_product_14_21_port, A(20) => 
                           predigest_product_14_20_port, A(19) => 
                           predigest_product_14_19_port, A(18) => 
                           predigest_product_14_18_port, A(17) => 
                           predigest_product_14_17_port, A(16) => 
                           predigest_product_14_16_port, A(15) => 
                           predigest_product_14_15_port, A(14) => 
                           predigest_product_14_14_port, A(13) => 
                           predigest_product_14_13_port, A(12) => 
                           predigest_product_14_12_port, A(11) => 
                           predigest_product_14_11_port, A(10) => 
                           predigest_product_14_10_port, A(9) => 
                           predigest_product_14_9_port, A(8) => 
                           predigest_product_14_8_port, A(7) => 
                           predigest_product_14_7_port, A(6) => 
                           predigest_product_14_6_port, A(5) => 
                           predigest_product_14_5_port, A(4) => 
                           predigest_product_14_4_port, A(3) => 
                           predigest_product_14_3_port, A(2) => 
                           predigest_product_14_2_port, A(1) => 
                           predigest_product_14_1_port, A(0) => 
                           predigest_product_14_0_port, B(63) => 
                           out_imux_15_63_port, B(62) => out_imux_15_62_port, 
                           B(61) => out_imux_15_61_port, B(60) => 
                           out_imux_15_60_port, B(59) => out_imux_15_59_port, 
                           B(58) => out_imux_15_58_port, B(57) => 
                           out_imux_15_57_port, B(56) => out_imux_15_56_port, 
                           B(55) => out_imux_15_55_port, B(54) => 
                           out_imux_15_54_port, B(53) => out_imux_15_53_port, 
                           B(52) => out_imux_15_52_port, B(51) => 
                           out_imux_15_51_port, B(50) => out_imux_15_50_port, 
                           B(49) => out_imux_15_49_port, B(48) => 
                           out_imux_15_48_port, B(47) => out_imux_15_47_port, 
                           B(46) => out_imux_15_46_port, B(45) => 
                           out_imux_15_45_port, B(44) => out_imux_15_44_port, 
                           B(43) => out_imux_15_43_port, B(42) => 
                           out_imux_15_42_port, B(41) => out_imux_15_41_port, 
                           B(40) => out_imux_15_40_port, B(39) => 
                           out_imux_15_39_port, B(38) => out_imux_15_38_port, 
                           B(37) => out_imux_15_37_port, B(36) => 
                           out_imux_15_36_port, B(35) => out_imux_15_35_port, 
                           B(34) => out_imux_15_34_port, B(33) => 
                           out_imux_15_33_port, B(32) => out_imux_15_32_port, 
                           B(31) => out_imux_15_31_port, B(30) => 
                           out_imux_15_30_port, B(29) => out_imux_15_29_port, 
                           B(28) => out_imux_15_28_port, B(27) => 
                           out_imux_15_27_port, B(26) => out_imux_15_26_port, 
                           B(25) => out_imux_15_25_port, B(24) => 
                           out_imux_15_24_port, B(23) => out_imux_15_23_port, 
                           B(22) => out_imux_15_22_port, B(21) => 
                           out_imux_15_21_port, B(20) => out_imux_15_20_port, 
                           B(19) => out_imux_15_19_port, B(18) => 
                           out_imux_15_18_port, B(17) => out_imux_15_17_port, 
                           B(16) => out_imux_15_16_port, B(15) => 
                           out_imux_15_15_port, B(14) => out_imux_15_14_port, 
                           B(13) => out_imux_15_13_port, B(12) => 
                           out_imux_15_12_port, B(11) => out_imux_15_11_port, 
                           B(10) => out_imux_15_10_port, B(9) => 
                           out_imux_15_9_port, B(8) => out_imux_15_8_port, B(7)
                           => out_imux_15_7_port, B(6) => out_imux_15_6_port, 
                           B(5) => out_imux_15_5_port, B(4) => 
                           out_imux_15_4_port, B(3) => out_imux_15_3_port, B(2)
                           => out_imux_15_2_port, B(1) => out_imux_15_1_port, 
                           B(0) => out_imux_15_0_port, Ci => X_Logic0_port, 
                           S(63) => P(63), S(62) => P(62), S(61) => P(61), 
                           S(60) => P(60), S(59) => P(59), S(58) => P(58), 
                           S(57) => P(57), S(56) => P(56), S(55) => P(55), 
                           S(54) => P(54), S(53) => P(53), S(52) => P(52), 
                           S(51) => P(51), S(50) => P(50), S(49) => P(49), 
                           S(48) => P(48), S(47) => P(47), S(46) => P(46), 
                           S(45) => P(45), S(44) => P(44), S(43) => P(43), 
                           S(42) => P(42), S(41) => P(41), S(40) => P(40), 
                           S(39) => P(39), S(38) => P(38), S(37) => P(37), 
                           S(36) => P(36), S(35) => P(35), S(34) => P(34), 
                           S(33) => P(33), S(32) => P(32), S(31) => P(31), 
                           S(30) => P(30), S(29) => P(29), S(28) => P(28), 
                           S(27) => P(27), S(26) => P(26), S(25) => P(25), 
                           S(24) => P(24), S(23) => P(23), S(22) => P(22), 
                           S(21) => P(21), S(20) => P(20), S(19) => P(19), 
                           S(18) => P(18), S(17) => P(17), S(16) => P(16), 
                           S(15) => P(15), S(14) => P(14), S(13) => P(13), 
                           S(12) => P(12), S(11) => P(11), S(10) => P(10), S(9)
                           => P(9), S(8) => P(8), S(7) => P(7), S(6) => P(6), 
                           S(5) => P(5), S(4) => P(4), S(3) => P(3), S(2) => 
                           P(2), S(1) => P(1), S(0) => P(0), Co => n_1106);
   add_66 : BOOTHMUL_NBIT32_DW01_inc_0 port map( A(63) => n39, A(62) => n39, 
                           A(61) => n39, A(60) => n39, A(59) => n39, A(58) => 
                           n39, A(57) => n39, A(56) => n39, A(55) => n39, A(54)
                           => n39, A(53) => n39, A(52) => n39, A(51) => n39, 
                           A(50) => n39, A(49) => n39, A(48) => n39, A(47) => 
                           n39, A(46) => n39, A(45) => n39, A(44) => n39, A(43)
                           => n39, A(42) => n39, A(41) => n39, A(40) => n39, 
                           A(39) => n39, A(38) => n39, A(37) => n39, A(36) => 
                           n39, A(35) => n39, A(34) => n39, A(33) => n39, A(32)
                           => n39, A(31) => n39, A(30) => n40, A(29) => n41, 
                           A(28) => n42, A(27) => n43, A(26) => n44, A(25) => 
                           n45, A(24) => n46, A(23) => n47, A(22) => n48, A(21)
                           => n49, A(20) => n50, A(19) => n51, A(18) => n52, 
                           A(17) => n53, A(16) => n54, A(15) => n55, A(14) => 
                           n56, A(13) => n57, A(12) => n58, A(11) => n59, A(10)
                           => n60, A(9) => n61, A(8) => n62, A(7) => n63, A(6) 
                           => n64, A(5) => n65, A(4) => n66, A(3) => n67, A(2) 
                           => n68, A(1) => n69, A(0) => n70, SUM(63) => 
                           negative_a_63_port, SUM(62) => negative_a_62_port, 
                           SUM(61) => negative_a_61_port, SUM(60) => 
                           negative_a_60_port, SUM(59) => negative_a_59_port, 
                           SUM(58) => negative_a_58_port, SUM(57) => 
                           negative_a_57_port, SUM(56) => negative_a_56_port, 
                           SUM(55) => negative_a_55_port, SUM(54) => 
                           negative_a_54_port, SUM(53) => negative_a_53_port, 
                           SUM(52) => negative_a_52_port, SUM(51) => 
                           negative_a_51_port, SUM(50) => negative_a_50_port, 
                           SUM(49) => negative_a_49_port, SUM(48) => 
                           negative_a_48_port, SUM(47) => negative_a_47_port, 
                           SUM(46) => negative_a_46_port, SUM(45) => 
                           negative_a_45_port, SUM(44) => negative_a_44_port, 
                           SUM(43) => negative_a_43_port, SUM(42) => 
                           negative_a_42_port, SUM(41) => negative_a_41_port, 
                           SUM(40) => negative_a_40_port, SUM(39) => 
                           negative_a_39_port, SUM(38) => negative_a_38_port, 
                           SUM(37) => negative_a_37_port, SUM(36) => 
                           negative_a_36_port, SUM(35) => negative_a_35_port, 
                           SUM(34) => negative_a_34_port, SUM(33) => 
                           negative_a_33_port, SUM(32) => negative_a_32_port, 
                           SUM(31) => negative_a_31_port, SUM(30) => 
                           negative_a_30_port, SUM(29) => negative_a_29_port, 
                           SUM(28) => negative_a_28_port, SUM(27) => 
                           negative_a_27_port, SUM(26) => negative_a_26_port, 
                           SUM(25) => negative_a_25_port, SUM(24) => 
                           negative_a_24_port, SUM(23) => negative_a_23_port, 
                           SUM(22) => negative_a_22_port, SUM(21) => 
                           negative_a_21_port, SUM(20) => negative_a_20_port, 
                           SUM(19) => negative_a_19_port, SUM(18) => 
                           negative_a_18_port, SUM(17) => negative_a_17_port, 
                           SUM(16) => negative_a_16_port, SUM(15) => 
                           negative_a_15_port, SUM(14) => negative_a_14_port, 
                           SUM(13) => negative_a_13_port, SUM(12) => 
                           negative_a_12_port, SUM(11) => negative_a_11_port, 
                           SUM(10) => negative_a_10_port, SUM(9) => 
                           negative_a_9_port, SUM(8) => negative_a_8_port, 
                           SUM(7) => negative_a_7_port, SUM(6) => 
                           negative_a_6_port, SUM(5) => negative_a_5_port, 
                           SUM(4) => negative_a_4_port, SUM(3) => 
                           negative_a_3_port, SUM(2) => negative_a_2_port, 
                           SUM(1) => negative_a_1_port, SUM(0) => 
                           negative_a_0_port);
   U35 : BUF_X1 port map( A => negative_a_32_port, Z => n33);
   U36 : BUF_X1 port map( A => negative_a_33_port, Z => n36);
   U37 : BUF_X1 port map( A => negative_a_32_port, Z => n34);
   U38 : BUF_X1 port map( A => negative_a_33_port, Z => n37);
   U39 : BUF_X1 port map( A => negative_a_32_port, Z => n35);
   U40 : BUF_X1 port map( A => negative_a_33_port, Z => n38);
   U41 : INV_X1 port map( A => A(31), ZN => n39);
   U42 : INV_X1 port map( A => A(30), ZN => n40);
   U43 : INV_X1 port map( A => A(29), ZN => n41);
   U44 : INV_X1 port map( A => A(28), ZN => n42);
   U45 : INV_X1 port map( A => A(27), ZN => n43);
   U46 : INV_X1 port map( A => A(26), ZN => n44);
   U47 : INV_X1 port map( A => A(25), ZN => n45);
   U48 : INV_X1 port map( A => A(24), ZN => n46);
   U49 : INV_X1 port map( A => A(23), ZN => n47);
   U50 : INV_X1 port map( A => A(22), ZN => n48);
   U51 : INV_X1 port map( A => A(21), ZN => n49);
   U52 : INV_X1 port map( A => A(20), ZN => n50);
   U53 : INV_X1 port map( A => A(19), ZN => n51);
   U54 : INV_X1 port map( A => A(18), ZN => n52);
   U55 : INV_X1 port map( A => A(17), ZN => n53);
   U56 : INV_X1 port map( A => A(16), ZN => n54);
   U57 : INV_X1 port map( A => A(15), ZN => n55);
   U58 : INV_X1 port map( A => A(14), ZN => n56);
   U59 : INV_X1 port map( A => A(13), ZN => n57);
   U60 : INV_X1 port map( A => A(12), ZN => n58);
   U61 : INV_X1 port map( A => A(11), ZN => n59);
   U62 : INV_X1 port map( A => A(10), ZN => n60);
   U63 : INV_X1 port map( A => A(9), ZN => n61);
   U64 : INV_X1 port map( A => A(8), ZN => n62);
   U65 : INV_X1 port map( A => A(7), ZN => n63);
   U66 : INV_X1 port map( A => A(6), ZN => n64);
   U67 : INV_X1 port map( A => A(5), ZN => n65);
   U68 : INV_X1 port map( A => A(4), ZN => n66);
   U69 : INV_X1 port map( A => A(3), ZN => n67);
   U70 : INV_X1 port map( A => A(2), ZN => n68);
   U71 : INV_X1 port map( A => A(1), ZN => n69);
   U72 : INV_X1 port map( A => A(0), ZN => n70);

end SYN_BOOTHMUL_STRUCT;
