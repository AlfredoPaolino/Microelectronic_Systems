
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_RF_generic_ADDR_BIT5_DATA_BIT32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_RF_generic_ADDR_BIT5_DATA_BIT32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_RF_generic_ADDR_BIT5_DATA_BIT32.all;

entity RF_generic_ADDR_BIT5_DATA_BIT32 is

   port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADDR_WR, ADDR_RD1, 
         ADDR_RD2 : in std_logic_vector (4 downto 0);  DATA_IN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_generic_ADDR_BIT5_DATA_BIT32;

architecture SYN_beh of RF_generic_ADDR_BIT5_DATA_BIT32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
      n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
      n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, 
      n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, 
      n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, 
      n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, 
      n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
      n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, 
      n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, 
      n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
      n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
      n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, 
      n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, 
      n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, 
      n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, 
      n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, 
      n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, 
      n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
      n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
      n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
      n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, 
      n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
      n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
      n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, 
      n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
      n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
      n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
      n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, 
      n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
      n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, 
      n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
      n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
      n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
      n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, 
      n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, 
      n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, 
      n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, 
      n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
      n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
      n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
      n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
      n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, 
      n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, 
      n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
      n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
      n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
      n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, 
      n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
      n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, 
      n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, 
      n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, 
      n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
      n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, 
      n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, 
      n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
      n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
      n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, 
      n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, 
      n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, 
      n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
      n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, 
      n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, 
      n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
      n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
      n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
      n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, 
      n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, 
      n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
      n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
      n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, 
      n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, 
      n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
      n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, 
      n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, 
      n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
      n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, 
      n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, 
      n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
      n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, 
      n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
      n6702, n6703, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, 
      n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, 
      n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, 
      n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8893, n8894, n8895, 
      n8896, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, 
      n8910, n8911, n8912, n8913, n8916, n8917, n8918, n8919, n8920, n8921, 
      n8922, n8923, n8924, n8927, n8928, n8929, n8930, n8933, n8934, n8935, 
      n8936, n8937, n8938, n8939, n8940, n8941, n8944, n8945, n8946, n8947, 
      n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8961, 
      n8962, n8963, n8964, n8967, n8968, n8969, n8970, n8971, n8972, n8973, 
      n8974, n8975, n8978, n8979, n8980, n8981, n8984, n8985, n8986, n8987, 
      n8988, n8989, n8990, n8991, n8992, n8995, n8996, n8997, n8998, n9001, 
      n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9012, n9013, 
      n9014, n9015, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9029, n9030, n9031, n9032, n9035, n9036, n9037, n9038, n9039, 
      n9040, n9041, n9042, n9043, n9046, n9047, n9048, n9049, n9052, n9053, 
      n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9063, n9064, n9065, 
      n9066, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, 
      n9080, n9081, n9082, n9083, n9086, n9087, n9088, n9089, n9090, n9091, 
      n9092, n9093, n9094, n9097, n9098, n9099, n9100, n9103, n9104, n9105, 
      n9106, n9107, n9108, n9109, n9110, n9111, n9114, n9115, n9116, n9117, 
      n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9131, 
      n9132, n9133, n9134, n9137, n9138, n9139, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9148, n9149, n9150, n9151, n9154, n9155, n9156, n9157, 
      n9158, n9159, n9160, n9161, n9162, n9165, n9166, n9167, n9168, n9171, 
      n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9182, n9183, 
      n9184, n9185, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, 
      n9196, n9199, n9200, n9201, n9202, n9205, n9206, n9207, n9208, n9209, 
      n9210, n9211, n9212, n9213, n9216, n9217, n9218, n9219, n9222, n9223, 
      n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9233, n9234, n9235, 
      n9236, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, 
      n9250, n9251, n9252, n9253, n9256, n9257, n9258, n9259, n9260, n9261, 
      n9262, n9263, n9264, n9267, n9268, n9269, n9270, n9273, n9274, n9275, 
      n9276, n9277, n9278, n9279, n9280, n9281, n9284, n9285, n9286, n9287, 
      n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9301, 
      n9302, n9303, n9304, n9307, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9318, n9319, n9320, n9321, n9324, n9325, n9326, n9327, 
      n9328, n9329, n9330, n9331, n9332, n9335, n9336, n9337, n9338, n9341, 
      n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9352, n9353, 
      n9354, n9355, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, 
      n9366, n9369, n9370, n9371, n9372, n9375, n9376, n9377, n9378, n9379, 
      n9380, n9381, n9382, n9383, n9386, n9387, n9388, n9389, n9392, n9393, 
      n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9403, n9404, n9405, 
      n9406, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, 
      n9420, n9421, n9422, n9423, n9426, n9427, n9428, n9429, n9430, n9431, 
      n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, 
      n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12674, n12675, 
      n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, 
      n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, 
      n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, 
      n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, 
      n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, 
      n12721, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, 
      n13567, n13568, n13569, n13570, n13571, n13572, n14597, n14598, n14599, 
      n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, 
      n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, 
      n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, 
      n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, 
      n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, 
      n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, 
      n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, 
      n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, 
      n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, 
      n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, 
      n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, 
      n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, 
      n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, 
      n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, 
      n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, 
      n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, 
      n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, 
      n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, 
      n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, 
      n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, 
      n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, 
      n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, 
      n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, 
      n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, 
      n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, 
      n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, 
      n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, 
      n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, 
      n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, 
      n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, 
      n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, 
      n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, 
      n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, 
      n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, 
      n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, 
      n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, 
      n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, 
      n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, 
      n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, 
      n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, 
      n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, 
      n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, 
      n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, 
      n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, 
      n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, 
      n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, 
      n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, 
      n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, 
      n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, 
      n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, 
      n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, 
      n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, 
      n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, 
      n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, 
      n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, 
      n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, 
      n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, 
      n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, 
      n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, 
      n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, 
      n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, 
      n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, 
      n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, 
      n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, 
      n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, 
      n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, 
      n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, 
      n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, 
      n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, 
      n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, 
      n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, 
      n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, 
      n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, 
      n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, 
      n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, 
      n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, 
      n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, 
      n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, 
      n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, 
      n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, 
      n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, 
      n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, 
      n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, 
      n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, 
      n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, 
      n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, 
      n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, 
      n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, 
      n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, 
      n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, 
      n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, 
      n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, 
      n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, 
      n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, 
      n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, 
      n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, 
      n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, 
      n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, 
      n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, 
      n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, 
      n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, 
      n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, 
      n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, 
      n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, 
      n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, 
      n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, 
      n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, 
      n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, 
      n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, 
      n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, 
      n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, 
      n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, 
      n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, 
      n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, 
      n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, 
      n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, 
      n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, 
      n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, 
      n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, 
      n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, 
      n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, 
      n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, 
      n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, 
      n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, 
      n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, 
      n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, 
      n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, 
      n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, 
      n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, 
      n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, 
      n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, 
      n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, 
      n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, 
      n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, 
      n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, 
      n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, 
      n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, 
      n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, 
      n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, 
      n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, 
      n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, 
      n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, 
      n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, 
      n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, 
      n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, 
      n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, 
      n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, 
      n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, 
      n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, 
      n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, 
      n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, 
      n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, 
      n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, 
      n15977, n15978, n15979, n15980, n16493, n16494, n16495, n16496, n16497, 
      n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, 
      n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, 
      n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, 
      n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, 
      n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, 
      n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, 
      n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, 
      n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, 
      n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, 
      n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, 
      n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, 
      n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, 
      n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, 
      n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, 
      n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, 
      n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, 
      n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, 
      n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, 
      n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, 
      n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, 
      n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, 
      n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, 
      n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, 
      n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, 
      n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, 
      n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, 
      n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, 
      n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, 
      n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, 
      n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, 
      n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, 
      n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, 
      n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, 
      n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, 
      n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, 
      n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, 
      n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, 
      n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, 
      n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, 
      n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, 
      n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, 
      n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, 
      n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, 
      n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, 
      n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, 
      n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, 
      n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, 
      n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, 
      n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, 
      n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, 
      n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, 
      n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, 
      n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, 
      n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, 
      n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, 
      n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, 
      n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, 
      n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, 
      n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, 
      n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, 
      n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, 
      n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, 
      n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, 
      n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, 
      n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, 
      n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, 
      n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, 
      n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, 
      n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, 
      n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, 
      n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, 
      n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, 
      n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, 
      n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, 
      n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, 
      n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, 
      n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, 
      n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, 
      n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, 
      n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, 
      n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, 
      n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, 
      n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, 
      n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, 
      n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, 
      n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, 
      n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, 
      n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, 
      n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, 
      n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, 
      n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, 
      n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, 
      n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, 
      n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, 
      n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, 
      n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, 
      n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, 
      n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, 
      n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, 
      n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, 
      n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, 
      n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, 
      n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, 
      n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, 
      n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, 
      n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, 
      n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, 
      n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, 
      n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, 
      n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, 
      n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, 
      n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, 
      n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, 
      n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, 
      n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, 
      n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, 
      n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, 
      n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, 
      n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, 
      n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, 
      n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, 
      n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, 
      n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, 
      n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, 
      n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, 
      n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, 
      n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, 
      n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, 
      n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, 
      n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, 
      n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, 
      n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, 
      n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, 
      n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, 
      n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, 
      n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, 
      n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, 
      n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, 
      n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, 
      n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, 
      n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, 
      n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, 
      n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, 
      n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, 
      n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, 
      n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, 
      n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, 
      n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, 
      n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, 
      n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, 
      n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, 
      n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, 
      n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, 
      n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, 
      n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, 
      n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, 
      n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, 
      n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, 
      n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, 
      n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, 
      n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, 
      n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, 
      n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, 
      n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, 
      n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, 
      n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, 
      n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, 
      n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, 
      n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, 
      n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, 
      n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, 
      n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, 
      n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, 
      n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, 
      n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, 
      n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, 
      n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, 
      n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, 
      n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, 
      n18109, n18110, n18111, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, 
      n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, 
      n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, 
      n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, 
      n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, 
      n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, 
      n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, 
      n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, 
      n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, 
      n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, 
      n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, 
      n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, 
      n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, 
      n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, 
      n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, 
      n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, 
      n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, 
      n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, 
      n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, 
      n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, 
      n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, 
      n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, 
      n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, 
      n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, 
      n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, 
      n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, 
      n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, 
      n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, 
      n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, 
      n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, 
      n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, 
      n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, 
      n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, 
      n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, 
      n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, 
      n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, 
      n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, 
      n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, 
      n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, 
      n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, 
      n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, 
      n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, 
      n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, 
      n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, 
      n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, 
      n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, 
      n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, 
      n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, 
      n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, 
      n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, 
      n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, 
      n_1510, n_1511 : std_logic;

begin
   
   OUT1_reg_31_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => OUT1(31), QN
                           => n8856);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => OUT1(30), QN
                           => n8857);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => OUT1(29), QN
                           => n8858);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => OUT1(28), QN
                           => n8859);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => OUT1(27), QN
                           => n8860);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => OUT1(26), QN
                           => n8861);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => OUT1(25), QN
                           => n8862);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => OUT1(24), QN
                           => n8863);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => OUT1(23), QN
                           => n8864);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => OUT1(22), QN
                           => n8865);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => OUT1(21), QN
                           => n8866);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => OUT1(20), QN
                           => n8867);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => OUT1(19), QN
                           => n8868);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => OUT1(18), QN
                           => n8869);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => OUT1(17), QN
                           => n8870);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => OUT1(16), QN
                           => n8871);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => OUT1(15), QN
                           => n8872);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => OUT1(14), QN
                           => n8873);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => OUT1(13), QN
                           => n8874);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => OUT1(12), QN
                           => n8875);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => OUT1(11), QN
                           => n8876);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => OUT1(10), QN
                           => n8877);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => OUT1(9), QN 
                           => n8878);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => OUT1(8), QN 
                           => n8879);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT1(7), QN 
                           => n8880);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => OUT1(6), QN 
                           => n8881);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT1(5), QN 
                           => n8882);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => OUT1(4), QN 
                           => n8883);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT1(3), QN 
                           => n8884);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => OUT1(2), QN 
                           => n8885);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT1(1), QN 
                           => n8886);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => OUT1(0), QN 
                           => n8887);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT2(31), QN
                           => n8888);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT2(30), QN
                           => n8905);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT2(29), QN
                           => n8922);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT2(28), QN
                           => n8939);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT2(27), QN
                           => n8956);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT2(26), QN
                           => n8973);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT2(25), QN
                           => n8990);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT2(24), QN
                           => n9007);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT2(23), QN
                           => n9024);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT2(22), QN
                           => n9041);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT2(21), QN
                           => n9058);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT2(20), QN
                           => n9075);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT2(19), QN
                           => n9092);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT2(18), QN
                           => n9109);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT2(17), QN
                           => n9126);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT2(16), QN
                           => n9143);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT2(15), QN
                           => n9160);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT2(14), QN
                           => n9177);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT2(13), QN
                           => n9194);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => OUT2(12), QN
                           => n9211);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT2(11), QN
                           => n9228);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT2(10), QN
                           => n9245);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT2(9), QN 
                           => n9262);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT2(8), QN 
                           => n9279);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT2(7), QN 
                           => n9296);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT2(6), QN 
                           => n9313);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT2(5), QN 
                           => n9330);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT2(4), QN 
                           => n9347);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT2(3), QN 
                           => n9364);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT2(2), QN 
                           => n9381);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT2(1), QN 
                           => n9398);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT2(0), QN 
                           => n9415);
   REGS_reg_17_31_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => n_1000, 
                           QN => n16652);
   REGS_reg_17_30_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => n_1001, 
                           QN => n16651);
   REGS_reg_17_29_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => n_1002, 
                           QN => n16650);
   REGS_reg_17_28_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => n_1003, 
                           QN => n16649);
   REGS_reg_17_27_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => n_1004, 
                           QN => n16648);
   REGS_reg_17_26_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => n_1005, 
                           QN => n16647);
   REGS_reg_17_25_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => n_1006, 
                           QN => n16646);
   REGS_reg_17_24_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => n_1007, 
                           QN => n16645);
   REGS_reg_16_30_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => n_1008, 
                           QN => n16811);
   REGS_reg_16_29_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => n_1009, 
                           QN => n16810);
   REGS_reg_16_28_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => n_1010, 
                           QN => n16809);
   REGS_reg_16_27_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => n_1011, 
                           QN => n16808);
   REGS_reg_16_26_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => n_1012, 
                           QN => n16807);
   REGS_reg_16_25_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => n_1013, 
                           QN => n16806);
   REGS_reg_16_24_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => n_1014, 
                           QN => n16805);
   REGS_reg_17_23_inst : DFF_X1 port map( D => n3064, CK => CLK, Q => n_1015, 
                           QN => n16644);
   REGS_reg_17_22_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => n_1016, 
                           QN => n16643);
   REGS_reg_17_21_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => n_1017, 
                           QN => n16642);
   REGS_reg_17_20_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => n_1018, 
                           QN => n16641);
   REGS_reg_17_19_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => n_1019, 
                           QN => n16640);
   REGS_reg_17_18_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => n_1020, 
                           QN => n16639);
   REGS_reg_17_17_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => n_1021, 
                           QN => n16638);
   REGS_reg_17_16_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => n_1022, 
                           QN => n16637);
   REGS_reg_17_15_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => n_1023, 
                           QN => n16636);
   REGS_reg_17_14_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => n_1024, 
                           QN => n16635);
   REGS_reg_17_13_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => n_1025, 
                           QN => n16634);
   REGS_reg_17_12_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => n_1026, 
                           QN => n16633);
   REGS_reg_17_11_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => n_1027, 
                           QN => n16748);
   REGS_reg_17_10_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => n_1028, 
                           QN => n16747);
   REGS_reg_17_9_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => n_1029, QN
                           => n16746);
   REGS_reg_17_8_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => n_1030, QN
                           => n16745);
   REGS_reg_17_7_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => n_1031, QN
                           => n16744);
   REGS_reg_17_6_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => n_1032, QN
                           => n16743);
   REGS_reg_17_5_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => n_1033, QN
                           => n16742);
   REGS_reg_17_4_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => n_1034, QN
                           => n16741);
   REGS_reg_17_3_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => n_1035, QN
                           => n16740);
   REGS_reg_17_2_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => n_1036, QN
                           => n16739);
   REGS_reg_17_1_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => n_1037, QN
                           => n16738);
   REGS_reg_17_0_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => n_1038, QN
                           => n16737);
   REGS_reg_16_23_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => n_1039, 
                           QN => n17244);
   REGS_reg_16_22_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => n_1040, 
                           QN => n17243);
   REGS_reg_16_21_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => n_1041, 
                           QN => n17242);
   REGS_reg_16_20_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => n_1042, 
                           QN => n17241);
   REGS_reg_16_19_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => n_1043, 
                           QN => n17240);
   REGS_reg_16_18_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => n_1044, 
                           QN => n17239);
   REGS_reg_16_17_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => n_1045, 
                           QN => n17238);
   REGS_reg_16_16_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => n_1046, 
                           QN => n17237);
   REGS_reg_16_15_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => n_1047, 
                           QN => n17236);
   REGS_reg_16_14_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => n_1048, 
                           QN => n17235);
   REGS_reg_16_13_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => n_1049, 
                           QN => n17234);
   REGS_reg_16_12_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => n_1050, 
                           QN => n17233);
   REGS_reg_16_11_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => n_1051, 
                           QN => n17232);
   REGS_reg_16_10_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => n_1052, 
                           QN => n17231);
   REGS_reg_16_9_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => n_1053, QN
                           => n17230);
   REGS_reg_16_8_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => n_1054, QN
                           => n17229);
   REGS_reg_16_7_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => n_1055, QN
                           => n17228);
   REGS_reg_16_6_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => n_1056, QN
                           => n17227);
   REGS_reg_16_5_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => n_1057, QN
                           => n17226);
   REGS_reg_16_4_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => n_1058, QN
                           => n17225);
   REGS_reg_16_3_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => n_1059, QN
                           => n17224);
   REGS_reg_16_2_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => n_1060, QN
                           => n17223);
   REGS_reg_16_1_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => n_1061, QN
                           => n17222);
   REGS_reg_16_0_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => n_1062, QN
                           => n17221);
   REGS_reg_31_31_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => n17276, 
                           QN => n8903);
   REGS_reg_31_30_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => n17275, 
                           QN => n8920);
   REGS_reg_31_29_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => n17274, 
                           QN => n8937);
   REGS_reg_31_28_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => n17273, 
                           QN => n8954);
   REGS_reg_31_27_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => n17272, 
                           QN => n8971);
   REGS_reg_31_26_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => n17271, 
                           QN => n8988);
   REGS_reg_31_25_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => n17270, 
                           QN => n9005);
   REGS_reg_31_24_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => n17269, 
                           QN => n9022);
   REGS_reg_31_23_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => n17268, 
                           QN => n9039);
   REGS_reg_31_22_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => n17267, 
                           QN => n9056);
   REGS_reg_31_21_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => n17266, 
                           QN => n9073);
   REGS_reg_31_20_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => n17265, 
                           QN => n9090);
   REGS_reg_31_19_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => n17264, 
                           QN => n9107);
   REGS_reg_31_18_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => n17263, 
                           QN => n9124);
   REGS_reg_31_17_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => n17262, 
                           QN => n9141);
   REGS_reg_31_16_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => n17261, 
                           QN => n9158);
   REGS_reg_31_15_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => n17260, 
                           QN => n9175);
   REGS_reg_31_14_inst : DFF_X1 port map( D => n2607, CK => CLK, Q => n17259, 
                           QN => n9192);
   REGS_reg_31_13_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => n17258, 
                           QN => n9209);
   REGS_reg_31_12_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => n17257, 
                           QN => n9226);
   REGS_reg_31_11_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => n17256, 
                           QN => n9243);
   REGS_reg_31_10_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => n17255, 
                           QN => n9260);
   REGS_reg_31_9_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => n17254, QN
                           => n9277);
   REGS_reg_31_8_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => n17253, QN
                           => n9294);
   REGS_reg_31_7_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => n17252, QN
                           => n9311);
   REGS_reg_31_6_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => n17251, QN
                           => n9328);
   REGS_reg_31_5_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => n17250, QN
                           => n9345);
   REGS_reg_31_4_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => n17249, QN
                           => n9362);
   REGS_reg_31_3_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => n17248, QN
                           => n9379);
   REGS_reg_31_2_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => n17247, QN
                           => n9396);
   REGS_reg_31_1_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => n17246, QN
                           => n9413);
   REGS_reg_31_0_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => n17245, QN
                           => n9430);
   REGS_reg_30_31_inst : DFF_X1 port map( D => n2656, CK => CLK, Q => n17027, 
                           QN => n8904);
   REGS_reg_30_30_inst : DFF_X1 port map( D => n2655, CK => CLK, Q => n17025, 
                           QN => n8921);
   REGS_reg_30_29_inst : DFF_X1 port map( D => n2654, CK => CLK, Q => n17023, 
                           QN => n8938);
   REGS_reg_30_28_inst : DFF_X1 port map( D => n2653, CK => CLK, Q => n17021, 
                           QN => n8955);
   REGS_reg_30_27_inst : DFF_X1 port map( D => n2652, CK => CLK, Q => n17019, 
                           QN => n8972);
   REGS_reg_30_26_inst : DFF_X1 port map( D => n2651, CK => CLK, Q => n17017, 
                           QN => n8989);
   REGS_reg_30_25_inst : DFF_X1 port map( D => n2650, CK => CLK, Q => n17015, 
                           QN => n9006);
   REGS_reg_30_24_inst : DFF_X1 port map( D => n2649, CK => CLK, Q => n17013, 
                           QN => n9023);
   REGS_reg_27_31_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => n17427, 
                           QN => n8901);
   REGS_reg_27_30_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => n17425, 
                           QN => n8918);
   REGS_reg_27_29_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => n17423, 
                           QN => n8935);
   REGS_reg_27_28_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => n17421, 
                           QN => n8952);
   REGS_reg_27_27_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => n17419, 
                           QN => n8969);
   REGS_reg_27_26_inst : DFF_X1 port map( D => n2747, CK => CLK, Q => n17417, 
                           QN => n8986);
   REGS_reg_27_25_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => n17415, 
                           QN => n9003);
   REGS_reg_27_24_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => n17413, 
                           QN => n9020);
   REGS_reg_26_31_inst : DFF_X1 port map( D => n2784, CK => CLK, Q => n16963, 
                           QN => n8902);
   REGS_reg_26_30_inst : DFF_X1 port map( D => n2783, CK => CLK, Q => n16961, 
                           QN => n8919);
   REGS_reg_26_29_inst : DFF_X1 port map( D => n2782, CK => CLK, Q => n16959, 
                           QN => n8936);
   REGS_reg_26_28_inst : DFF_X1 port map( D => n2781, CK => CLK, Q => n16957, 
                           QN => n8953);
   REGS_reg_26_27_inst : DFF_X1 port map( D => n2780, CK => CLK, Q => n16955, 
                           QN => n8970);
   REGS_reg_26_26_inst : DFF_X1 port map( D => n2779, CK => CLK, Q => n16953, 
                           QN => n8987);
   REGS_reg_26_25_inst : DFF_X1 port map( D => n2778, CK => CLK, Q => n16951, 
                           QN => n9004);
   REGS_reg_26_24_inst : DFF_X1 port map( D => n2777, CK => CLK, Q => n16949, 
                           QN => n9021);
   REGS_reg_21_31_inst : DFF_X1 port map( D => n2944, CK => CLK, Q => n17468, 
                           QN => n8899);
   REGS_reg_21_30_inst : DFF_X1 port map( D => n2943, CK => CLK, Q => n17467, 
                           QN => n8916);
   REGS_reg_21_29_inst : DFF_X1 port map( D => n2942, CK => CLK, Q => n17466, 
                           QN => n8933);
   REGS_reg_21_28_inst : DFF_X1 port map( D => n2941, CK => CLK, Q => n17465, 
                           QN => n8950);
   REGS_reg_21_27_inst : DFF_X1 port map( D => n2940, CK => CLK, Q => n17464, 
                           QN => n8967);
   REGS_reg_21_26_inst : DFF_X1 port map( D => n2939, CK => CLK, Q => n17463, 
                           QN => n8984);
   REGS_reg_21_25_inst : DFF_X1 port map( D => n2938, CK => CLK, Q => n17462, 
                           QN => n9001);
   REGS_reg_21_24_inst : DFF_X1 port map( D => n2937, CK => CLK, Q => n17461, 
                           QN => n9018);
   REGS_reg_20_31_inst : DFF_X1 port map( D => n2976, CK => CLK, Q => n17036, 
                           QN => n8900);
   REGS_reg_20_30_inst : DFF_X1 port map( D => n2975, CK => CLK, Q => n17035, 
                           QN => n8917);
   REGS_reg_20_29_inst : DFF_X1 port map( D => n2974, CK => CLK, Q => n17034, 
                           QN => n8934);
   REGS_reg_20_28_inst : DFF_X1 port map( D => n2973, CK => CLK, Q => n17033, 
                           QN => n8951);
   REGS_reg_20_27_inst : DFF_X1 port map( D => n2972, CK => CLK, Q => n17032, 
                           QN => n8968);
   REGS_reg_20_26_inst : DFF_X1 port map( D => n2971, CK => CLK, Q => n17031, 
                           QN => n8985);
   REGS_reg_20_25_inst : DFF_X1 port map( D => n2970, CK => CLK, Q => n17030, 
                           QN => n9002);
   REGS_reg_20_24_inst : DFF_X1 port map( D => n2969, CK => CLK, Q => n17029, 
                           QN => n9019);
   REGS_reg_13_31_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => n17460, 
                           QN => n8895);
   REGS_reg_13_30_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => n17459, 
                           QN => n8912);
   REGS_reg_13_29_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => n17458, 
                           QN => n8929);
   REGS_reg_13_28_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => n17457, 
                           QN => n8946);
   REGS_reg_13_27_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => n17456, 
                           QN => n8963);
   REGS_reg_13_26_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => n17455, 
                           QN => n8980);
   REGS_reg_13_25_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => n17454, 
                           QN => n8997);
   REGS_reg_13_24_inst : DFF_X1 port map( D => n3193, CK => CLK, Q => n17453, 
                           QN => n9014);
   REGS_reg_12_31_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => n17028, 
                           QN => n8896);
   REGS_reg_12_30_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => n17026, 
                           QN => n8913);
   REGS_reg_12_29_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => n17024, 
                           QN => n8930);
   REGS_reg_12_28_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => n17022, 
                           QN => n8947);
   REGS_reg_12_27_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => n17020, 
                           QN => n8964);
   REGS_reg_12_26_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => n17018, 
                           QN => n8981);
   REGS_reg_12_25_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => n17016, 
                           QN => n8998);
   REGS_reg_12_24_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => n17014, 
                           QN => n9015);
   REGS_reg_9_31_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => n17428, QN
                           => n8893);
   REGS_reg_9_30_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => n17426, QN
                           => n8910);
   REGS_reg_9_29_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => n17424, QN
                           => n8927);
   REGS_reg_9_28_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => n17422, QN
                           => n8944);
   REGS_reg_9_27_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => n17420, QN
                           => n8961);
   REGS_reg_9_26_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => n17418, QN
                           => n8978);
   REGS_reg_9_25_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => n17416, QN
                           => n8995);
   REGS_reg_9_24_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => n17414, QN
                           => n9012);
   REGS_reg_8_31_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => n16964, QN
                           => n8894);
   REGS_reg_8_30_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => n16962, QN
                           => n8911);
   REGS_reg_8_29_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => n16960, QN
                           => n8928);
   REGS_reg_8_28_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => n16958, QN
                           => n8945);
   REGS_reg_8_27_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => n16956, QN
                           => n8962);
   REGS_reg_8_26_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => n16954, QN
                           => n8979);
   REGS_reg_8_25_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => n16952, QN
                           => n8996);
   REGS_reg_8_24_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => n16950, QN
                           => n9013);
   REGS_reg_5_31_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => n17364, QN
                           => n6672);
   REGS_reg_5_30_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => n17363, QN
                           => n6673);
   REGS_reg_5_29_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => n17362, QN
                           => n6674);
   REGS_reg_5_28_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => n17361, QN
                           => n6675);
   REGS_reg_5_27_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => n17360, QN
                           => n6676);
   REGS_reg_5_26_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => n17359, QN
                           => n6677);
   REGS_reg_5_25_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => n17358, QN
                           => n6678);
   REGS_reg_5_24_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => n17357, QN
                           => n6679);
   REGS_reg_4_31_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => n16900, QN
                           => n6640);
   REGS_reg_4_30_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => n16899, QN
                           => n6641);
   REGS_reg_4_29_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => n16898, QN
                           => n6642);
   REGS_reg_4_28_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => n16897, QN
                           => n6643);
   REGS_reg_4_27_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => n16896, QN
                           => n6644);
   REGS_reg_4_26_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => n16895, QN
                           => n6645);
   REGS_reg_4_25_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => n16894, QN
                           => n6646);
   REGS_reg_4_24_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => n16893, QN
                           => n6647);
   REGS_reg_3_31_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => n16844, QN
                           => n8890);
   REGS_reg_3_30_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => n16843, QN
                           => n8907);
   REGS_reg_3_29_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => n16842, QN
                           => n8924);
   REGS_reg_3_28_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => n16841, QN
                           => n8941);
   REGS_reg_3_27_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => n16840, QN
                           => n8958);
   REGS_reg_3_26_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => n16839, QN
                           => n8975);
   REGS_reg_3_25_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => n16838, QN
                           => n8992);
   REGS_reg_3_24_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => n16837, QN
                           => n9009);
   REGS_reg_2_31_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => n17308, QN
                           => n8889);
   REGS_reg_2_30_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => n17307, QN
                           => n8906);
   REGS_reg_2_29_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => n17306, QN
                           => n8923);
   REGS_reg_2_28_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => n17305, QN
                           => n8940);
   REGS_reg_2_27_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => n17304, QN
                           => n8957);
   REGS_reg_2_26_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => n17303, QN
                           => n8974);
   REGS_reg_2_25_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => n17302, QN
                           => n8991);
   REGS_reg_2_24_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => n17301, QN
                           => n9008);
   REGS_reg_30_23_inst : DFF_X1 port map( D => n2648, CK => CLK, Q => n17011, 
                           QN => n9040);
   REGS_reg_30_22_inst : DFF_X1 port map( D => n2647, CK => CLK, Q => n17009, 
                           QN => n9057);
   REGS_reg_30_21_inst : DFF_X1 port map( D => n2646, CK => CLK, Q => n17007, 
                           QN => n9074);
   REGS_reg_30_20_inst : DFF_X1 port map( D => n2645, CK => CLK, Q => n17005, 
                           QN => n9091);
   REGS_reg_30_19_inst : DFF_X1 port map( D => n2644, CK => CLK, Q => n17003, 
                           QN => n9108);
   REGS_reg_30_18_inst : DFF_X1 port map( D => n2643, CK => CLK, Q => n17001, 
                           QN => n9125);
   REGS_reg_30_17_inst : DFF_X1 port map( D => n2642, CK => CLK, Q => n16999, 
                           QN => n9142);
   REGS_reg_30_16_inst : DFF_X1 port map( D => n2641, CK => CLK, Q => n16997, 
                           QN => n9159);
   REGS_reg_30_15_inst : DFF_X1 port map( D => n2640, CK => CLK, Q => n16995, 
                           QN => n9176);
   REGS_reg_30_14_inst : DFF_X1 port map( D => n2639, CK => CLK, Q => n16993, 
                           QN => n9193);
   REGS_reg_30_13_inst : DFF_X1 port map( D => n2638, CK => CLK, Q => n16991, 
                           QN => n9210);
   REGS_reg_30_12_inst : DFF_X1 port map( D => n2637, CK => CLK, Q => n16989, 
                           QN => n9227);
   REGS_reg_30_11_inst : DFF_X1 port map( D => n2636, CK => CLK, Q => n16987, 
                           QN => n9244);
   REGS_reg_30_10_inst : DFF_X1 port map( D => n2635, CK => CLK, Q => n16985, 
                           QN => n9261);
   REGS_reg_30_9_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => n16983, QN
                           => n9278);
   REGS_reg_30_8_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => n16981, QN
                           => n9295);
   REGS_reg_30_7_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => n16979, QN
                           => n9312);
   REGS_reg_30_6_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => n16977, QN
                           => n9329);
   REGS_reg_30_5_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => n16975, QN
                           => n9346);
   REGS_reg_30_4_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => n16973, QN
                           => n9363);
   REGS_reg_30_3_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => n16971, QN
                           => n9380);
   REGS_reg_30_2_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => n16969, QN
                           => n9397);
   REGS_reg_30_1_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => n16967, QN
                           => n9414);
   REGS_reg_30_0_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => n16965, QN
                           => n9431);
   REGS_reg_27_23_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => n17411, 
                           QN => n9037);
   REGS_reg_27_22_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => n17409, 
                           QN => n9054);
   REGS_reg_27_21_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => n17407, 
                           QN => n9071);
   REGS_reg_27_20_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => n17405, 
                           QN => n9088);
   REGS_reg_27_19_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => n17403, 
                           QN => n9105);
   REGS_reg_27_18_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => n17401, 
                           QN => n9122);
   REGS_reg_27_17_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => n17399, 
                           QN => n9139);
   REGS_reg_27_16_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => n17397, 
                           QN => n9156);
   REGS_reg_27_15_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => n17395, 
                           QN => n9173);
   REGS_reg_27_14_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => n17393, 
                           QN => n9190);
   REGS_reg_27_13_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => n17391, 
                           QN => n9207);
   REGS_reg_27_12_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => n17389, 
                           QN => n9224);
   REGS_reg_27_11_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => n17387, 
                           QN => n9241);
   REGS_reg_27_10_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => n17385, 
                           QN => n9258);
   REGS_reg_27_9_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => n17383, QN
                           => n9275);
   REGS_reg_27_8_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => n17381, QN
                           => n9292);
   REGS_reg_27_7_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => n17379, QN
                           => n9309);
   REGS_reg_27_6_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => n17377, QN
                           => n9326);
   REGS_reg_27_5_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => n17375, QN
                           => n9343);
   REGS_reg_27_4_inst : DFF_X1 port map( D => n2725, CK => CLK, Q => n17373, QN
                           => n9360);
   REGS_reg_27_3_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => n17371, QN
                           => n9377);
   REGS_reg_27_2_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => n17369, QN
                           => n9394);
   REGS_reg_27_1_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => n17367, QN
                           => n9411);
   REGS_reg_27_0_inst : DFF_X1 port map( D => n2721, CK => CLK, Q => n17365, QN
                           => n9428);
   REGS_reg_26_23_inst : DFF_X1 port map( D => n2776, CK => CLK, Q => n16947, 
                           QN => n9038);
   REGS_reg_26_22_inst : DFF_X1 port map( D => n2775, CK => CLK, Q => n16945, 
                           QN => n9055);
   REGS_reg_26_21_inst : DFF_X1 port map( D => n2774, CK => CLK, Q => n16943, 
                           QN => n9072);
   REGS_reg_26_20_inst : DFF_X1 port map( D => n2773, CK => CLK, Q => n16941, 
                           QN => n9089);
   REGS_reg_26_19_inst : DFF_X1 port map( D => n2772, CK => CLK, Q => n16939, 
                           QN => n9106);
   REGS_reg_26_18_inst : DFF_X1 port map( D => n2771, CK => CLK, Q => n16937, 
                           QN => n9123);
   REGS_reg_26_17_inst : DFF_X1 port map( D => n2770, CK => CLK, Q => n16935, 
                           QN => n9140);
   REGS_reg_26_16_inst : DFF_X1 port map( D => n2769, CK => CLK, Q => n16933, 
                           QN => n9157);
   REGS_reg_26_15_inst : DFF_X1 port map( D => n2768, CK => CLK, Q => n16931, 
                           QN => n9174);
   REGS_reg_26_14_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => n16929, 
                           QN => n9191);
   REGS_reg_26_13_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => n16927, 
                           QN => n9208);
   REGS_reg_26_12_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => n16925, 
                           QN => n9225);
   REGS_reg_26_11_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => n16923, 
                           QN => n9242);
   REGS_reg_26_10_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => n16921, 
                           QN => n9259);
   REGS_reg_26_9_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => n16919, QN
                           => n9276);
   REGS_reg_26_8_inst : DFF_X1 port map( D => n2761, CK => CLK, Q => n16917, QN
                           => n9293);
   REGS_reg_26_7_inst : DFF_X1 port map( D => n2760, CK => CLK, Q => n16915, QN
                           => n9310);
   REGS_reg_26_6_inst : DFF_X1 port map( D => n2759, CK => CLK, Q => n16913, QN
                           => n9327);
   REGS_reg_26_5_inst : DFF_X1 port map( D => n2758, CK => CLK, Q => n16911, QN
                           => n9344);
   REGS_reg_26_4_inst : DFF_X1 port map( D => n2757, CK => CLK, Q => n16909, QN
                           => n9361);
   REGS_reg_26_3_inst : DFF_X1 port map( D => n2756, CK => CLK, Q => n16907, QN
                           => n9378);
   REGS_reg_26_2_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => n16905, QN
                           => n9395);
   REGS_reg_26_1_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => n16903, QN
                           => n9412);
   REGS_reg_26_0_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => n16901, QN
                           => n9429);
   REGS_reg_21_23_inst : DFF_X1 port map( D => n2936, CK => CLK, Q => n17355, 
                           QN => n9035);
   REGS_reg_21_22_inst : DFF_X1 port map( D => n2935, CK => CLK, Q => n17353, 
                           QN => n9052);
   REGS_reg_21_21_inst : DFF_X1 port map( D => n2934, CK => CLK, Q => n17351, 
                           QN => n9069);
   REGS_reg_21_20_inst : DFF_X1 port map( D => n2933, CK => CLK, Q => n17349, 
                           QN => n9086);
   REGS_reg_21_19_inst : DFF_X1 port map( D => n2932, CK => CLK, Q => n17347, 
                           QN => n9103);
   REGS_reg_21_18_inst : DFF_X1 port map( D => n2931, CK => CLK, Q => n17345, 
                           QN => n9120);
   REGS_reg_21_17_inst : DFF_X1 port map( D => n2930, CK => CLK, Q => n17343, 
                           QN => n9137);
   REGS_reg_21_16_inst : DFF_X1 port map( D => n2929, CK => CLK, Q => n17341, 
                           QN => n9154);
   REGS_reg_21_15_inst : DFF_X1 port map( D => n2928, CK => CLK, Q => n17339, 
                           QN => n9171);
   REGS_reg_21_14_inst : DFF_X1 port map( D => n2927, CK => CLK, Q => n17337, 
                           QN => n9188);
   REGS_reg_21_13_inst : DFF_X1 port map( D => n2926, CK => CLK, Q => n17335, 
                           QN => n9205);
   REGS_reg_21_12_inst : DFF_X1 port map( D => n2925, CK => CLK, Q => n17333, 
                           QN => n9222);
   REGS_reg_21_11_inst : DFF_X1 port map( D => n2924, CK => CLK, Q => n17331, 
                           QN => n9239);
   REGS_reg_21_10_inst : DFF_X1 port map( D => n2923, CK => CLK, Q => n17329, 
                           QN => n9256);
   REGS_reg_21_9_inst : DFF_X1 port map( D => n2922, CK => CLK, Q => n17327, QN
                           => n9273);
   REGS_reg_21_8_inst : DFF_X1 port map( D => n2921, CK => CLK, Q => n17325, QN
                           => n9290);
   REGS_reg_21_7_inst : DFF_X1 port map( D => n2920, CK => CLK, Q => n17323, QN
                           => n9307);
   REGS_reg_21_6_inst : DFF_X1 port map( D => n2919, CK => CLK, Q => n17321, QN
                           => n9324);
   REGS_reg_21_5_inst : DFF_X1 port map( D => n2918, CK => CLK, Q => n17319, QN
                           => n9341);
   REGS_reg_21_4_inst : DFF_X1 port map( D => n2917, CK => CLK, Q => n17317, QN
                           => n9358);
   REGS_reg_21_3_inst : DFF_X1 port map( D => n2916, CK => CLK, Q => n17315, QN
                           => n9375);
   REGS_reg_21_2_inst : DFF_X1 port map( D => n2915, CK => CLK, Q => n17313, QN
                           => n9392);
   REGS_reg_21_1_inst : DFF_X1 port map( D => n2914, CK => CLK, Q => n17311, QN
                           => n9409);
   REGS_reg_21_0_inst : DFF_X1 port map( D => n2913, CK => CLK, Q => n17309, QN
                           => n9426);
   REGS_reg_20_23_inst : DFF_X1 port map( D => n2968, CK => CLK, Q => n16891, 
                           QN => n9036);
   REGS_reg_20_22_inst : DFF_X1 port map( D => n2967, CK => CLK, Q => n16889, 
                           QN => n9053);
   REGS_reg_20_21_inst : DFF_X1 port map( D => n2966, CK => CLK, Q => n16887, 
                           QN => n9070);
   REGS_reg_20_20_inst : DFF_X1 port map( D => n2965, CK => CLK, Q => n16885, 
                           QN => n9087);
   REGS_reg_20_19_inst : DFF_X1 port map( D => n2964, CK => CLK, Q => n16883, 
                           QN => n9104);
   REGS_reg_20_18_inst : DFF_X1 port map( D => n2963, CK => CLK, Q => n16881, 
                           QN => n9121);
   REGS_reg_20_17_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => n16879, 
                           QN => n9138);
   REGS_reg_20_16_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => n16877, 
                           QN => n9155);
   REGS_reg_20_15_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => n16875, 
                           QN => n9172);
   REGS_reg_20_14_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => n16873, 
                           QN => n9189);
   REGS_reg_20_13_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => n16871, 
                           QN => n9206);
   REGS_reg_20_12_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => n16869, 
                           QN => n9223);
   REGS_reg_20_11_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => n16867, 
                           QN => n9240);
   REGS_reg_20_10_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => n16865, 
                           QN => n9257);
   REGS_reg_20_9_inst : DFF_X1 port map( D => n2954, CK => CLK, Q => n16863, QN
                           => n9274);
   REGS_reg_20_8_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => n16861, QN
                           => n9291);
   REGS_reg_20_7_inst : DFF_X1 port map( D => n2952, CK => CLK, Q => n16859, QN
                           => n9308);
   REGS_reg_20_6_inst : DFF_X1 port map( D => n2951, CK => CLK, Q => n16857, QN
                           => n9325);
   REGS_reg_20_5_inst : DFF_X1 port map( D => n2950, CK => CLK, Q => n16855, QN
                           => n9342);
   REGS_reg_20_4_inst : DFF_X1 port map( D => n2949, CK => CLK, Q => n16853, QN
                           => n9359);
   REGS_reg_20_3_inst : DFF_X1 port map( D => n2948, CK => CLK, Q => n16851, QN
                           => n9376);
   REGS_reg_20_2_inst : DFF_X1 port map( D => n2947, CK => CLK, Q => n16849, QN
                           => n9393);
   REGS_reg_20_1_inst : DFF_X1 port map( D => n2946, CK => CLK, Q => n16847, QN
                           => n9410);
   REGS_reg_20_0_inst : DFF_X1 port map( D => n2945, CK => CLK, Q => n16845, QN
                           => n9427);
   REGS_reg_13_23_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => n17452, 
                           QN => n9031);
   REGS_reg_13_22_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => n17451, 
                           QN => n9048);
   REGS_reg_13_21_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => n17450, 
                           QN => n9065);
   REGS_reg_13_20_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => n17449, 
                           QN => n9082);
   REGS_reg_13_19_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => n17448, 
                           QN => n9099);
   REGS_reg_13_18_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => n17447, 
                           QN => n9116);
   REGS_reg_13_17_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => n17446, 
                           QN => n9133);
   REGS_reg_13_16_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => n17445, 
                           QN => n9150);
   REGS_reg_13_15_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => n17444, 
                           QN => n9167);
   REGS_reg_13_14_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => n17443, 
                           QN => n9184);
   REGS_reg_13_13_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => n17442, 
                           QN => n9201);
   REGS_reg_13_12_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => n17441, 
                           QN => n9218);
   REGS_reg_13_11_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => n17440, 
                           QN => n9235);
   REGS_reg_13_10_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => n17439, 
                           QN => n9252);
   REGS_reg_13_9_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => n17438, QN
                           => n9269);
   REGS_reg_13_8_inst : DFF_X1 port map( D => n3177, CK => CLK, Q => n17437, QN
                           => n9286);
   REGS_reg_13_7_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => n17436, QN
                           => n9303);
   REGS_reg_13_6_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => n17435, QN
                           => n9320);
   REGS_reg_13_5_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => n17434, QN
                           => n9337);
   REGS_reg_13_4_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => n17433, QN
                           => n9354);
   REGS_reg_13_3_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => n17432, QN
                           => n9371);
   REGS_reg_13_2_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => n17431, QN
                           => n9388);
   REGS_reg_13_1_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => n17430, QN
                           => n9405);
   REGS_reg_13_0_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => n17429, QN
                           => n9422);
   REGS_reg_12_23_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => n17012, 
                           QN => n9032);
   REGS_reg_12_22_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => n17010, 
                           QN => n9049);
   REGS_reg_12_21_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => n17008, 
                           QN => n9066);
   REGS_reg_12_20_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => n17006, 
                           QN => n9083);
   REGS_reg_12_19_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => n17004, 
                           QN => n9100);
   REGS_reg_12_18_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => n17002, 
                           QN => n9117);
   REGS_reg_12_17_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => n17000, 
                           QN => n9134);
   REGS_reg_12_16_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => n16998, 
                           QN => n9151);
   REGS_reg_12_15_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => n16996, 
                           QN => n9168);
   REGS_reg_12_14_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => n16994, 
                           QN => n9185);
   REGS_reg_12_13_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => n16992, 
                           QN => n9202);
   REGS_reg_12_12_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => n16990, 
                           QN => n9219);
   REGS_reg_12_11_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => n16988, 
                           QN => n9236);
   REGS_reg_12_10_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => n16986, 
                           QN => n9253);
   REGS_reg_12_9_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => n16984, QN
                           => n9270);
   REGS_reg_12_8_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => n16982, QN
                           => n9287);
   REGS_reg_12_7_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => n16980, QN
                           => n9304);
   REGS_reg_12_6_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => n16978, QN
                           => n9321);
   REGS_reg_12_5_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => n16976, QN
                           => n9338);
   REGS_reg_12_4_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => n16974, QN
                           => n9355);
   REGS_reg_12_3_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => n16972, QN
                           => n9372);
   REGS_reg_12_2_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => n16970, QN
                           => n9389);
   REGS_reg_12_1_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => n16968, QN
                           => n9406);
   REGS_reg_12_0_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => n16966, QN
                           => n9423);
   REGS_reg_9_23_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => n17412, QN
                           => n9029);
   REGS_reg_9_22_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => n17410, QN
                           => n9046);
   REGS_reg_9_21_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => n17408, QN
                           => n9063);
   REGS_reg_9_20_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => n17406, QN
                           => n9080);
   REGS_reg_9_19_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => n17404, QN
                           => n9097);
   REGS_reg_9_18_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => n17402, QN
                           => n9114);
   REGS_reg_9_17_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => n17400, QN
                           => n9131);
   REGS_reg_9_16_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => n17398, QN
                           => n9148);
   REGS_reg_9_15_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => n17396, QN
                           => n9165);
   REGS_reg_9_14_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => n17394, QN
                           => n9182);
   REGS_reg_9_13_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => n17392, QN
                           => n9199);
   REGS_reg_9_12_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => n17390, QN
                           => n9216);
   REGS_reg_9_11_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => n17388, QN
                           => n9233);
   REGS_reg_9_10_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => n17386, QN
                           => n9250);
   REGS_reg_9_9_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => n17384, QN 
                           => n9267);
   REGS_reg_9_8_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => n17382, QN 
                           => n9284);
   REGS_reg_9_7_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => n17380, QN 
                           => n9301);
   REGS_reg_9_6_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => n17378, QN 
                           => n9318);
   REGS_reg_9_5_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => n17376, QN 
                           => n9335);
   REGS_reg_9_4_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => n17374, QN 
                           => n9352);
   REGS_reg_9_3_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => n17372, QN 
                           => n9369);
   REGS_reg_9_2_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => n17370, QN 
                           => n9386);
   REGS_reg_9_1_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => n17368, QN 
                           => n9403);
   REGS_reg_9_0_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => n17366, QN 
                           => n9420);
   REGS_reg_8_23_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => n16948, QN
                           => n9030);
   REGS_reg_8_22_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => n16946, QN
                           => n9047);
   REGS_reg_8_21_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => n16944, QN
                           => n9064);
   REGS_reg_8_20_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => n16942, QN
                           => n9081);
   REGS_reg_8_19_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => n16940, QN
                           => n9098);
   REGS_reg_8_18_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => n16938, QN
                           => n9115);
   REGS_reg_8_17_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => n16936, QN
                           => n9132);
   REGS_reg_8_16_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => n16934, QN
                           => n9149);
   REGS_reg_8_15_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => n16932, QN
                           => n9166);
   REGS_reg_8_14_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => n16930, QN
                           => n9183);
   REGS_reg_8_13_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => n16928, QN
                           => n9200);
   REGS_reg_8_12_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => n16926, QN
                           => n9217);
   REGS_reg_8_11_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => n16924, QN
                           => n9234);
   REGS_reg_8_10_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => n16922, QN
                           => n9251);
   REGS_reg_8_9_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => n16920, QN 
                           => n9268);
   REGS_reg_8_8_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => n16918, QN 
                           => n9285);
   REGS_reg_8_7_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => n16916, QN 
                           => n9302);
   REGS_reg_8_6_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => n16914, QN 
                           => n9319);
   REGS_reg_8_5_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => n16912, QN 
                           => n9336);
   REGS_reg_8_4_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => n16910, QN 
                           => n9353);
   REGS_reg_8_3_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => n16908, QN 
                           => n9370);
   REGS_reg_8_2_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => n16906, QN 
                           => n9387);
   REGS_reg_8_1_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => n16904, QN 
                           => n9404);
   REGS_reg_8_0_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => n16902, QN 
                           => n9421);
   REGS_reg_5_23_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => n17356, QN
                           => n6680);
   REGS_reg_5_22_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => n17354, QN
                           => n6681);
   REGS_reg_5_21_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => n17352, QN
                           => n6682);
   REGS_reg_5_20_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => n17350, QN
                           => n6683);
   REGS_reg_5_19_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => n17348, QN
                           => n6684);
   REGS_reg_5_18_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => n17346, QN
                           => n6685);
   REGS_reg_5_17_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => n17344, QN
                           => n6686);
   REGS_reg_5_16_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => n17342, QN
                           => n6687);
   REGS_reg_5_15_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => n17340, QN
                           => n6688);
   REGS_reg_5_14_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => n17338, QN
                           => n6689);
   REGS_reg_5_13_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => n17336, QN
                           => n6690);
   REGS_reg_5_12_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => n17334, QN
                           => n6691);
   REGS_reg_5_11_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => n17332, QN
                           => n6692);
   REGS_reg_5_10_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => n17330, QN
                           => n6693);
   REGS_reg_5_9_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => n17328, QN 
                           => n6694);
   REGS_reg_5_8_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => n17326, QN 
                           => n6695);
   REGS_reg_5_7_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => n17324, QN 
                           => n6696);
   REGS_reg_5_6_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => n17322, QN 
                           => n6697);
   REGS_reg_5_5_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => n17320, QN 
                           => n6698);
   REGS_reg_5_4_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => n17318, QN 
                           => n6699);
   REGS_reg_5_3_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => n17316, QN 
                           => n6700);
   REGS_reg_5_2_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => n17314, QN 
                           => n6701);
   REGS_reg_5_1_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => n17312, QN 
                           => n6702);
   REGS_reg_5_0_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => n17310, QN 
                           => n6703);
   REGS_reg_4_23_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => n16892, QN
                           => n6648);
   REGS_reg_4_22_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => n16890, QN
                           => n6649);
   REGS_reg_4_21_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => n16888, QN
                           => n6650);
   REGS_reg_4_20_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => n16886, QN
                           => n6651);
   REGS_reg_4_19_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => n16884, QN
                           => n6652);
   REGS_reg_4_18_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => n16882, QN
                           => n6653);
   REGS_reg_4_17_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => n16880, QN
                           => n6654);
   REGS_reg_4_16_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => n16878, QN
                           => n6655);
   REGS_reg_4_15_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => n16876, QN
                           => n6656);
   REGS_reg_4_14_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => n16874, QN
                           => n6657);
   REGS_reg_4_13_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => n16872, QN
                           => n6658);
   REGS_reg_4_12_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => n16870, QN
                           => n6659);
   REGS_reg_4_11_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => n16868, QN
                           => n6660);
   REGS_reg_4_10_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => n16866, QN
                           => n6661);
   REGS_reg_4_9_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => n16864, QN 
                           => n6662);
   REGS_reg_4_8_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => n16862, QN 
                           => n6663);
   REGS_reg_4_7_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => n16860, QN 
                           => n6664);
   REGS_reg_4_6_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => n16858, QN 
                           => n6665);
   REGS_reg_4_5_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => n16856, QN 
                           => n6666);
   REGS_reg_4_4_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => n16854, QN 
                           => n6667);
   REGS_reg_4_3_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => n16852, QN 
                           => n6668);
   REGS_reg_4_2_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => n16850, QN 
                           => n6669);
   REGS_reg_4_1_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => n16848, QN 
                           => n6670);
   REGS_reg_4_0_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => n16846, QN 
                           => n6671);
   REGS_reg_3_23_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => n16836, QN
                           => n9026);
   REGS_reg_3_22_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => n16835, QN
                           => n9043);
   REGS_reg_3_21_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => n16834, QN
                           => n9060);
   REGS_reg_3_20_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => n16833, QN
                           => n9077);
   REGS_reg_3_19_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => n16832, QN
                           => n9094);
   REGS_reg_3_18_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => n16831, QN
                           => n9111);
   REGS_reg_3_17_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => n16830, QN
                           => n9128);
   REGS_reg_3_16_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => n16829, QN
                           => n9145);
   REGS_reg_3_15_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => n16828, QN
                           => n9162);
   REGS_reg_3_14_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => n16827, QN
                           => n9179);
   REGS_reg_3_13_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => n16826, QN
                           => n9196);
   REGS_reg_3_12_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => n16825, QN
                           => n9213);
   REGS_reg_3_11_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => n16824, QN
                           => n9230);
   REGS_reg_3_10_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => n16823, QN
                           => n9247);
   REGS_reg_3_9_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => n16822, QN 
                           => n9264);
   REGS_reg_3_8_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => n16821, QN 
                           => n9281);
   REGS_reg_3_7_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => n16820, QN 
                           => n9298);
   REGS_reg_3_6_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => n16819, QN 
                           => n9315);
   REGS_reg_3_5_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => n16818, QN 
                           => n9332);
   REGS_reg_3_4_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => n16817, QN 
                           => n9349);
   REGS_reg_3_3_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => n16816, QN 
                           => n9366);
   REGS_reg_3_2_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => n16815, QN 
                           => n9383);
   REGS_reg_3_1_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => n16814, QN 
                           => n9400);
   REGS_reg_3_0_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => n16813, QN 
                           => n9417);
   REGS_reg_2_23_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => n17300, QN
                           => n9025);
   REGS_reg_2_22_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => n17299, QN
                           => n9042);
   REGS_reg_2_21_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => n17298, QN
                           => n9059);
   REGS_reg_2_20_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => n17297, QN
                           => n9076);
   REGS_reg_2_19_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => n17296, QN
                           => n9093);
   REGS_reg_2_18_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => n17295, QN
                           => n9110);
   REGS_reg_2_17_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => n17294, QN
                           => n9127);
   REGS_reg_2_16_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => n17293, QN
                           => n9144);
   REGS_reg_2_15_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => n17292, QN
                           => n9161);
   REGS_reg_2_14_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => n17291, QN
                           => n9178);
   REGS_reg_2_13_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => n17290, QN
                           => n9195);
   REGS_reg_2_12_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => n17289, QN
                           => n9212);
   REGS_reg_2_11_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => n17288, QN
                           => n9229);
   REGS_reg_2_10_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => n17287, QN
                           => n9246);
   REGS_reg_2_9_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => n17286, QN 
                           => n9263);
   REGS_reg_2_8_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => n17285, QN 
                           => n9280);
   REGS_reg_2_7_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => n17284, QN 
                           => n9297);
   REGS_reg_2_6_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => n17283, QN 
                           => n9314);
   REGS_reg_2_5_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => n17282, QN 
                           => n9331);
   REGS_reg_2_4_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => n17281, QN 
                           => n9348);
   REGS_reg_2_3_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => n17280, QN 
                           => n9365);
   REGS_reg_2_2_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => n17279, QN 
                           => n9382);
   REGS_reg_2_1_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => n17278, QN 
                           => n9399);
   REGS_reg_2_0_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => n17277, QN 
                           => n9416);
   REGS_reg_16_31_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => n_1063, 
                           QN => n16812);
   REGS_reg_28_31_inst : DFF_X1 port map( D => n2720, CK => CLK, Q => n_1064, 
                           QN => n16804);
   REGS_reg_28_30_inst : DFF_X1 port map( D => n2719, CK => CLK, Q => n_1065, 
                           QN => n16803);
   REGS_reg_28_29_inst : DFF_X1 port map( D => n2718, CK => CLK, Q => n_1066, 
                           QN => n16802);
   REGS_reg_28_28_inst : DFF_X1 port map( D => n2717, CK => CLK, Q => n_1067, 
                           QN => n16801);
   REGS_reg_28_27_inst : DFF_X1 port map( D => n2716, CK => CLK, Q => n_1068, 
                           QN => n16800);
   REGS_reg_28_26_inst : DFF_X1 port map( D => n2715, CK => CLK, Q => n_1069, 
                           QN => n16799);
   REGS_reg_28_25_inst : DFF_X1 port map( D => n2714, CK => CLK, Q => n_1070, 
                           QN => n16798);
   REGS_reg_28_24_inst : DFF_X1 port map( D => n2713, CK => CLK, Q => n_1071, 
                           QN => n16797);
   REGS_reg_24_31_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => n_1072, 
                           QN => n16796);
   REGS_reg_24_30_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => n_1073, 
                           QN => n16795);
   REGS_reg_24_29_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => n_1074, 
                           QN => n16794);
   REGS_reg_24_28_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => n_1075, 
                           QN => n16793);
   REGS_reg_24_27_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => n_1076, 
                           QN => n16792);
   REGS_reg_24_26_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => n_1077, 
                           QN => n16791);
   REGS_reg_24_25_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => n_1078, 
                           QN => n16790);
   REGS_reg_24_24_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => n_1079, 
                           QN => n16789);
   REGS_reg_22_31_inst : DFF_X1 port map( D => n2912, CK => CLK, Q => n_1080, 
                           QN => n16788);
   REGS_reg_22_30_inst : DFF_X1 port map( D => n2911, CK => CLK, Q => n_1081, 
                           QN => n16787);
   REGS_reg_22_29_inst : DFF_X1 port map( D => n2910, CK => CLK, Q => n_1082, 
                           QN => n16786);
   REGS_reg_22_28_inst : DFF_X1 port map( D => n2909, CK => CLK, Q => n_1083, 
                           QN => n16785);
   REGS_reg_22_27_inst : DFF_X1 port map( D => n2908, CK => CLK, Q => n_1084, 
                           QN => n16784);
   REGS_reg_22_26_inst : DFF_X1 port map( D => n2907, CK => CLK, Q => n_1085, 
                           QN => n16783);
   REGS_reg_22_25_inst : DFF_X1 port map( D => n2906, CK => CLK, Q => n_1086, 
                           QN => n16782);
   REGS_reg_22_24_inst : DFF_X1 port map( D => n2905, CK => CLK, Q => n_1087, 
                           QN => n16781);
   REGS_reg_14_31_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => n_1088, 
                           QN => n16780);
   REGS_reg_14_30_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => n_1089, 
                           QN => n16779);
   REGS_reg_14_29_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => n_1090, 
                           QN => n16778);
   REGS_reg_14_28_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => n_1091, 
                           QN => n16777);
   REGS_reg_14_27_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => n_1092, 
                           QN => n16776);
   REGS_reg_14_26_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => n_1093, 
                           QN => n16775);
   REGS_reg_14_25_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => n_1094, 
                           QN => n16774);
   REGS_reg_14_24_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => n_1095, 
                           QN => n16773);
   REGS_reg_10_31_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => n_1096, 
                           QN => n16772);
   REGS_reg_10_30_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => n_1097, 
                           QN => n16771);
   REGS_reg_10_29_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => n_1098, 
                           QN => n16770);
   REGS_reg_10_28_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => n_1099, 
                           QN => n16769);
   REGS_reg_10_27_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => n_1100, 
                           QN => n16768);
   REGS_reg_10_26_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => n_1101, 
                           QN => n16767);
   REGS_reg_10_25_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => n_1102, 
                           QN => n16766);
   REGS_reg_10_24_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => n_1103, 
                           QN => n16765);
   REGS_reg_6_31_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => n_1104, QN
                           => n16764);
   REGS_reg_6_30_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => n_1105, QN
                           => n16763);
   REGS_reg_6_29_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => n_1106, QN
                           => n16762);
   REGS_reg_6_28_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => n_1107, QN
                           => n16761);
   REGS_reg_6_27_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => n_1108, QN
                           => n16760);
   REGS_reg_6_26_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => n_1109, QN
                           => n16759);
   REGS_reg_6_25_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => n_1110, QN
                           => n16758);
   REGS_reg_6_24_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => n_1111, QN
                           => n16757);
   REGS_reg_1_31_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => n_1112, QN
                           => n16756);
   REGS_reg_1_30_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => n_1113, QN
                           => n16755);
   REGS_reg_1_29_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => n_1114, QN
                           => n16754);
   REGS_reg_1_28_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => n_1115, QN
                           => n16753);
   REGS_reg_1_27_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => n_1116, QN
                           => n16752);
   REGS_reg_1_26_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => n_1117, QN
                           => n16751);
   REGS_reg_1_25_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => n_1118, QN
                           => n16750);
   REGS_reg_1_24_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => n_1119, QN
                           => n16749);
   REGS_reg_29_31_inst : DFF_X1 port map( D => n2688, CK => CLK, Q => n_1120, 
                           QN => n16548);
   REGS_reg_29_30_inst : DFF_X1 port map( D => n2687, CK => CLK, Q => n_1121, 
                           QN => n16547);
   REGS_reg_29_29_inst : DFF_X1 port map( D => n2686, CK => CLK, Q => n_1122, 
                           QN => n16546);
   REGS_reg_29_28_inst : DFF_X1 port map( D => n2685, CK => CLK, Q => n_1123, 
                           QN => n16545);
   REGS_reg_29_27_inst : DFF_X1 port map( D => n2684, CK => CLK, Q => n_1124, 
                           QN => n16544);
   REGS_reg_29_26_inst : DFF_X1 port map( D => n2683, CK => CLK, Q => n_1125, 
                           QN => n16543);
   REGS_reg_29_25_inst : DFF_X1 port map( D => n2682, CK => CLK, Q => n_1126, 
                           QN => n16542);
   REGS_reg_29_24_inst : DFF_X1 port map( D => n2681, CK => CLK, Q => n_1127, 
                           QN => n16541);
   REGS_reg_25_31_inst : DFF_X1 port map( D => n2816, CK => CLK, Q => n_1128, 
                           QN => n16540);
   REGS_reg_25_30_inst : DFF_X1 port map( D => n2815, CK => CLK, Q => n_1129, 
                           QN => n16539);
   REGS_reg_25_29_inst : DFF_X1 port map( D => n2814, CK => CLK, Q => n_1130, 
                           QN => n16538);
   REGS_reg_25_28_inst : DFF_X1 port map( D => n2813, CK => CLK, Q => n_1131, 
                           QN => n16537);
   REGS_reg_25_27_inst : DFF_X1 port map( D => n2812, CK => CLK, Q => n_1132, 
                           QN => n16536);
   REGS_reg_25_26_inst : DFF_X1 port map( D => n2811, CK => CLK, Q => n_1133, 
                           QN => n16535);
   REGS_reg_25_25_inst : DFF_X1 port map( D => n2810, CK => CLK, Q => n_1134, 
                           QN => n16534);
   REGS_reg_25_24_inst : DFF_X1 port map( D => n2809, CK => CLK, Q => n_1135, 
                           QN => n16533);
   REGS_reg_23_31_inst : DFF_X1 port map( D => n2880, CK => CLK, Q => n_1136, 
                           QN => n16532);
   REGS_reg_23_30_inst : DFF_X1 port map( D => n2879, CK => CLK, Q => n_1137, 
                           QN => n16531);
   REGS_reg_23_29_inst : DFF_X1 port map( D => n2878, CK => CLK, Q => n_1138, 
                           QN => n16530);
   REGS_reg_23_28_inst : DFF_X1 port map( D => n2877, CK => CLK, Q => n_1139, 
                           QN => n16529);
   REGS_reg_23_27_inst : DFF_X1 port map( D => n2876, CK => CLK, Q => n_1140, 
                           QN => n16528);
   REGS_reg_23_26_inst : DFF_X1 port map( D => n2875, CK => CLK, Q => n_1141, 
                           QN => n16527);
   REGS_reg_23_25_inst : DFF_X1 port map( D => n2874, CK => CLK, Q => n_1142, 
                           QN => n16526);
   REGS_reg_23_24_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => n_1143, 
                           QN => n16525);
   REGS_reg_15_31_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => n_1144, 
                           QN => n16524);
   REGS_reg_15_30_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => n_1145, 
                           QN => n16523);
   REGS_reg_15_29_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => n_1146, 
                           QN => n16522);
   REGS_reg_15_28_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => n_1147, 
                           QN => n16521);
   REGS_reg_15_27_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => n_1148, 
                           QN => n16520);
   REGS_reg_15_26_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => n_1149, 
                           QN => n16519);
   REGS_reg_15_25_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => n_1150, 
                           QN => n16518);
   REGS_reg_15_24_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => n_1151, 
                           QN => n16517);
   REGS_reg_11_31_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => n_1152, 
                           QN => n16516);
   REGS_reg_11_30_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => n_1153, 
                           QN => n16515);
   REGS_reg_11_29_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => n_1154, 
                           QN => n16514);
   REGS_reg_11_28_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => n_1155, 
                           QN => n16513);
   REGS_reg_11_27_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => n_1156, 
                           QN => n16512);
   REGS_reg_11_26_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => n_1157, 
                           QN => n16511);
   REGS_reg_11_25_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => n_1158, 
                           QN => n16510);
   REGS_reg_11_24_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => n_1159, 
                           QN => n16509);
   REGS_reg_7_31_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => n_1160, QN
                           => n16508);
   REGS_reg_7_30_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => n_1161, QN
                           => n16507);
   REGS_reg_7_29_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => n_1162, QN
                           => n16506);
   REGS_reg_7_28_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => n_1163, QN
                           => n16505);
   REGS_reg_7_27_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => n_1164, QN
                           => n16504);
   REGS_reg_7_26_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => n_1165, QN
                           => n16503);
   REGS_reg_7_25_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => n_1166, QN
                           => n16502);
   REGS_reg_7_24_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => n_1167, QN
                           => n16501);
   REGS_reg_0_31_inst : DFF_X1 port map( D => n3616, CK => CLK, Q => n_1168, QN
                           => n16500);
   REGS_reg_0_30_inst : DFF_X1 port map( D => n3615, CK => CLK, Q => n_1169, QN
                           => n16499);
   REGS_reg_0_29_inst : DFF_X1 port map( D => n3614, CK => CLK, Q => n_1170, QN
                           => n16498);
   REGS_reg_0_28_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => n_1171, QN
                           => n16497);
   REGS_reg_0_27_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => n_1172, QN
                           => n16496);
   REGS_reg_0_26_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => n_1173, QN
                           => n16495);
   REGS_reg_0_25_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => n_1174, QN
                           => n16494);
   REGS_reg_0_24_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => n_1175, QN
                           => n16493);
   REGS_reg_28_23_inst : DFF_X1 port map( D => n2712, CK => CLK, Q => n_1176, 
                           QN => n17220);
   REGS_reg_28_22_inst : DFF_X1 port map( D => n2711, CK => CLK, Q => n_1177, 
                           QN => n17219);
   REGS_reg_28_21_inst : DFF_X1 port map( D => n2710, CK => CLK, Q => n_1178, 
                           QN => n17218);
   REGS_reg_28_20_inst : DFF_X1 port map( D => n2709, CK => CLK, Q => n_1179, 
                           QN => n17217);
   REGS_reg_28_19_inst : DFF_X1 port map( D => n2708, CK => CLK, Q => n_1180, 
                           QN => n17216);
   REGS_reg_28_18_inst : DFF_X1 port map( D => n2707, CK => CLK, Q => n_1181, 
                           QN => n17215);
   REGS_reg_28_17_inst : DFF_X1 port map( D => n2706, CK => CLK, Q => n_1182, 
                           QN => n17214);
   REGS_reg_28_16_inst : DFF_X1 port map( D => n2705, CK => CLK, Q => n_1183, 
                           QN => n17213);
   REGS_reg_28_15_inst : DFF_X1 port map( D => n2704, CK => CLK, Q => n_1184, 
                           QN => n17212);
   REGS_reg_28_14_inst : DFF_X1 port map( D => n2703, CK => CLK, Q => n_1185, 
                           QN => n17211);
   REGS_reg_28_13_inst : DFF_X1 port map( D => n2702, CK => CLK, Q => n_1186, 
                           QN => n17210);
   REGS_reg_28_12_inst : DFF_X1 port map( D => n2701, CK => CLK, Q => n_1187, 
                           QN => n17209);
   REGS_reg_28_11_inst : DFF_X1 port map( D => n2700, CK => CLK, Q => n_1188, 
                           QN => n17208);
   REGS_reg_28_10_inst : DFF_X1 port map( D => n2699, CK => CLK, Q => n_1189, 
                           QN => n17207);
   REGS_reg_28_9_inst : DFF_X1 port map( D => n2698, CK => CLK, Q => n_1190, QN
                           => n17206);
   REGS_reg_28_8_inst : DFF_X1 port map( D => n2697, CK => CLK, Q => n_1191, QN
                           => n17205);
   REGS_reg_28_7_inst : DFF_X1 port map( D => n2696, CK => CLK, Q => n_1192, QN
                           => n17204);
   REGS_reg_28_6_inst : DFF_X1 port map( D => n2695, CK => CLK, Q => n_1193, QN
                           => n17203);
   REGS_reg_28_5_inst : DFF_X1 port map( D => n2694, CK => CLK, Q => n_1194, QN
                           => n17202);
   REGS_reg_28_4_inst : DFF_X1 port map( D => n2693, CK => CLK, Q => n_1195, QN
                           => n17201);
   REGS_reg_28_3_inst : DFF_X1 port map( D => n2692, CK => CLK, Q => n_1196, QN
                           => n17200);
   REGS_reg_28_2_inst : DFF_X1 port map( D => n2691, CK => CLK, Q => n_1197, QN
                           => n17199);
   REGS_reg_28_1_inst : DFF_X1 port map( D => n2690, CK => CLK, Q => n_1198, QN
                           => n17198);
   REGS_reg_28_0_inst : DFF_X1 port map( D => n2689, CK => CLK, Q => n_1199, QN
                           => n17197);
   REGS_reg_24_23_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => n_1200, 
                           QN => n17196);
   REGS_reg_24_22_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => n_1201, 
                           QN => n17195);
   REGS_reg_24_21_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => n_1202, 
                           QN => n17194);
   REGS_reg_24_20_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => n_1203, 
                           QN => n17193);
   REGS_reg_24_19_inst : DFF_X1 port map( D => n2836, CK => CLK, Q => n_1204, 
                           QN => n17192);
   REGS_reg_24_18_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => n_1205, 
                           QN => n17191);
   REGS_reg_24_17_inst : DFF_X1 port map( D => n2834, CK => CLK, Q => n_1206, 
                           QN => n17190);
   REGS_reg_24_16_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => n_1207, 
                           QN => n17189);
   REGS_reg_24_15_inst : DFF_X1 port map( D => n2832, CK => CLK, Q => n_1208, 
                           QN => n17188);
   REGS_reg_24_14_inst : DFF_X1 port map( D => n2831, CK => CLK, Q => n_1209, 
                           QN => n17187);
   REGS_reg_24_13_inst : DFF_X1 port map( D => n2830, CK => CLK, Q => n_1210, 
                           QN => n17186);
   REGS_reg_24_12_inst : DFF_X1 port map( D => n2829, CK => CLK, Q => n_1211, 
                           QN => n17185);
   REGS_reg_24_11_inst : DFF_X1 port map( D => n2828, CK => CLK, Q => n_1212, 
                           QN => n17184);
   REGS_reg_24_10_inst : DFF_X1 port map( D => n2827, CK => CLK, Q => n_1213, 
                           QN => n17183);
   REGS_reg_24_9_inst : DFF_X1 port map( D => n2826, CK => CLK, Q => n_1214, QN
                           => n17182);
   REGS_reg_24_8_inst : DFF_X1 port map( D => n2825, CK => CLK, Q => n_1215, QN
                           => n17181);
   REGS_reg_24_7_inst : DFF_X1 port map( D => n2824, CK => CLK, Q => n_1216, QN
                           => n17180);
   REGS_reg_24_6_inst : DFF_X1 port map( D => n2823, CK => CLK, Q => n_1217, QN
                           => n17179);
   REGS_reg_24_5_inst : DFF_X1 port map( D => n2822, CK => CLK, Q => n_1218, QN
                           => n17178);
   REGS_reg_24_4_inst : DFF_X1 port map( D => n2821, CK => CLK, Q => n_1219, QN
                           => n17177);
   REGS_reg_24_3_inst : DFF_X1 port map( D => n2820, CK => CLK, Q => n_1220, QN
                           => n17176);
   REGS_reg_24_2_inst : DFF_X1 port map( D => n2819, CK => CLK, Q => n_1221, QN
                           => n17175);
   REGS_reg_24_1_inst : DFF_X1 port map( D => n2818, CK => CLK, Q => n_1222, QN
                           => n17174);
   REGS_reg_24_0_inst : DFF_X1 port map( D => n2817, CK => CLK, Q => n_1223, QN
                           => n17173);
   REGS_reg_22_23_inst : DFF_X1 port map( D => n2904, CK => CLK, Q => n_1224, 
                           QN => n17172);
   REGS_reg_22_22_inst : DFF_X1 port map( D => n2903, CK => CLK, Q => n_1225, 
                           QN => n17171);
   REGS_reg_22_21_inst : DFF_X1 port map( D => n2902, CK => CLK, Q => n_1226, 
                           QN => n17170);
   REGS_reg_22_20_inst : DFF_X1 port map( D => n2901, CK => CLK, Q => n_1227, 
                           QN => n17169);
   REGS_reg_22_19_inst : DFF_X1 port map( D => n2900, CK => CLK, Q => n_1228, 
                           QN => n17168);
   REGS_reg_22_18_inst : DFF_X1 port map( D => n2899, CK => CLK, Q => n_1229, 
                           QN => n17167);
   REGS_reg_22_17_inst : DFF_X1 port map( D => n2898, CK => CLK, Q => n_1230, 
                           QN => n17166);
   REGS_reg_22_16_inst : DFF_X1 port map( D => n2897, CK => CLK, Q => n_1231, 
                           QN => n17165);
   REGS_reg_22_15_inst : DFF_X1 port map( D => n2896, CK => CLK, Q => n_1232, 
                           QN => n17164);
   REGS_reg_22_14_inst : DFF_X1 port map( D => n2895, CK => CLK, Q => n_1233, 
                           QN => n17163);
   REGS_reg_22_13_inst : DFF_X1 port map( D => n2894, CK => CLK, Q => n_1234, 
                           QN => n17162);
   REGS_reg_22_12_inst : DFF_X1 port map( D => n2893, CK => CLK, Q => n_1235, 
                           QN => n17161);
   REGS_reg_22_11_inst : DFF_X1 port map( D => n2892, CK => CLK, Q => n_1236, 
                           QN => n17160);
   REGS_reg_22_10_inst : DFF_X1 port map( D => n2891, CK => CLK, Q => n_1237, 
                           QN => n17159);
   REGS_reg_22_9_inst : DFF_X1 port map( D => n2890, CK => CLK, Q => n_1238, QN
                           => n17158);
   REGS_reg_22_8_inst : DFF_X1 port map( D => n2889, CK => CLK, Q => n_1239, QN
                           => n17157);
   REGS_reg_22_7_inst : DFF_X1 port map( D => n2888, CK => CLK, Q => n_1240, QN
                           => n17156);
   REGS_reg_22_6_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => n_1241, QN
                           => n17155);
   REGS_reg_22_5_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => n_1242, QN
                           => n17154);
   REGS_reg_22_4_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => n_1243, QN
                           => n17153);
   REGS_reg_22_3_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => n_1244, QN
                           => n17152);
   REGS_reg_22_2_inst : DFF_X1 port map( D => n2883, CK => CLK, Q => n_1245, QN
                           => n17151);
   REGS_reg_22_1_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => n_1246, QN
                           => n17150);
   REGS_reg_22_0_inst : DFF_X1 port map( D => n2881, CK => CLK, Q => n_1247, QN
                           => n17149);
   REGS_reg_14_23_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => n_1248, 
                           QN => n17148);
   REGS_reg_14_22_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => n_1249, 
                           QN => n17147);
   REGS_reg_14_21_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => n_1250, 
                           QN => n17146);
   REGS_reg_14_20_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => n_1251, 
                           QN => n17145);
   REGS_reg_14_19_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => n_1252, 
                           QN => n17144);
   REGS_reg_14_18_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => n_1253, 
                           QN => n17143);
   REGS_reg_14_17_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => n_1254, 
                           QN => n17142);
   REGS_reg_14_16_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => n_1255, 
                           QN => n17141);
   REGS_reg_14_15_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => n_1256, 
                           QN => n17140);
   REGS_reg_14_14_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => n_1257, 
                           QN => n17139);
   REGS_reg_14_13_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => n_1258, 
                           QN => n17138);
   REGS_reg_14_12_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => n_1259, 
                           QN => n17137);
   REGS_reg_14_11_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => n_1260, 
                           QN => n17136);
   REGS_reg_14_10_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => n_1261, 
                           QN => n17135);
   REGS_reg_14_9_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => n_1262, QN
                           => n17134);
   REGS_reg_14_8_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => n_1263, QN
                           => n17133);
   REGS_reg_14_7_inst : DFF_X1 port map( D => n3144, CK => CLK, Q => n_1264, QN
                           => n17132);
   REGS_reg_14_6_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => n_1265, QN
                           => n17131);
   REGS_reg_14_5_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => n_1266, QN
                           => n17130);
   REGS_reg_14_4_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => n_1267, QN
                           => n17129);
   REGS_reg_14_3_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => n_1268, QN
                           => n17128);
   REGS_reg_14_2_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => n_1269, QN
                           => n17127);
   REGS_reg_14_1_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => n_1270, QN
                           => n17126);
   REGS_reg_14_0_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => n_1271, QN
                           => n17125);
   REGS_reg_10_23_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => n_1272, 
                           QN => n17124);
   REGS_reg_10_22_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => n_1273, 
                           QN => n17123);
   REGS_reg_10_21_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => n_1274, 
                           QN => n17122);
   REGS_reg_10_20_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => n_1275, 
                           QN => n17121);
   REGS_reg_10_19_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => n_1276, 
                           QN => n17120);
   REGS_reg_10_18_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => n_1277, 
                           QN => n17119);
   REGS_reg_10_17_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => n_1278, 
                           QN => n17118);
   REGS_reg_10_16_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => n_1279, 
                           QN => n17117);
   REGS_reg_10_15_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => n_1280, 
                           QN => n17116);
   REGS_reg_10_14_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => n_1281, 
                           QN => n17115);
   REGS_reg_10_13_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => n_1282, 
                           QN => n17114);
   REGS_reg_10_12_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => n_1283, 
                           QN => n17113);
   REGS_reg_10_11_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => n_1284, 
                           QN => n17112);
   REGS_reg_10_10_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => n_1285, 
                           QN => n17111);
   REGS_reg_10_9_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => n_1286, QN
                           => n17110);
   REGS_reg_10_8_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => n_1287, QN
                           => n17109);
   REGS_reg_10_7_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => n_1288, QN
                           => n17108);
   REGS_reg_10_6_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => n_1289, QN
                           => n17107);
   REGS_reg_10_5_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => n_1290, QN
                           => n17106);
   REGS_reg_10_4_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => n_1291, QN
                           => n17105);
   REGS_reg_10_3_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => n_1292, QN
                           => n17104);
   REGS_reg_10_2_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => n_1293, QN
                           => n17103);
   REGS_reg_10_1_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => n_1294, QN
                           => n17102);
   REGS_reg_10_0_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => n_1295, QN
                           => n17101);
   REGS_reg_6_23_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => n_1296, QN
                           => n17100);
   REGS_reg_6_22_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => n_1297, QN
                           => n17099);
   REGS_reg_6_21_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => n_1298, QN
                           => n17098);
   REGS_reg_6_20_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => n_1299, QN
                           => n17097);
   REGS_reg_6_19_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => n_1300, QN
                           => n17096);
   REGS_reg_6_18_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => n_1301, QN
                           => n17095);
   REGS_reg_6_17_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => n_1302, QN
                           => n17094);
   REGS_reg_6_16_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => n_1303, QN
                           => n17093);
   REGS_reg_6_15_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => n_1304, QN
                           => n17092);
   REGS_reg_6_14_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => n_1305, QN
                           => n17091);
   REGS_reg_6_13_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => n_1306, QN
                           => n17090);
   REGS_reg_6_12_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => n_1307, QN
                           => n17089);
   REGS_reg_6_11_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => n_1308, QN
                           => n17088);
   REGS_reg_6_10_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => n_1309, QN
                           => n17087);
   REGS_reg_6_9_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => n_1310, QN 
                           => n17086);
   REGS_reg_6_8_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => n_1311, QN 
                           => n17085);
   REGS_reg_6_7_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => n_1312, QN 
                           => n17084);
   REGS_reg_6_6_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => n_1313, QN 
                           => n17083);
   REGS_reg_6_5_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => n_1314, QN 
                           => n17082);
   REGS_reg_6_4_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => n_1315, QN 
                           => n17081);
   REGS_reg_6_3_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => n_1316, QN 
                           => n17080);
   REGS_reg_6_2_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => n_1317, QN 
                           => n17079);
   REGS_reg_6_1_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => n_1318, QN 
                           => n17078);
   REGS_reg_6_0_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => n_1319, QN 
                           => n17077);
   REGS_reg_1_23_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => n_1320, QN
                           => n17076);
   REGS_reg_1_22_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => n_1321, QN
                           => n17075);
   REGS_reg_1_21_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => n_1322, QN
                           => n17074);
   REGS_reg_1_20_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => n_1323, QN
                           => n17073);
   REGS_reg_1_19_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => n_1324, QN
                           => n17072);
   REGS_reg_1_18_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => n_1325, QN
                           => n17071);
   REGS_reg_1_17_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => n_1326, QN
                           => n17070);
   REGS_reg_1_16_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => n_1327, QN
                           => n17069);
   REGS_reg_1_15_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => n_1328, QN
                           => n17068);
   REGS_reg_1_14_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => n_1329, QN
                           => n17067);
   REGS_reg_1_13_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => n_1330, QN
                           => n17066);
   REGS_reg_1_12_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => n_1331, QN
                           => n17065);
   REGS_reg_1_11_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => n_1332, QN
                           => n17064);
   REGS_reg_1_10_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => n_1333, QN
                           => n17063);
   REGS_reg_1_9_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => n_1334, QN 
                           => n17062);
   REGS_reg_1_8_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => n_1335, QN 
                           => n17061);
   REGS_reg_1_7_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => n_1336, QN 
                           => n17060);
   REGS_reg_1_6_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => n_1337, QN 
                           => n17059);
   REGS_reg_1_5_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => n_1338, QN 
                           => n17058);
   REGS_reg_1_4_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => n_1339, QN 
                           => n17057);
   REGS_reg_1_3_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => n_1340, QN 
                           => n17056);
   REGS_reg_1_2_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => n_1341, QN 
                           => n17055);
   REGS_reg_1_1_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => n_1342, QN 
                           => n17054);
   REGS_reg_1_0_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => n_1343, QN 
                           => n17053);
   REGS_reg_29_23_inst : DFF_X1 port map( D => n2680, CK => CLK, Q => n_1344, 
                           QN => n16632);
   REGS_reg_29_22_inst : DFF_X1 port map( D => n2679, CK => CLK, Q => n_1345, 
                           QN => n16631);
   REGS_reg_29_21_inst : DFF_X1 port map( D => n2678, CK => CLK, Q => n_1346, 
                           QN => n16630);
   REGS_reg_29_20_inst : DFF_X1 port map( D => n2677, CK => CLK, Q => n_1347, 
                           QN => n16629);
   REGS_reg_29_19_inst : DFF_X1 port map( D => n2676, CK => CLK, Q => n_1348, 
                           QN => n16628);
   REGS_reg_29_18_inst : DFF_X1 port map( D => n2675, CK => CLK, Q => n_1349, 
                           QN => n16627);
   REGS_reg_29_17_inst : DFF_X1 port map( D => n2674, CK => CLK, Q => n_1350, 
                           QN => n16626);
   REGS_reg_29_16_inst : DFF_X1 port map( D => n2673, CK => CLK, Q => n_1351, 
                           QN => n16625);
   REGS_reg_29_15_inst : DFF_X1 port map( D => n2672, CK => CLK, Q => n_1352, 
                           QN => n16624);
   REGS_reg_29_14_inst : DFF_X1 port map( D => n2671, CK => CLK, Q => n_1353, 
                           QN => n16623);
   REGS_reg_29_13_inst : DFF_X1 port map( D => n2670, CK => CLK, Q => n_1354, 
                           QN => n16622);
   REGS_reg_29_12_inst : DFF_X1 port map( D => n2669, CK => CLK, Q => n_1355, 
                           QN => n16621);
   REGS_reg_29_11_inst : DFF_X1 port map( D => n2668, CK => CLK, Q => n_1356, 
                           QN => n16736);
   REGS_reg_29_10_inst : DFF_X1 port map( D => n2667, CK => CLK, Q => n_1357, 
                           QN => n16735);
   REGS_reg_29_9_inst : DFF_X1 port map( D => n2666, CK => CLK, Q => n_1358, QN
                           => n16734);
   REGS_reg_29_8_inst : DFF_X1 port map( D => n2665, CK => CLK, Q => n_1359, QN
                           => n16733);
   REGS_reg_29_7_inst : DFF_X1 port map( D => n2664, CK => CLK, Q => n_1360, QN
                           => n16732);
   REGS_reg_29_6_inst : DFF_X1 port map( D => n2663, CK => CLK, Q => n_1361, QN
                           => n16731);
   REGS_reg_29_5_inst : DFF_X1 port map( D => n2662, CK => CLK, Q => n_1362, QN
                           => n16730);
   REGS_reg_29_4_inst : DFF_X1 port map( D => n2661, CK => CLK, Q => n_1363, QN
                           => n16729);
   REGS_reg_29_3_inst : DFF_X1 port map( D => n2660, CK => CLK, Q => n_1364, QN
                           => n16728);
   REGS_reg_29_2_inst : DFF_X1 port map( D => n2659, CK => CLK, Q => n_1365, QN
                           => n16727);
   REGS_reg_29_1_inst : DFF_X1 port map( D => n2658, CK => CLK, Q => n_1366, QN
                           => n16726);
   REGS_reg_29_0_inst : DFF_X1 port map( D => n2657, CK => CLK, Q => n_1367, QN
                           => n16725);
   REGS_reg_25_23_inst : DFF_X1 port map( D => n2808, CK => CLK, Q => n_1368, 
                           QN => n16620);
   REGS_reg_25_22_inst : DFF_X1 port map( D => n2807, CK => CLK, Q => n_1369, 
                           QN => n16619);
   REGS_reg_25_21_inst : DFF_X1 port map( D => n2806, CK => CLK, Q => n_1370, 
                           QN => n16618);
   REGS_reg_25_20_inst : DFF_X1 port map( D => n2805, CK => CLK, Q => n_1371, 
                           QN => n16617);
   REGS_reg_25_19_inst : DFF_X1 port map( D => n2804, CK => CLK, Q => n_1372, 
                           QN => n16616);
   REGS_reg_25_18_inst : DFF_X1 port map( D => n2803, CK => CLK, Q => n_1373, 
                           QN => n16615);
   REGS_reg_25_17_inst : DFF_X1 port map( D => n2802, CK => CLK, Q => n_1374, 
                           QN => n16614);
   REGS_reg_25_16_inst : DFF_X1 port map( D => n2801, CK => CLK, Q => n_1375, 
                           QN => n16613);
   REGS_reg_25_15_inst : DFF_X1 port map( D => n2800, CK => CLK, Q => n_1376, 
                           QN => n16612);
   REGS_reg_25_14_inst : DFF_X1 port map( D => n2799, CK => CLK, Q => n_1377, 
                           QN => n16611);
   REGS_reg_25_13_inst : DFF_X1 port map( D => n2798, CK => CLK, Q => n_1378, 
                           QN => n16610);
   REGS_reg_25_12_inst : DFF_X1 port map( D => n2797, CK => CLK, Q => n_1379, 
                           QN => n16609);
   REGS_reg_25_11_inst : DFF_X1 port map( D => n2796, CK => CLK, Q => n_1380, 
                           QN => n16724);
   REGS_reg_25_10_inst : DFF_X1 port map( D => n2795, CK => CLK, Q => n_1381, 
                           QN => n16723);
   REGS_reg_25_9_inst : DFF_X1 port map( D => n2794, CK => CLK, Q => n_1382, QN
                           => n16722);
   REGS_reg_25_8_inst : DFF_X1 port map( D => n2793, CK => CLK, Q => n_1383, QN
                           => n16721);
   REGS_reg_25_7_inst : DFF_X1 port map( D => n2792, CK => CLK, Q => n_1384, QN
                           => n16720);
   REGS_reg_25_6_inst : DFF_X1 port map( D => n2791, CK => CLK, Q => n_1385, QN
                           => n16719);
   REGS_reg_25_5_inst : DFF_X1 port map( D => n2790, CK => CLK, Q => n_1386, QN
                           => n16718);
   REGS_reg_25_4_inst : DFF_X1 port map( D => n2789, CK => CLK, Q => n_1387, QN
                           => n16717);
   REGS_reg_25_3_inst : DFF_X1 port map( D => n2788, CK => CLK, Q => n_1388, QN
                           => n16716);
   REGS_reg_25_2_inst : DFF_X1 port map( D => n2787, CK => CLK, Q => n_1389, QN
                           => n16715);
   REGS_reg_25_1_inst : DFF_X1 port map( D => n2786, CK => CLK, Q => n_1390, QN
                           => n16714);
   REGS_reg_25_0_inst : DFF_X1 port map( D => n2785, CK => CLK, Q => n_1391, QN
                           => n16713);
   REGS_reg_23_23_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => n_1392, 
                           QN => n16608);
   REGS_reg_23_22_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => n_1393, 
                           QN => n16607);
   REGS_reg_23_21_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => n_1394, 
                           QN => n16606);
   REGS_reg_23_20_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => n_1395, 
                           QN => n16605);
   REGS_reg_23_19_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => n_1396, 
                           QN => n16604);
   REGS_reg_23_18_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => n_1397, 
                           QN => n16603);
   REGS_reg_23_17_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => n_1398, 
                           QN => n16602);
   REGS_reg_23_16_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => n_1399, 
                           QN => n16601);
   REGS_reg_23_15_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => n_1400, 
                           QN => n16600);
   REGS_reg_23_14_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => n_1401, 
                           QN => n16599);
   REGS_reg_23_13_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => n_1402, 
                           QN => n16598);
   REGS_reg_23_12_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => n_1403, 
                           QN => n16597);
   REGS_reg_23_11_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => n_1404, 
                           QN => n16712);
   REGS_reg_23_10_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => n_1405, 
                           QN => n16711);
   REGS_reg_23_9_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => n_1406, QN
                           => n16710);
   REGS_reg_23_8_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => n_1407, QN
                           => n16709);
   REGS_reg_23_7_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => n_1408, QN
                           => n16708);
   REGS_reg_23_6_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => n_1409, QN
                           => n16707);
   REGS_reg_23_5_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => n_1410, QN
                           => n16706);
   REGS_reg_23_4_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => n_1411, QN
                           => n16705);
   REGS_reg_23_3_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => n_1412, QN
                           => n16704);
   REGS_reg_23_2_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => n_1413, QN
                           => n16703);
   REGS_reg_23_1_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => n_1414, QN
                           => n16702);
   REGS_reg_23_0_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => n_1415, QN
                           => n16701);
   REGS_reg_15_23_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => n_1416, 
                           QN => n16596);
   REGS_reg_15_22_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => n_1417, 
                           QN => n16595);
   REGS_reg_15_21_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => n_1418, 
                           QN => n16594);
   REGS_reg_15_20_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => n_1419, 
                           QN => n16593);
   REGS_reg_15_19_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => n_1420, 
                           QN => n16592);
   REGS_reg_15_18_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => n_1421, 
                           QN => n16591);
   REGS_reg_15_17_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => n_1422, 
                           QN => n16590);
   REGS_reg_15_16_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => n_1423, 
                           QN => n16589);
   REGS_reg_15_15_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => n_1424, 
                           QN => n16588);
   REGS_reg_15_14_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => n_1425, 
                           QN => n16587);
   REGS_reg_15_13_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => n_1426, 
                           QN => n16586);
   REGS_reg_15_12_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => n_1427, 
                           QN => n16585);
   REGS_reg_15_11_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => n_1428, 
                           QN => n16700);
   REGS_reg_15_10_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => n_1429, 
                           QN => n16699);
   REGS_reg_15_9_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => n_1430, QN
                           => n16698);
   REGS_reg_15_8_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => n_1431, QN
                           => n16697);
   REGS_reg_15_7_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => n_1432, QN
                           => n16696);
   REGS_reg_15_6_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => n_1433, QN
                           => n16695);
   REGS_reg_15_5_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => n_1434, QN
                           => n16694);
   REGS_reg_15_4_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => n_1435, QN
                           => n16693);
   REGS_reg_15_3_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => n_1436, QN
                           => n16692);
   REGS_reg_15_2_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => n_1437, QN
                           => n16691);
   REGS_reg_15_1_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => n_1438, QN
                           => n16690);
   REGS_reg_15_0_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => n_1439, QN
                           => n16689);
   REGS_reg_11_23_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => n_1440, 
                           QN => n16584);
   REGS_reg_11_22_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => n_1441, 
                           QN => n16583);
   REGS_reg_11_21_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => n_1442, 
                           QN => n16582);
   REGS_reg_11_20_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => n_1443, 
                           QN => n16581);
   REGS_reg_11_19_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => n_1444, 
                           QN => n16580);
   REGS_reg_11_18_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => n_1445, 
                           QN => n16579);
   REGS_reg_11_17_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => n_1446, 
                           QN => n16578);
   REGS_reg_11_16_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => n_1447, 
                           QN => n16577);
   REGS_reg_11_15_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => n_1448, 
                           QN => n16576);
   REGS_reg_11_14_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => n_1449, 
                           QN => n16575);
   REGS_reg_11_13_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => n_1450, 
                           QN => n16574);
   REGS_reg_11_12_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => n_1451, 
                           QN => n16573);
   REGS_reg_11_11_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => n_1452, 
                           QN => n16688);
   REGS_reg_11_10_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => n_1453, 
                           QN => n16687);
   REGS_reg_11_9_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => n_1454, QN
                           => n16686);
   REGS_reg_11_8_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => n_1455, QN
                           => n16685);
   REGS_reg_11_7_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => n_1456, QN
                           => n16684);
   REGS_reg_11_6_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => n_1457, QN
                           => n16683);
   REGS_reg_11_5_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => n_1458, QN
                           => n16682);
   REGS_reg_11_4_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => n_1459, QN
                           => n16681);
   REGS_reg_11_3_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => n_1460, QN
                           => n16680);
   REGS_reg_11_2_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => n_1461, QN
                           => n16679);
   REGS_reg_11_1_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => n_1462, QN
                           => n16678);
   REGS_reg_11_0_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => n_1463, QN
                           => n16677);
   REGS_reg_7_23_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => n_1464, QN
                           => n16572);
   REGS_reg_7_22_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => n_1465, QN
                           => n16571);
   REGS_reg_7_21_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => n_1466, QN
                           => n16570);
   REGS_reg_7_20_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => n_1467, QN
                           => n16569);
   REGS_reg_7_19_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => n_1468, QN
                           => n16568);
   REGS_reg_7_18_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => n_1469, QN
                           => n16567);
   REGS_reg_7_17_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => n_1470, QN
                           => n16566);
   REGS_reg_7_16_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => n_1471, QN
                           => n16565);
   REGS_reg_7_15_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => n_1472, QN
                           => n16564);
   REGS_reg_7_14_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => n_1473, QN
                           => n16563);
   REGS_reg_7_13_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => n_1474, QN
                           => n16562);
   REGS_reg_7_12_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => n_1475, QN
                           => n16561);
   REGS_reg_7_11_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => n_1476, QN
                           => n16676);
   REGS_reg_7_10_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => n_1477, QN
                           => n16675);
   REGS_reg_7_9_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => n_1478, QN 
                           => n16674);
   REGS_reg_7_8_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => n_1479, QN 
                           => n16673);
   REGS_reg_7_7_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => n_1480, QN 
                           => n16672);
   REGS_reg_7_6_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => n_1481, QN 
                           => n16671);
   REGS_reg_7_5_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => n_1482, QN 
                           => n16670);
   REGS_reg_7_4_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => n_1483, QN 
                           => n16669);
   REGS_reg_7_3_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => n_1484, QN 
                           => n16668);
   REGS_reg_7_2_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => n_1485, QN 
                           => n16667);
   REGS_reg_7_1_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => n_1486, QN 
                           => n16666);
   REGS_reg_7_0_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => n_1487, QN 
                           => n16665);
   REGS_reg_0_23_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => n_1488, QN
                           => n16560);
   REGS_reg_0_22_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => n_1489, QN
                           => n16559);
   REGS_reg_0_21_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => n_1490, QN
                           => n16558);
   REGS_reg_0_20_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => n_1491, QN
                           => n16557);
   REGS_reg_0_19_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => n_1492, QN
                           => n16556);
   REGS_reg_0_18_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => n_1493, QN
                           => n16555);
   REGS_reg_0_17_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => n_1494, QN
                           => n16554);
   REGS_reg_0_16_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => n_1495, QN
                           => n16553);
   REGS_reg_0_15_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => n_1496, QN
                           => n16552);
   REGS_reg_0_14_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => n_1497, QN
                           => n16551);
   REGS_reg_0_13_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => n_1498, QN
                           => n16550);
   REGS_reg_0_12_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => n_1499, QN
                           => n16549);
   REGS_reg_0_11_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => n_1500, QN
                           => n16664);
   REGS_reg_0_10_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => n_1501, QN
                           => n16663);
   REGS_reg_0_9_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => n_1502, QN 
                           => n16662);
   REGS_reg_0_8_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => n_1503, QN 
                           => n16661);
   REGS_reg_0_7_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => n_1504, QN 
                           => n16660);
   REGS_reg_0_6_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => n_1505, QN 
                           => n16659);
   REGS_reg_0_5_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => n_1506, QN 
                           => n16658);
   REGS_reg_0_4_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => n_1507, QN 
                           => n16657);
   REGS_reg_0_3_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => n_1508, QN 
                           => n16656);
   REGS_reg_0_2_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => n_1509, QN 
                           => n16655);
   REGS_reg_0_1_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => n_1510, QN 
                           => n16654);
   REGS_reg_0_0_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => n_1511, QN 
                           => n16653);
   REGS_reg_18_31_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => n12483, 
                           QN => n17044);
   REGS_reg_18_30_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => n12482, 
                           QN => n17043);
   REGS_reg_18_29_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => n12481, 
                           QN => n17042);
   REGS_reg_18_28_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => n12480, 
                           QN => n17041);
   REGS_reg_18_27_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => n12479, 
                           QN => n17040);
   REGS_reg_18_26_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => n12478, 
                           QN => n17039);
   REGS_reg_18_25_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => n12477, 
                           QN => n17038);
   REGS_reg_18_24_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => n12476, 
                           QN => n17037);
   REGS_reg_18_23_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => n12721, 
                           QN => n17492);
   REGS_reg_18_22_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => n12720, 
                           QN => n17491);
   REGS_reg_18_21_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => n12719, 
                           QN => n17490);
   REGS_reg_18_20_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => n12718, 
                           QN => n17489);
   REGS_reg_18_19_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => n12717, 
                           QN => n17488);
   REGS_reg_18_18_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => n12716, 
                           QN => n17487);
   REGS_reg_18_17_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => n12715, 
                           QN => n17486);
   REGS_reg_18_16_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => n12714, 
                           QN => n17485);
   REGS_reg_18_15_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => n12713, 
                           QN => n17484);
   REGS_reg_18_14_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => n12712, 
                           QN => n17483);
   REGS_reg_18_13_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => n12711, 
                           QN => n17482);
   REGS_reg_18_12_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => n12710, 
                           QN => n17481);
   REGS_reg_18_11_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => n12709, 
                           QN => n17480);
   REGS_reg_18_10_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => n12708, 
                           QN => n17479);
   REGS_reg_18_9_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => n12707, QN
                           => n17478);
   REGS_reg_18_8_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => n12706, QN
                           => n17477);
   REGS_reg_18_7_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => n12705, QN
                           => n17476);
   REGS_reg_18_6_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => n12704, QN
                           => n17475);
   REGS_reg_18_5_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => n12703, QN
                           => n17474);
   REGS_reg_18_4_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => n12702, QN
                           => n17473);
   REGS_reg_18_3_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => n12701, QN
                           => n17472);
   REGS_reg_18_2_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => n12700, QN
                           => n17471);
   REGS_reg_18_1_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => n12699, QN
                           => n17470);
   REGS_reg_18_0_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => n12698, QN
                           => n17469);
   REGS_reg_19_31_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => n12475, 
                           QN => n17052);
   REGS_reg_19_30_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => n12474, 
                           QN => n17051);
   REGS_reg_19_29_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => n12473, 
                           QN => n17050);
   REGS_reg_19_28_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => n12472, 
                           QN => n17049);
   REGS_reg_19_27_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => n12471, 
                           QN => n17048);
   REGS_reg_19_26_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => n12470, 
                           QN => n17047);
   REGS_reg_19_25_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => n12469, 
                           QN => n17046);
   REGS_reg_19_24_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => n12468, 
                           QN => n17045);
   REGS_reg_19_23_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => n12697, 
                           QN => n17516);
   REGS_reg_19_22_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => n12696, 
                           QN => n17515);
   REGS_reg_19_21_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => n12695, 
                           QN => n17514);
   REGS_reg_19_20_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => n12694, 
                           QN => n17513);
   REGS_reg_19_19_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => n12693, 
                           QN => n17512);
   REGS_reg_19_18_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => n12692, 
                           QN => n17511);
   REGS_reg_19_17_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => n12691, 
                           QN => n17510);
   REGS_reg_19_16_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => n12690, 
                           QN => n17509);
   REGS_reg_19_15_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => n12689, 
                           QN => n17508);
   REGS_reg_19_14_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => n12688, 
                           QN => n17507);
   REGS_reg_19_13_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => n12687, 
                           QN => n17506);
   REGS_reg_19_12_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => n12686, 
                           QN => n17505);
   REGS_reg_19_11_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => n12685, 
                           QN => n17504);
   REGS_reg_19_10_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => n12684, 
                           QN => n17503);
   REGS_reg_19_9_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => n12683, QN
                           => n17502);
   REGS_reg_19_8_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => n12682, QN
                           => n17501);
   REGS_reg_19_7_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => n12681, QN
                           => n17500);
   REGS_reg_19_6_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => n12680, QN
                           => n17499);
   REGS_reg_19_5_inst : DFF_X1 port map( D => n2982, CK => CLK, Q => n12679, QN
                           => n17498);
   REGS_reg_19_4_inst : DFF_X1 port map( D => n2981, CK => CLK, Q => n12678, QN
                           => n17497);
   REGS_reg_19_3_inst : DFF_X1 port map( D => n2980, CK => CLK, Q => n12677, QN
                           => n17496);
   REGS_reg_19_2_inst : DFF_X1 port map( D => n2979, CK => CLK, Q => n12676, QN
                           => n17495);
   REGS_reg_19_1_inst : DFF_X1 port map( D => n2978, CK => CLK, Q => n12675, QN
                           => n17494);
   REGS_reg_19_0_inst : DFF_X1 port map( D => n2977, CK => CLK, Q => n12674, QN
                           => n17493);
   U13060 : NAND3_X1 port map( A1 => n13561, A2 => n13560, A3 => n14647, ZN => 
                           n14630);
   U13061 : NAND3_X1 port map( A1 => n14647, A2 => n13560, A3 => ADDR_WR(3), ZN
                           => n14649);
   U13062 : NAND3_X1 port map( A1 => n14647, A2 => n13561, A3 => ADDR_WR(4), ZN
                           => n14658);
   U13063 : NAND3_X1 port map( A1 => n13563, A2 => n13562, A3 => n13564, ZN => 
                           n14631);
   U13064 : NAND3_X1 port map( A1 => n13563, A2 => n13562, A3 => ADDR_WR(0), ZN
                           => n14634);
   U13065 : NAND3_X1 port map( A1 => n13564, A2 => n13562, A3 => ADDR_WR(1), ZN
                           => n14636);
   U13066 : NAND3_X1 port map( A1 => ADDR_WR(0), A2 => n13562, A3 => ADDR_WR(1)
                           , ZN => n14638);
   U13067 : NAND3_X1 port map( A1 => n13564, A2 => n13563, A3 => ADDR_WR(2), ZN
                           => n14640);
   U13068 : NAND3_X1 port map( A1 => ADDR_WR(0), A2 => n13563, A3 => ADDR_WR(2)
                           , ZN => n14642);
   U13069 : NAND3_X1 port map( A1 => ADDR_WR(1), A2 => n13564, A3 => ADDR_WR(2)
                           , ZN => n14644);
   U13070 : NAND3_X1 port map( A1 => ADDR_WR(3), A2 => n14647, A3 => ADDR_WR(4)
                           , ZN => n14667);
   U13071 : NAND3_X1 port map( A1 => ADDR_WR(1), A2 => ADDR_WR(0), A3 => 
                           ADDR_WR(2), ZN => n14646);
   U13072 : NOR2_X1 port map( A1 => ADDR_RD2(1), A2 => ADDR_RD2(2), ZN => 
                           n15959);
   U13073 : NOR2_X1 port map( A1 => ADDR_RD1(1), A2 => ADDR_RD1(2), ZN => 
                           n15306);
   U13074 : INV_X1 port map( A => n18104, ZN => n18097);
   U13075 : INV_X1 port map( A => n17990, ZN => n17983);
   U13076 : INV_X1 port map( A => n17981, ZN => n17974);
   U13077 : INV_X1 port map( A => n17972, ZN => n17965);
   U13078 : INV_X1 port map( A => n17963, ZN => n17956);
   U13079 : INV_X1 port map( A => n17936, ZN => n17929);
   U13080 : INV_X1 port map( A => n17927, ZN => n17920);
   U13081 : INV_X1 port map( A => n17900, ZN => n17893);
   U13082 : INV_X1 port map( A => n17891, ZN => n17884);
   U13083 : INV_X1 port map( A => n17828, ZN => n17821);
   U13084 : INV_X1 port map( A => n17819, ZN => n17812);
   U13085 : INV_X1 port map( A => n17774, ZN => n17767);
   U13086 : INV_X1 port map( A => n17765, ZN => n17758);
   U13087 : INV_X1 port map( A => n17738, ZN => n17731);
   U13088 : INV_X1 port map( A => n17837, ZN => n17830);
   U13089 : INV_X1 port map( A => n17846, ZN => n17839);
   U13090 : INV_X1 port map( A => n17945, ZN => n17938);
   U13091 : INV_X1 port map( A => n17909, ZN => n17902);
   U13092 : INV_X1 port map( A => n17873, ZN => n17866);
   U13093 : INV_X1 port map( A => n17801, ZN => n17794);
   U13094 : INV_X1 port map( A => n17783, ZN => n17776);
   U13095 : INV_X1 port map( A => n17747, ZN => n17740);
   U13096 : INV_X1 port map( A => n17999, ZN => n17992);
   U13097 : INV_X1 port map( A => n17954, ZN => n17947);
   U13098 : INV_X1 port map( A => n17918, ZN => n17911);
   U13099 : INV_X1 port map( A => n17882, ZN => n17875);
   U13100 : INV_X1 port map( A => n17810, ZN => n17803);
   U13101 : INV_X1 port map( A => n17792, ZN => n17785);
   U13102 : INV_X1 port map( A => n17756, ZN => n17749);
   U13103 : INV_X1 port map( A => n17864, ZN => n17857);
   U13104 : INV_X1 port map( A => n17855, ZN => n17848);
   U13105 : BUF_X1 port map( A => n18105, Z => n18098);
   U13106 : BUF_X1 port map( A => n18105, Z => n18099);
   U13107 : BUF_X1 port map( A => n18105, Z => n18100);
   U13108 : BUF_X1 port map( A => n18105, Z => n18101);
   U13109 : BUF_X1 port map( A => n18105, Z => n18102);
   U13110 : BUF_X1 port map( A => n18105, Z => n18103);
   U13111 : BUF_X1 port map( A => n18105, Z => n18104);
   U13112 : BUF_X1 port map( A => n17730, Z => n17722);
   U13113 : BUF_X1 port map( A => n17730, Z => n17723);
   U13114 : BUF_X1 port map( A => n17730, Z => n17724);
   U13115 : BUF_X1 port map( A => n17730, Z => n17725);
   U13116 : BUF_X1 port map( A => n17730, Z => n17726);
   U13117 : BUF_X1 port map( A => n17730, Z => n17727);
   U13118 : BUF_X1 port map( A => n17727, Z => n17728);
   U13119 : BUF_X1 port map( A => n17722, Z => n17729);
   U13120 : BUF_X1 port map( A => n15339, Z => n17604);
   U13121 : BUF_X1 port map( A => n15344, Z => n17592);
   U13122 : BUF_X1 port map( A => n15349, Z => n17580);
   U13123 : BUF_X1 port map( A => n15354, Z => n17568);
   U13124 : BUF_X1 port map( A => n15363, Z => n17556);
   U13125 : BUF_X1 port map( A => n15368, Z => n17544);
   U13126 : BUF_X1 port map( A => n15373, Z => n17532);
   U13127 : BUF_X1 port map( A => n15378, Z => n17520);
   U13128 : BUF_X1 port map( A => n15339, Z => n17605);
   U13129 : BUF_X1 port map( A => n15344, Z => n17593);
   U13130 : BUF_X1 port map( A => n15349, Z => n17581);
   U13131 : BUF_X1 port map( A => n15354, Z => n17569);
   U13132 : BUF_X1 port map( A => n15363, Z => n17557);
   U13133 : BUF_X1 port map( A => n15368, Z => n17545);
   U13134 : BUF_X1 port map( A => n15373, Z => n17533);
   U13135 : BUF_X1 port map( A => n15378, Z => n17521);
   U13136 : BUF_X1 port map( A => n14686, Z => n17706);
   U13137 : BUF_X1 port map( A => n14691, Z => n17694);
   U13138 : BUF_X1 port map( A => n14696, Z => n17682);
   U13139 : BUF_X1 port map( A => n14701, Z => n17670);
   U13140 : BUF_X1 port map( A => n14710, Z => n17658);
   U13141 : BUF_X1 port map( A => n14715, Z => n17646);
   U13142 : BUF_X1 port map( A => n14720, Z => n17634);
   U13143 : BUF_X1 port map( A => n14725, Z => n17622);
   U13144 : BUF_X1 port map( A => n14686, Z => n17707);
   U13145 : BUF_X1 port map( A => n14691, Z => n17695);
   U13146 : BUF_X1 port map( A => n14696, Z => n17683);
   U13147 : BUF_X1 port map( A => n14701, Z => n17671);
   U13148 : BUF_X1 port map( A => n14710, Z => n17659);
   U13149 : BUF_X1 port map( A => n14715, Z => n17647);
   U13150 : BUF_X1 port map( A => n14720, Z => n17635);
   U13151 : BUF_X1 port map( A => n14725, Z => n17623);
   U13152 : BUF_X1 port map( A => n15340, Z => n17601);
   U13153 : BUF_X1 port map( A => n15345, Z => n17589);
   U13154 : BUF_X1 port map( A => n15350, Z => n17577);
   U13155 : BUF_X1 port map( A => n15355, Z => n17565);
   U13156 : BUF_X1 port map( A => n15364, Z => n17553);
   U13157 : BUF_X1 port map( A => n15369, Z => n17541);
   U13158 : BUF_X1 port map( A => n15374, Z => n17529);
   U13159 : BUF_X1 port map( A => n15379, Z => n17517);
   U13160 : BUF_X1 port map( A => n15340, Z => n17602);
   U13161 : BUF_X1 port map( A => n15345, Z => n17590);
   U13162 : BUF_X1 port map( A => n15350, Z => n17578);
   U13163 : BUF_X1 port map( A => n15355, Z => n17566);
   U13164 : BUF_X1 port map( A => n15364, Z => n17554);
   U13165 : BUF_X1 port map( A => n15369, Z => n17542);
   U13166 : BUF_X1 port map( A => n15374, Z => n17530);
   U13167 : BUF_X1 port map( A => n15379, Z => n17518);
   U13168 : BUF_X1 port map( A => n14687, Z => n17703);
   U13169 : BUF_X1 port map( A => n14692, Z => n17691);
   U13170 : BUF_X1 port map( A => n14697, Z => n17679);
   U13171 : BUF_X1 port map( A => n14702, Z => n17667);
   U13172 : BUF_X1 port map( A => n14711, Z => n17655);
   U13173 : BUF_X1 port map( A => n14716, Z => n17643);
   U13174 : BUF_X1 port map( A => n14721, Z => n17631);
   U13175 : BUF_X1 port map( A => n14726, Z => n17619);
   U13176 : BUF_X1 port map( A => n14687, Z => n17704);
   U13177 : BUF_X1 port map( A => n14692, Z => n17692);
   U13178 : BUF_X1 port map( A => n14697, Z => n17680);
   U13179 : BUF_X1 port map( A => n14702, Z => n17668);
   U13180 : BUF_X1 port map( A => n14711, Z => n17656);
   U13181 : BUF_X1 port map( A => n14716, Z => n17644);
   U13182 : BUF_X1 port map( A => n14721, Z => n17632);
   U13183 : BUF_X1 port map( A => n14726, Z => n17620);
   U13184 : BUF_X1 port map( A => n15336, Z => n17610);
   U13185 : BUF_X1 port map( A => n15341, Z => n17598);
   U13186 : BUF_X1 port map( A => n15346, Z => n17586);
   U13187 : BUF_X1 port map( A => n15351, Z => n17574);
   U13188 : BUF_X1 port map( A => n15360, Z => n17562);
   U13189 : BUF_X1 port map( A => n15365, Z => n17550);
   U13190 : BUF_X1 port map( A => n15370, Z => n17538);
   U13191 : BUF_X1 port map( A => n15375, Z => n17526);
   U13192 : BUF_X1 port map( A => n15336, Z => n17611);
   U13193 : BUF_X1 port map( A => n15341, Z => n17599);
   U13194 : BUF_X1 port map( A => n15346, Z => n17587);
   U13195 : BUF_X1 port map( A => n15351, Z => n17575);
   U13196 : BUF_X1 port map( A => n15360, Z => n17563);
   U13197 : BUF_X1 port map( A => n15365, Z => n17551);
   U13198 : BUF_X1 port map( A => n15370, Z => n17539);
   U13199 : BUF_X1 port map( A => n15375, Z => n17527);
   U13200 : BUF_X1 port map( A => n14683, Z => n17712);
   U13201 : BUF_X1 port map( A => n14688, Z => n17700);
   U13202 : BUF_X1 port map( A => n14693, Z => n17688);
   U13203 : BUF_X1 port map( A => n14698, Z => n17676);
   U13204 : BUF_X1 port map( A => n14707, Z => n17664);
   U13205 : BUF_X1 port map( A => n14712, Z => n17652);
   U13206 : BUF_X1 port map( A => n14717, Z => n17640);
   U13207 : BUF_X1 port map( A => n14722, Z => n17628);
   U13208 : BUF_X1 port map( A => n14683, Z => n17713);
   U13209 : BUF_X1 port map( A => n14688, Z => n17701);
   U13210 : BUF_X1 port map( A => n14693, Z => n17689);
   U13211 : BUF_X1 port map( A => n14698, Z => n17677);
   U13212 : BUF_X1 port map( A => n14707, Z => n17665);
   U13213 : BUF_X1 port map( A => n14712, Z => n17653);
   U13214 : BUF_X1 port map( A => n14717, Z => n17641);
   U13215 : BUF_X1 port map( A => n14722, Z => n17629);
   U13216 : BUF_X1 port map( A => n15337, Z => n17607);
   U13217 : BUF_X1 port map( A => n15342, Z => n17595);
   U13218 : BUF_X1 port map( A => n15347, Z => n17583);
   U13219 : BUF_X1 port map( A => n15352, Z => n17571);
   U13220 : BUF_X1 port map( A => n15361, Z => n17559);
   U13221 : BUF_X1 port map( A => n15366, Z => n17547);
   U13222 : BUF_X1 port map( A => n15371, Z => n17535);
   U13223 : BUF_X1 port map( A => n15376, Z => n17523);
   U13224 : BUF_X1 port map( A => n15337, Z => n17608);
   U13225 : BUF_X1 port map( A => n15342, Z => n17596);
   U13226 : BUF_X1 port map( A => n15347, Z => n17584);
   U13227 : BUF_X1 port map( A => n15352, Z => n17572);
   U13228 : BUF_X1 port map( A => n15361, Z => n17560);
   U13229 : BUF_X1 port map( A => n15366, Z => n17548);
   U13230 : BUF_X1 port map( A => n15371, Z => n17536);
   U13231 : BUF_X1 port map( A => n15376, Z => n17524);
   U13232 : BUF_X1 port map( A => n14684, Z => n17709);
   U13233 : BUF_X1 port map( A => n14689, Z => n17697);
   U13234 : BUF_X1 port map( A => n14694, Z => n17685);
   U13235 : BUF_X1 port map( A => n14699, Z => n17673);
   U13236 : BUF_X1 port map( A => n14708, Z => n17661);
   U13237 : BUF_X1 port map( A => n14713, Z => n17649);
   U13238 : BUF_X1 port map( A => n14718, Z => n17637);
   U13239 : BUF_X1 port map( A => n14723, Z => n17625);
   U13240 : BUF_X1 port map( A => n14684, Z => n17710);
   U13241 : BUF_X1 port map( A => n14689, Z => n17698);
   U13242 : BUF_X1 port map( A => n14694, Z => n17686);
   U13243 : BUF_X1 port map( A => n14699, Z => n17674);
   U13244 : BUF_X1 port map( A => n14708, Z => n17662);
   U13245 : BUF_X1 port map( A => n14713, Z => n17650);
   U13246 : BUF_X1 port map( A => n14718, Z => n17638);
   U13247 : BUF_X1 port map( A => n14723, Z => n17626);
   U13248 : BUF_X1 port map( A => n15339, Z => n17606);
   U13249 : BUF_X1 port map( A => n15344, Z => n17594);
   U13250 : BUF_X1 port map( A => n15349, Z => n17582);
   U13251 : BUF_X1 port map( A => n15354, Z => n17570);
   U13252 : BUF_X1 port map( A => n15363, Z => n17558);
   U13253 : BUF_X1 port map( A => n15368, Z => n17546);
   U13254 : BUF_X1 port map( A => n15373, Z => n17534);
   U13255 : BUF_X1 port map( A => n15378, Z => n17522);
   U13256 : BUF_X1 port map( A => n14686, Z => n17708);
   U13257 : BUF_X1 port map( A => n14691, Z => n17696);
   U13258 : BUF_X1 port map( A => n14696, Z => n17684);
   U13259 : BUF_X1 port map( A => n14701, Z => n17672);
   U13260 : BUF_X1 port map( A => n14710, Z => n17660);
   U13261 : BUF_X1 port map( A => n14715, Z => n17648);
   U13262 : BUF_X1 port map( A => n14720, Z => n17636);
   U13263 : BUF_X1 port map( A => n14725, Z => n17624);
   U13264 : BUF_X1 port map( A => n15340, Z => n17603);
   U13265 : BUF_X1 port map( A => n15345, Z => n17591);
   U13266 : BUF_X1 port map( A => n15350, Z => n17579);
   U13267 : BUF_X1 port map( A => n15355, Z => n17567);
   U13268 : BUF_X1 port map( A => n15364, Z => n17555);
   U13269 : BUF_X1 port map( A => n15369, Z => n17543);
   U13270 : BUF_X1 port map( A => n15374, Z => n17531);
   U13271 : BUF_X1 port map( A => n15379, Z => n17519);
   U13272 : BUF_X1 port map( A => n14687, Z => n17705);
   U13273 : BUF_X1 port map( A => n14692, Z => n17693);
   U13274 : BUF_X1 port map( A => n14697, Z => n17681);
   U13275 : BUF_X1 port map( A => n14702, Z => n17669);
   U13276 : BUF_X1 port map( A => n14711, Z => n17657);
   U13277 : BUF_X1 port map( A => n14716, Z => n17645);
   U13278 : BUF_X1 port map( A => n14721, Z => n17633);
   U13279 : BUF_X1 port map( A => n14726, Z => n17621);
   U13280 : BUF_X1 port map( A => n15336, Z => n17612);
   U13281 : BUF_X1 port map( A => n15341, Z => n17600);
   U13282 : BUF_X1 port map( A => n15346, Z => n17588);
   U13283 : BUF_X1 port map( A => n15351, Z => n17576);
   U13284 : BUF_X1 port map( A => n15360, Z => n17564);
   U13285 : BUF_X1 port map( A => n15365, Z => n17552);
   U13286 : BUF_X1 port map( A => n15370, Z => n17540);
   U13287 : BUF_X1 port map( A => n15375, Z => n17528);
   U13288 : BUF_X1 port map( A => n14683, Z => n17714);
   U13289 : BUF_X1 port map( A => n14688, Z => n17702);
   U13290 : BUF_X1 port map( A => n14693, Z => n17690);
   U13291 : BUF_X1 port map( A => n14698, Z => n17678);
   U13292 : BUF_X1 port map( A => n14707, Z => n17666);
   U13293 : BUF_X1 port map( A => n14712, Z => n17654);
   U13294 : BUF_X1 port map( A => n14717, Z => n17642);
   U13295 : BUF_X1 port map( A => n14722, Z => n17630);
   U13296 : BUF_X1 port map( A => n15337, Z => n17609);
   U13297 : BUF_X1 port map( A => n15342, Z => n17597);
   U13298 : BUF_X1 port map( A => n15347, Z => n17585);
   U13299 : BUF_X1 port map( A => n15352, Z => n17573);
   U13300 : BUF_X1 port map( A => n15361, Z => n17561);
   U13301 : BUF_X1 port map( A => n15366, Z => n17549);
   U13302 : BUF_X1 port map( A => n15371, Z => n17537);
   U13303 : BUF_X1 port map( A => n15376, Z => n17525);
   U13304 : BUF_X1 port map( A => n14684, Z => n17711);
   U13305 : BUF_X1 port map( A => n14689, Z => n17699);
   U13306 : BUF_X1 port map( A => n14694, Z => n17687);
   U13307 : BUF_X1 port map( A => n14699, Z => n17675);
   U13308 : BUF_X1 port map( A => n14708, Z => n17663);
   U13309 : BUF_X1 port map( A => n14713, Z => n17651);
   U13310 : BUF_X1 port map( A => n14718, Z => n17639);
   U13311 : BUF_X1 port map( A => n14723, Z => n17627);
   U13312 : BUF_X1 port map( A => n17838, Z => n17831);
   U13313 : BUF_X1 port map( A => n17838, Z => n17832);
   U13314 : BUF_X1 port map( A => n17838, Z => n17833);
   U13315 : BUF_X1 port map( A => n17838, Z => n17834);
   U13316 : BUF_X1 port map( A => n17838, Z => n17835);
   U13317 : BUF_X1 port map( A => n17838, Z => n17836);
   U13318 : BUF_X1 port map( A => n17847, Z => n17840);
   U13319 : BUF_X1 port map( A => n17847, Z => n17841);
   U13320 : BUF_X1 port map( A => n17847, Z => n17842);
   U13321 : BUF_X1 port map( A => n17847, Z => n17843);
   U13322 : BUF_X1 port map( A => n17847, Z => n17844);
   U13323 : BUF_X1 port map( A => n17847, Z => n17845);
   U13324 : BUF_X1 port map( A => n17910, Z => n17903);
   U13325 : BUF_X1 port map( A => n17910, Z => n17904);
   U13326 : BUF_X1 port map( A => n17910, Z => n17905);
   U13327 : BUF_X1 port map( A => n17910, Z => n17906);
   U13328 : BUF_X1 port map( A => n17874, Z => n17867);
   U13329 : BUF_X1 port map( A => n17874, Z => n17868);
   U13330 : BUF_X1 port map( A => n17874, Z => n17869);
   U13331 : BUF_X1 port map( A => n17874, Z => n17870);
   U13332 : BUF_X1 port map( A => n17802, Z => n17795);
   U13333 : BUF_X1 port map( A => n17802, Z => n17796);
   U13334 : BUF_X1 port map( A => n17802, Z => n17797);
   U13335 : BUF_X1 port map( A => n17802, Z => n17798);
   U13336 : BUF_X1 port map( A => n17784, Z => n17777);
   U13337 : BUF_X1 port map( A => n17784, Z => n17778);
   U13338 : BUF_X1 port map( A => n17784, Z => n17779);
   U13339 : BUF_X1 port map( A => n17784, Z => n17780);
   U13340 : BUF_X1 port map( A => n17748, Z => n17741);
   U13341 : BUF_X1 port map( A => n17748, Z => n17742);
   U13342 : BUF_X1 port map( A => n17748, Z => n17743);
   U13343 : BUF_X1 port map( A => n17748, Z => n17744);
   U13344 : BUF_X1 port map( A => n17919, Z => n17912);
   U13345 : BUF_X1 port map( A => n17919, Z => n17913);
   U13346 : BUF_X1 port map( A => n17919, Z => n17914);
   U13347 : BUF_X1 port map( A => n17919, Z => n17915);
   U13348 : BUF_X1 port map( A => n17883, Z => n17876);
   U13349 : BUF_X1 port map( A => n17883, Z => n17877);
   U13350 : BUF_X1 port map( A => n17883, Z => n17878);
   U13351 : BUF_X1 port map( A => n17883, Z => n17879);
   U13352 : BUF_X1 port map( A => n17811, Z => n17804);
   U13353 : BUF_X1 port map( A => n17811, Z => n17805);
   U13354 : BUF_X1 port map( A => n17811, Z => n17806);
   U13355 : BUF_X1 port map( A => n17811, Z => n17807);
   U13356 : BUF_X1 port map( A => n17793, Z => n17786);
   U13357 : BUF_X1 port map( A => n17793, Z => n17787);
   U13358 : BUF_X1 port map( A => n17793, Z => n17788);
   U13359 : BUF_X1 port map( A => n17793, Z => n17789);
   U13360 : BUF_X1 port map( A => n17757, Z => n17750);
   U13361 : BUF_X1 port map( A => n17757, Z => n17751);
   U13362 : BUF_X1 port map( A => n17757, Z => n17752);
   U13363 : BUF_X1 port map( A => n17757, Z => n17753);
   U13364 : BUF_X1 port map( A => n17910, Z => n17907);
   U13365 : BUF_X1 port map( A => n17910, Z => n17908);
   U13366 : BUF_X1 port map( A => n17874, Z => n17871);
   U13367 : BUF_X1 port map( A => n17874, Z => n17872);
   U13368 : BUF_X1 port map( A => n17802, Z => n17799);
   U13369 : BUF_X1 port map( A => n17802, Z => n17800);
   U13370 : BUF_X1 port map( A => n17784, Z => n17781);
   U13371 : BUF_X1 port map( A => n17784, Z => n17782);
   U13372 : BUF_X1 port map( A => n17748, Z => n17745);
   U13373 : BUF_X1 port map( A => n17748, Z => n17746);
   U13374 : BUF_X1 port map( A => n17919, Z => n17916);
   U13375 : BUF_X1 port map( A => n17919, Z => n17917);
   U13376 : BUF_X1 port map( A => n17883, Z => n17880);
   U13377 : BUF_X1 port map( A => n17883, Z => n17881);
   U13378 : BUF_X1 port map( A => n17811, Z => n17808);
   U13379 : BUF_X1 port map( A => n17811, Z => n17809);
   U13380 : BUF_X1 port map( A => n17793, Z => n17790);
   U13381 : BUF_X1 port map( A => n17793, Z => n17791);
   U13382 : BUF_X1 port map( A => n17757, Z => n17754);
   U13383 : BUF_X1 port map( A => n17757, Z => n17755);
   U13384 : BUF_X1 port map( A => n17937, Z => n17930);
   U13385 : BUF_X1 port map( A => n17937, Z => n17931);
   U13386 : BUF_X1 port map( A => n17937, Z => n17932);
   U13387 : BUF_X1 port map( A => n17937, Z => n17933);
   U13388 : BUF_X1 port map( A => n17928, Z => n17921);
   U13389 : BUF_X1 port map( A => n17928, Z => n17922);
   U13390 : BUF_X1 port map( A => n17928, Z => n17923);
   U13391 : BUF_X1 port map( A => n17928, Z => n17924);
   U13392 : BUF_X1 port map( A => n17901, Z => n17894);
   U13393 : BUF_X1 port map( A => n17901, Z => n17895);
   U13394 : BUF_X1 port map( A => n17901, Z => n17896);
   U13395 : BUF_X1 port map( A => n17901, Z => n17897);
   U13396 : BUF_X1 port map( A => n17892, Z => n17885);
   U13397 : BUF_X1 port map( A => n17892, Z => n17886);
   U13398 : BUF_X1 port map( A => n17892, Z => n17887);
   U13399 : BUF_X1 port map( A => n17892, Z => n17888);
   U13400 : BUF_X1 port map( A => n17829, Z => n17822);
   U13401 : BUF_X1 port map( A => n17829, Z => n17823);
   U13402 : BUF_X1 port map( A => n17829, Z => n17824);
   U13403 : BUF_X1 port map( A => n17829, Z => n17825);
   U13404 : BUF_X1 port map( A => n17820, Z => n17813);
   U13405 : BUF_X1 port map( A => n17820, Z => n17814);
   U13406 : BUF_X1 port map( A => n17820, Z => n17815);
   U13407 : BUF_X1 port map( A => n17820, Z => n17816);
   U13408 : BUF_X1 port map( A => n17775, Z => n17768);
   U13409 : BUF_X1 port map( A => n17775, Z => n17769);
   U13410 : BUF_X1 port map( A => n17775, Z => n17770);
   U13411 : BUF_X1 port map( A => n17775, Z => n17771);
   U13412 : BUF_X1 port map( A => n17766, Z => n17759);
   U13413 : BUF_X1 port map( A => n17766, Z => n17760);
   U13414 : BUF_X1 port map( A => n17766, Z => n17761);
   U13415 : BUF_X1 port map( A => n17766, Z => n17762);
   U13416 : BUF_X1 port map( A => n17739, Z => n17732);
   U13417 : BUF_X1 port map( A => n17739, Z => n17733);
   U13418 : BUF_X1 port map( A => n17739, Z => n17734);
   U13419 : BUF_X1 port map( A => n17739, Z => n17735);
   U13420 : BUF_X1 port map( A => n17937, Z => n17934);
   U13421 : BUF_X1 port map( A => n17937, Z => n17935);
   U13422 : BUF_X1 port map( A => n17928, Z => n17925);
   U13423 : BUF_X1 port map( A => n17928, Z => n17926);
   U13424 : BUF_X1 port map( A => n17901, Z => n17898);
   U13425 : BUF_X1 port map( A => n17901, Z => n17899);
   U13426 : BUF_X1 port map( A => n17892, Z => n17889);
   U13427 : BUF_X1 port map( A => n17892, Z => n17890);
   U13428 : BUF_X1 port map( A => n17829, Z => n17826);
   U13429 : BUF_X1 port map( A => n17829, Z => n17827);
   U13430 : BUF_X1 port map( A => n17820, Z => n17817);
   U13431 : BUF_X1 port map( A => n17820, Z => n17818);
   U13432 : BUF_X1 port map( A => n17775, Z => n17772);
   U13433 : BUF_X1 port map( A => n17775, Z => n17773);
   U13434 : BUF_X1 port map( A => n17766, Z => n17763);
   U13435 : BUF_X1 port map( A => n17766, Z => n17764);
   U13436 : BUF_X1 port map( A => n17739, Z => n17736);
   U13437 : BUF_X1 port map( A => n17739, Z => n17737);
   U13438 : BUF_X1 port map( A => n17865, Z => n17858);
   U13439 : BUF_X1 port map( A => n17865, Z => n17859);
   U13440 : BUF_X1 port map( A => n17865, Z => n17860);
   U13441 : BUF_X1 port map( A => n17865, Z => n17861);
   U13442 : BUF_X1 port map( A => n17856, Z => n17849);
   U13443 : BUF_X1 port map( A => n17856, Z => n17850);
   U13444 : BUF_X1 port map( A => n17856, Z => n17851);
   U13445 : BUF_X1 port map( A => n17856, Z => n17852);
   U13446 : BUF_X1 port map( A => n17865, Z => n17862);
   U13447 : BUF_X1 port map( A => n17865, Z => n17863);
   U13448 : BUF_X1 port map( A => n17856, Z => n17853);
   U13449 : BUF_X1 port map( A => n17856, Z => n17854);
   U13450 : BUF_X1 port map( A => n17946, Z => n17939);
   U13451 : BUF_X1 port map( A => n17946, Z => n17940);
   U13452 : BUF_X1 port map( A => n17946, Z => n17941);
   U13453 : BUF_X1 port map( A => n17946, Z => n17942);
   U13454 : BUF_X1 port map( A => n18000, Z => n17993);
   U13455 : BUF_X1 port map( A => n18000, Z => n17994);
   U13456 : BUF_X1 port map( A => n18000, Z => n17995);
   U13457 : BUF_X1 port map( A => n18000, Z => n17996);
   U13458 : BUF_X1 port map( A => n17955, Z => n17948);
   U13459 : BUF_X1 port map( A => n17955, Z => n17949);
   U13460 : BUF_X1 port map( A => n17955, Z => n17950);
   U13461 : BUF_X1 port map( A => n17955, Z => n17951);
   U13462 : BUF_X1 port map( A => n17946, Z => n17943);
   U13463 : BUF_X1 port map( A => n17946, Z => n17944);
   U13464 : BUF_X1 port map( A => n18000, Z => n17997);
   U13465 : BUF_X1 port map( A => n18000, Z => n17998);
   U13466 : BUF_X1 port map( A => n17955, Z => n17952);
   U13467 : BUF_X1 port map( A => n17955, Z => n17953);
   U13468 : BUF_X1 port map( A => n17991, Z => n17984);
   U13469 : BUF_X1 port map( A => n17991, Z => n17985);
   U13470 : BUF_X1 port map( A => n17991, Z => n17986);
   U13471 : BUF_X1 port map( A => n17991, Z => n17987);
   U13472 : BUF_X1 port map( A => n17982, Z => n17975);
   U13473 : BUF_X1 port map( A => n17982, Z => n17976);
   U13474 : BUF_X1 port map( A => n17982, Z => n17977);
   U13475 : BUF_X1 port map( A => n17982, Z => n17978);
   U13476 : BUF_X1 port map( A => n17973, Z => n17966);
   U13477 : BUF_X1 port map( A => n17973, Z => n17967);
   U13478 : BUF_X1 port map( A => n17973, Z => n17968);
   U13479 : BUF_X1 port map( A => n17973, Z => n17969);
   U13480 : BUF_X1 port map( A => n17964, Z => n17957);
   U13481 : BUF_X1 port map( A => n17964, Z => n17958);
   U13482 : BUF_X1 port map( A => n17964, Z => n17959);
   U13483 : BUF_X1 port map( A => n17964, Z => n17960);
   U13484 : BUF_X1 port map( A => n17991, Z => n17988);
   U13485 : BUF_X1 port map( A => n17991, Z => n17989);
   U13486 : BUF_X1 port map( A => n17982, Z => n17979);
   U13487 : BUF_X1 port map( A => n17982, Z => n17980);
   U13488 : BUF_X1 port map( A => n17973, Z => n17970);
   U13489 : BUF_X1 port map( A => n17973, Z => n17971);
   U13490 : BUF_X1 port map( A => n17964, Z => n17961);
   U13491 : BUF_X1 port map( A => n17964, Z => n17962);
   U13492 : BUF_X1 port map( A => n17838, Z => n17837);
   U13493 : BUF_X1 port map( A => n17847, Z => n17846);
   U13494 : BUF_X1 port map( A => n17910, Z => n17909);
   U13495 : BUF_X1 port map( A => n17874, Z => n17873);
   U13496 : BUF_X1 port map( A => n17802, Z => n17801);
   U13497 : BUF_X1 port map( A => n17784, Z => n17783);
   U13498 : BUF_X1 port map( A => n17748, Z => n17747);
   U13499 : BUF_X1 port map( A => n17919, Z => n17918);
   U13500 : BUF_X1 port map( A => n17883, Z => n17882);
   U13501 : BUF_X1 port map( A => n17811, Z => n17810);
   U13502 : BUF_X1 port map( A => n17793, Z => n17792);
   U13503 : BUF_X1 port map( A => n17757, Z => n17756);
   U13504 : BUF_X1 port map( A => n17937, Z => n17936);
   U13505 : BUF_X1 port map( A => n17928, Z => n17927);
   U13506 : BUF_X1 port map( A => n17901, Z => n17900);
   U13507 : BUF_X1 port map( A => n17892, Z => n17891);
   U13508 : BUF_X1 port map( A => n17829, Z => n17828);
   U13509 : BUF_X1 port map( A => n17820, Z => n17819);
   U13510 : BUF_X1 port map( A => n17775, Z => n17774);
   U13511 : BUF_X1 port map( A => n17766, Z => n17765);
   U13512 : BUF_X1 port map( A => n17739, Z => n17738);
   U13513 : BUF_X1 port map( A => n17865, Z => n17864);
   U13514 : BUF_X1 port map( A => n17856, Z => n17855);
   U13515 : BUF_X1 port map( A => n17946, Z => n17945);
   U13516 : BUF_X1 port map( A => n18000, Z => n17999);
   U13517 : BUF_X1 port map( A => n17955, Z => n17954);
   U13518 : BUF_X1 port map( A => n17991, Z => n17990);
   U13519 : BUF_X1 port map( A => n17982, Z => n17981);
   U13520 : BUF_X1 port map( A => n17973, Z => n17972);
   U13521 : BUF_X1 port map( A => n17964, Z => n17963);
   U13522 : INV_X1 port map( A => n14598, ZN => n18105);
   U13523 : OAI21_X1 port map( B1 => n14630, B2 => n14631, A => n18003, ZN => 
                           n14598);
   U13524 : INV_X1 port map( A => n17721, ZN => n17730);
   U13525 : AOI221_X1 port map( B1 => n17562, B2 => n17277, C1 => n17559, C2 =>
                           n16813, A => n15973, ZN => n15972);
   U13526 : OAI22_X1 port map( A1 => n16653, A2 => n17556, B1 => n17053, B2 => 
                           n17553, ZN => n15973);
   U13527 : AOI221_X1 port map( B1 => n17562, B2 => n17278, C1 => n17559, C2 =>
                           n16814, A => n15946, ZN => n15945);
   U13528 : OAI22_X1 port map( A1 => n16654, A2 => n17556, B1 => n17054, B2 => 
                           n17553, ZN => n15946);
   U13529 : AOI221_X1 port map( B1 => n17562, B2 => n17279, C1 => n17559, C2 =>
                           n16815, A => n15927, ZN => n15926);
   U13530 : OAI22_X1 port map( A1 => n16655, A2 => n17556, B1 => n17055, B2 => 
                           n17553, ZN => n15927);
   U13531 : AOI221_X1 port map( B1 => n17562, B2 => n17280, C1 => n17559, C2 =>
                           n16816, A => n15908, ZN => n15907);
   U13532 : OAI22_X1 port map( A1 => n16656, A2 => n17556, B1 => n17056, B2 => 
                           n17553, ZN => n15908);
   U13533 : AOI221_X1 port map( B1 => n17562, B2 => n17281, C1 => n17559, C2 =>
                           n16817, A => n15889, ZN => n15888);
   U13534 : OAI22_X1 port map( A1 => n16657, A2 => n17556, B1 => n17057, B2 => 
                           n17553, ZN => n15889);
   U13535 : AOI221_X1 port map( B1 => n17562, B2 => n17282, C1 => n17559, C2 =>
                           n16818, A => n15870, ZN => n15869);
   U13536 : OAI22_X1 port map( A1 => n16658, A2 => n17556, B1 => n17058, B2 => 
                           n17553, ZN => n15870);
   U13537 : AOI221_X1 port map( B1 => n17562, B2 => n17283, C1 => n17559, C2 =>
                           n16819, A => n15851, ZN => n15850);
   U13538 : OAI22_X1 port map( A1 => n16659, A2 => n17556, B1 => n17059, B2 => 
                           n17553, ZN => n15851);
   U13539 : AOI221_X1 port map( B1 => n17562, B2 => n17284, C1 => n17559, C2 =>
                           n16820, A => n15832, ZN => n15831);
   U13540 : OAI22_X1 port map( A1 => n16660, A2 => n17556, B1 => n17060, B2 => 
                           n17553, ZN => n15832);
   U13541 : AOI221_X1 port map( B1 => n17562, B2 => n17285, C1 => n17559, C2 =>
                           n16821, A => n15813, ZN => n15812);
   U13542 : OAI22_X1 port map( A1 => n16661, A2 => n17556, B1 => n17061, B2 => 
                           n17553, ZN => n15813);
   U13543 : AOI221_X1 port map( B1 => n17562, B2 => n17286, C1 => n17559, C2 =>
                           n16822, A => n15794, ZN => n15793);
   U13544 : OAI22_X1 port map( A1 => n16662, A2 => n17556, B1 => n17062, B2 => 
                           n17553, ZN => n15794);
   U13545 : AOI221_X1 port map( B1 => n17562, B2 => n17287, C1 => n17559, C2 =>
                           n16823, A => n15775, ZN => n15774);
   U13546 : OAI22_X1 port map( A1 => n16663, A2 => n17556, B1 => n17063, B2 => 
                           n17553, ZN => n15775);
   U13547 : AOI221_X1 port map( B1 => n17562, B2 => n17288, C1 => n17559, C2 =>
                           n16824, A => n15756, ZN => n15755);
   U13548 : OAI22_X1 port map( A1 => n16664, A2 => n17556, B1 => n17064, B2 => 
                           n17553, ZN => n15756);
   U13549 : AOI221_X1 port map( B1 => n17563, B2 => n17289, C1 => n17560, C2 =>
                           n16825, A => n15737, ZN => n15736);
   U13550 : OAI22_X1 port map( A1 => n16549, A2 => n17557, B1 => n17065, B2 => 
                           n17554, ZN => n15737);
   U13551 : AOI221_X1 port map( B1 => n17563, B2 => n17290, C1 => n17560, C2 =>
                           n16826, A => n15718, ZN => n15717);
   U13552 : OAI22_X1 port map( A1 => n16550, A2 => n17557, B1 => n17066, B2 => 
                           n17554, ZN => n15718);
   U13553 : AOI221_X1 port map( B1 => n17563, B2 => n17291, C1 => n17560, C2 =>
                           n16827, A => n15699, ZN => n15698);
   U13554 : OAI22_X1 port map( A1 => n16551, A2 => n17557, B1 => n17067, B2 => 
                           n17554, ZN => n15699);
   U13555 : AOI221_X1 port map( B1 => n17563, B2 => n17292, C1 => n17560, C2 =>
                           n16828, A => n15680, ZN => n15679);
   U13556 : OAI22_X1 port map( A1 => n16552, A2 => n17557, B1 => n17068, B2 => 
                           n17554, ZN => n15680);
   U13557 : AOI221_X1 port map( B1 => n17563, B2 => n17293, C1 => n17560, C2 =>
                           n16829, A => n15661, ZN => n15660);
   U13558 : OAI22_X1 port map( A1 => n16553, A2 => n17557, B1 => n17069, B2 => 
                           n17554, ZN => n15661);
   U13559 : AOI221_X1 port map( B1 => n17563, B2 => n17294, C1 => n17560, C2 =>
                           n16830, A => n15642, ZN => n15641);
   U13560 : OAI22_X1 port map( A1 => n16554, A2 => n17557, B1 => n17070, B2 => 
                           n17554, ZN => n15642);
   U13561 : AOI221_X1 port map( B1 => n17563, B2 => n17295, C1 => n17560, C2 =>
                           n16831, A => n15623, ZN => n15622);
   U13562 : OAI22_X1 port map( A1 => n16555, A2 => n17557, B1 => n17071, B2 => 
                           n17554, ZN => n15623);
   U13563 : AOI221_X1 port map( B1 => n17563, B2 => n17296, C1 => n17560, C2 =>
                           n16832, A => n15604, ZN => n15603);
   U13564 : OAI22_X1 port map( A1 => n16556, A2 => n17557, B1 => n17072, B2 => 
                           n17554, ZN => n15604);
   U13565 : AOI221_X1 port map( B1 => n17563, B2 => n17297, C1 => n17560, C2 =>
                           n16833, A => n15585, ZN => n15584);
   U13566 : OAI22_X1 port map( A1 => n16557, A2 => n17557, B1 => n17073, B2 => 
                           n17554, ZN => n15585);
   U13567 : AOI221_X1 port map( B1 => n17563, B2 => n17298, C1 => n17560, C2 =>
                           n16834, A => n15566, ZN => n15565);
   U13568 : OAI22_X1 port map( A1 => n16558, A2 => n17557, B1 => n17074, B2 => 
                           n17554, ZN => n15566);
   U13569 : AOI221_X1 port map( B1 => n17563, B2 => n17299, C1 => n17560, C2 =>
                           n16835, A => n15547, ZN => n15546);
   U13570 : OAI22_X1 port map( A1 => n16559, A2 => n17557, B1 => n17075, B2 => 
                           n17554, ZN => n15547);
   U13571 : AOI221_X1 port map( B1 => n17563, B2 => n17300, C1 => n17560, C2 =>
                           n16836, A => n15528, ZN => n15527);
   U13572 : OAI22_X1 port map( A1 => n16560, A2 => n17557, B1 => n17076, B2 => 
                           n17554, ZN => n15528);
   U13573 : AOI221_X1 port map( B1 => n17564, B2 => n17301, C1 => n17561, C2 =>
                           n16837, A => n15509, ZN => n15508);
   U13574 : OAI22_X1 port map( A1 => n16493, A2 => n17558, B1 => n16749, B2 => 
                           n17555, ZN => n15509);
   U13575 : AOI221_X1 port map( B1 => n17564, B2 => n17302, C1 => n17561, C2 =>
                           n16838, A => n15490, ZN => n15489);
   U13576 : OAI22_X1 port map( A1 => n16494, A2 => n17558, B1 => n16750, B2 => 
                           n17555, ZN => n15490);
   U13577 : AOI221_X1 port map( B1 => n17564, B2 => n17303, C1 => n17561, C2 =>
                           n16839, A => n15471, ZN => n15470);
   U13578 : OAI22_X1 port map( A1 => n16495, A2 => n17558, B1 => n16751, B2 => 
                           n17555, ZN => n15471);
   U13579 : AOI221_X1 port map( B1 => n17564, B2 => n17304, C1 => n17561, C2 =>
                           n16840, A => n15452, ZN => n15451);
   U13580 : OAI22_X1 port map( A1 => n16496, A2 => n17558, B1 => n16752, B2 => 
                           n17555, ZN => n15452);
   U13581 : AOI221_X1 port map( B1 => n17564, B2 => n17305, C1 => n17561, C2 =>
                           n16841, A => n15433, ZN => n15432);
   U13582 : OAI22_X1 port map( A1 => n16497, A2 => n17558, B1 => n16753, B2 => 
                           n17555, ZN => n15433);
   U13583 : AOI221_X1 port map( B1 => n17564, B2 => n17306, C1 => n17561, C2 =>
                           n16842, A => n15414, ZN => n15413);
   U13584 : OAI22_X1 port map( A1 => n16498, A2 => n17558, B1 => n16754, B2 => 
                           n17555, ZN => n15414);
   U13585 : AOI221_X1 port map( B1 => n17564, B2 => n17307, C1 => n17561, C2 =>
                           n16843, A => n15395, ZN => n15394);
   U13586 : OAI22_X1 port map( A1 => n16499, A2 => n17558, B1 => n16755, B2 => 
                           n17555, ZN => n15395);
   U13587 : AOI221_X1 port map( B1 => n17564, B2 => n17308, C1 => n17561, C2 =>
                           n16844, A => n15362, ZN => n15359);
   U13588 : OAI22_X1 port map( A1 => n16500, A2 => n17558, B1 => n16756, B2 => 
                           n17555, ZN => n15362);
   U13589 : AOI221_X1 port map( B1 => n17664, B2 => n17277, C1 => n17661, C2 =>
                           n16813, A => n15320, ZN => n15319);
   U13590 : OAI22_X1 port map( A1 => n16653, A2 => n17658, B1 => n17053, B2 => 
                           n17655, ZN => n15320);
   U13591 : AOI221_X1 port map( B1 => n17664, B2 => n17278, C1 => n17661, C2 =>
                           n16814, A => n15293, ZN => n15292);
   U13592 : OAI22_X1 port map( A1 => n16654, A2 => n17658, B1 => n17054, B2 => 
                           n17655, ZN => n15293);
   U13593 : AOI221_X1 port map( B1 => n17664, B2 => n17279, C1 => n17661, C2 =>
                           n16815, A => n15274, ZN => n15273);
   U13594 : OAI22_X1 port map( A1 => n16655, A2 => n17658, B1 => n17055, B2 => 
                           n17655, ZN => n15274);
   U13595 : AOI221_X1 port map( B1 => n17664, B2 => n17280, C1 => n17661, C2 =>
                           n16816, A => n15255, ZN => n15254);
   U13596 : OAI22_X1 port map( A1 => n16656, A2 => n17658, B1 => n17056, B2 => 
                           n17655, ZN => n15255);
   U13597 : AOI221_X1 port map( B1 => n17664, B2 => n17281, C1 => n17661, C2 =>
                           n16817, A => n15236, ZN => n15235);
   U13598 : OAI22_X1 port map( A1 => n16657, A2 => n17658, B1 => n17057, B2 => 
                           n17655, ZN => n15236);
   U13599 : AOI221_X1 port map( B1 => n17664, B2 => n17282, C1 => n17661, C2 =>
                           n16818, A => n15217, ZN => n15216);
   U13600 : OAI22_X1 port map( A1 => n16658, A2 => n17658, B1 => n17058, B2 => 
                           n17655, ZN => n15217);
   U13601 : AOI221_X1 port map( B1 => n17664, B2 => n17283, C1 => n17661, C2 =>
                           n16819, A => n15198, ZN => n15197);
   U13602 : OAI22_X1 port map( A1 => n16659, A2 => n17658, B1 => n17059, B2 => 
                           n17655, ZN => n15198);
   U13603 : AOI221_X1 port map( B1 => n17664, B2 => n17284, C1 => n17661, C2 =>
                           n16820, A => n15179, ZN => n15178);
   U13604 : OAI22_X1 port map( A1 => n16660, A2 => n17658, B1 => n17060, B2 => 
                           n17655, ZN => n15179);
   U13605 : AOI221_X1 port map( B1 => n17664, B2 => n17285, C1 => n17661, C2 =>
                           n16821, A => n15160, ZN => n15159);
   U13606 : OAI22_X1 port map( A1 => n16661, A2 => n17658, B1 => n17061, B2 => 
                           n17655, ZN => n15160);
   U13607 : AOI221_X1 port map( B1 => n17664, B2 => n17286, C1 => n17661, C2 =>
                           n16822, A => n15141, ZN => n15140);
   U13608 : OAI22_X1 port map( A1 => n16662, A2 => n17658, B1 => n17062, B2 => 
                           n17655, ZN => n15141);
   U13609 : AOI221_X1 port map( B1 => n17664, B2 => n17287, C1 => n17661, C2 =>
                           n16823, A => n15122, ZN => n15121);
   U13610 : OAI22_X1 port map( A1 => n16663, A2 => n17658, B1 => n17063, B2 => 
                           n17655, ZN => n15122);
   U13611 : AOI221_X1 port map( B1 => n17664, B2 => n17288, C1 => n17661, C2 =>
                           n16824, A => n15103, ZN => n15102);
   U13612 : OAI22_X1 port map( A1 => n16664, A2 => n17658, B1 => n17064, B2 => 
                           n17655, ZN => n15103);
   U13613 : AOI221_X1 port map( B1 => n17665, B2 => n17289, C1 => n17662, C2 =>
                           n16825, A => n15084, ZN => n15083);
   U13614 : OAI22_X1 port map( A1 => n16549, A2 => n17659, B1 => n17065, B2 => 
                           n17656, ZN => n15084);
   U13615 : AOI221_X1 port map( B1 => n17665, B2 => n17290, C1 => n17662, C2 =>
                           n16826, A => n15065, ZN => n15064);
   U13616 : OAI22_X1 port map( A1 => n16550, A2 => n17659, B1 => n17066, B2 => 
                           n17656, ZN => n15065);
   U13617 : AOI221_X1 port map( B1 => n17665, B2 => n17291, C1 => n17662, C2 =>
                           n16827, A => n15046, ZN => n15045);
   U13618 : OAI22_X1 port map( A1 => n16551, A2 => n17659, B1 => n17067, B2 => 
                           n17656, ZN => n15046);
   U13619 : AOI221_X1 port map( B1 => n17665, B2 => n17292, C1 => n17662, C2 =>
                           n16828, A => n15027, ZN => n15026);
   U13620 : OAI22_X1 port map( A1 => n16552, A2 => n17659, B1 => n17068, B2 => 
                           n17656, ZN => n15027);
   U13621 : AOI221_X1 port map( B1 => n17665, B2 => n17293, C1 => n17662, C2 =>
                           n16829, A => n15008, ZN => n15007);
   U13622 : OAI22_X1 port map( A1 => n16553, A2 => n17659, B1 => n17069, B2 => 
                           n17656, ZN => n15008);
   U13623 : AOI221_X1 port map( B1 => n17665, B2 => n17294, C1 => n17662, C2 =>
                           n16830, A => n14989, ZN => n14988);
   U13624 : OAI22_X1 port map( A1 => n16554, A2 => n17659, B1 => n17070, B2 => 
                           n17656, ZN => n14989);
   U13625 : AOI221_X1 port map( B1 => n17665, B2 => n17295, C1 => n17662, C2 =>
                           n16831, A => n14970, ZN => n14969);
   U13626 : OAI22_X1 port map( A1 => n16555, A2 => n17659, B1 => n17071, B2 => 
                           n17656, ZN => n14970);
   U13627 : AOI221_X1 port map( B1 => n17665, B2 => n17296, C1 => n17662, C2 =>
                           n16832, A => n14951, ZN => n14950);
   U13628 : OAI22_X1 port map( A1 => n16556, A2 => n17659, B1 => n17072, B2 => 
                           n17656, ZN => n14951);
   U13629 : AOI221_X1 port map( B1 => n17665, B2 => n17297, C1 => n17662, C2 =>
                           n16833, A => n14932, ZN => n14931);
   U13630 : OAI22_X1 port map( A1 => n16557, A2 => n17659, B1 => n17073, B2 => 
                           n17656, ZN => n14932);
   U13631 : AOI221_X1 port map( B1 => n17665, B2 => n17298, C1 => n17662, C2 =>
                           n16834, A => n14913, ZN => n14912);
   U13632 : OAI22_X1 port map( A1 => n16558, A2 => n17659, B1 => n17074, B2 => 
                           n17656, ZN => n14913);
   U13633 : AOI221_X1 port map( B1 => n17665, B2 => n17299, C1 => n17662, C2 =>
                           n16835, A => n14894, ZN => n14893);
   U13634 : OAI22_X1 port map( A1 => n16559, A2 => n17659, B1 => n17075, B2 => 
                           n17656, ZN => n14894);
   U13635 : AOI221_X1 port map( B1 => n17665, B2 => n17300, C1 => n17662, C2 =>
                           n16836, A => n14875, ZN => n14874);
   U13636 : OAI22_X1 port map( A1 => n16560, A2 => n17659, B1 => n17076, B2 => 
                           n17656, ZN => n14875);
   U13637 : AOI221_X1 port map( B1 => n17666, B2 => n17301, C1 => n17663, C2 =>
                           n16837, A => n14856, ZN => n14855);
   U13638 : OAI22_X1 port map( A1 => n16493, A2 => n17660, B1 => n16749, B2 => 
                           n17657, ZN => n14856);
   U13639 : AOI221_X1 port map( B1 => n17666, B2 => n17302, C1 => n17663, C2 =>
                           n16838, A => n14837, ZN => n14836);
   U13640 : OAI22_X1 port map( A1 => n16494, A2 => n17660, B1 => n16750, B2 => 
                           n17657, ZN => n14837);
   U13641 : AOI221_X1 port map( B1 => n17666, B2 => n17303, C1 => n17663, C2 =>
                           n16839, A => n14818, ZN => n14817);
   U13642 : OAI22_X1 port map( A1 => n16495, A2 => n17660, B1 => n16751, B2 => 
                           n17657, ZN => n14818);
   U13643 : AOI221_X1 port map( B1 => n17666, B2 => n17304, C1 => n17663, C2 =>
                           n16840, A => n14799, ZN => n14798);
   U13644 : OAI22_X1 port map( A1 => n16496, A2 => n17660, B1 => n16752, B2 => 
                           n17657, ZN => n14799);
   U13645 : AOI221_X1 port map( B1 => n17666, B2 => n17305, C1 => n17663, C2 =>
                           n16841, A => n14780, ZN => n14779);
   U13646 : OAI22_X1 port map( A1 => n16497, A2 => n17660, B1 => n16753, B2 => 
                           n17657, ZN => n14780);
   U13647 : AOI221_X1 port map( B1 => n17666, B2 => n17306, C1 => n17663, C2 =>
                           n16842, A => n14761, ZN => n14760);
   U13648 : OAI22_X1 port map( A1 => n16498, A2 => n17660, B1 => n16754, B2 => 
                           n17657, ZN => n14761);
   U13649 : AOI221_X1 port map( B1 => n17666, B2 => n17307, C1 => n17663, C2 =>
                           n16843, A => n14742, ZN => n14741);
   U13650 : OAI22_X1 port map( A1 => n16499, A2 => n17660, B1 => n16755, B2 => 
                           n17657, ZN => n14742);
   U13651 : AOI221_X1 port map( B1 => n17666, B2 => n17308, C1 => n17663, C2 =>
                           n16844, A => n14709, ZN => n14706);
   U13652 : OAI22_X1 port map( A1 => n16500, A2 => n17660, B1 => n16756, B2 => 
                           n17657, ZN => n14709);
   U13653 : AOI221_X1 port map( B1 => n17598, B2 => n17309, C1 => n17595, C2 =>
                           n16845, A => n15962, ZN => n15955);
   U13654 : OAI22_X1 port map( A1 => n16701, A2 => n17592, B1 => n17149, B2 => 
                           n17589, ZN => n15962);
   U13655 : AOI221_X1 port map( B1 => n17550, B2 => n17310, C1 => n17547, C2 =>
                           n16846, A => n15976, ZN => n15971);
   U13656 : OAI22_X1 port map( A1 => n16665, A2 => n17544, B1 => n17077, B2 => 
                           n17541, ZN => n15976);
   U13657 : AOI221_X1 port map( B1 => n17598, B2 => n17311, C1 => n17595, C2 =>
                           n16847, A => n15939, ZN => n15936);
   U13658 : OAI22_X1 port map( A1 => n16702, A2 => n17592, B1 => n17150, B2 => 
                           n17589, ZN => n15939);
   U13659 : AOI221_X1 port map( B1 => n17550, B2 => n17312, C1 => n17547, C2 =>
                           n16848, A => n15947, ZN => n15944);
   U13660 : OAI22_X1 port map( A1 => n16666, A2 => n17544, B1 => n17078, B2 => 
                           n17541, ZN => n15947);
   U13661 : AOI221_X1 port map( B1 => n17598, B2 => n17313, C1 => n17595, C2 =>
                           n16849, A => n15920, ZN => n15917);
   U13662 : OAI22_X1 port map( A1 => n16703, A2 => n17592, B1 => n17151, B2 => 
                           n17589, ZN => n15920);
   U13663 : AOI221_X1 port map( B1 => n17550, B2 => n17314, C1 => n17547, C2 =>
                           n16850, A => n15928, ZN => n15925);
   U13664 : OAI22_X1 port map( A1 => n16667, A2 => n17544, B1 => n17079, B2 => 
                           n17541, ZN => n15928);
   U13665 : AOI221_X1 port map( B1 => n17598, B2 => n17315, C1 => n17595, C2 =>
                           n16851, A => n15901, ZN => n15898);
   U13666 : OAI22_X1 port map( A1 => n16704, A2 => n17592, B1 => n17152, B2 => 
                           n17589, ZN => n15901);
   U13667 : AOI221_X1 port map( B1 => n17550, B2 => n17316, C1 => n17547, C2 =>
                           n16852, A => n15909, ZN => n15906);
   U13668 : OAI22_X1 port map( A1 => n16668, A2 => n17544, B1 => n17080, B2 => 
                           n17541, ZN => n15909);
   U13669 : AOI221_X1 port map( B1 => n17598, B2 => n17317, C1 => n17595, C2 =>
                           n16853, A => n15882, ZN => n15879);
   U13670 : OAI22_X1 port map( A1 => n16705, A2 => n17592, B1 => n17153, B2 => 
                           n17589, ZN => n15882);
   U13671 : AOI221_X1 port map( B1 => n17550, B2 => n17318, C1 => n17547, C2 =>
                           n16854, A => n15890, ZN => n15887);
   U13672 : OAI22_X1 port map( A1 => n16669, A2 => n17544, B1 => n17081, B2 => 
                           n17541, ZN => n15890);
   U13673 : AOI221_X1 port map( B1 => n17598, B2 => n17319, C1 => n17595, C2 =>
                           n16855, A => n15863, ZN => n15860);
   U13674 : OAI22_X1 port map( A1 => n16706, A2 => n17592, B1 => n17154, B2 => 
                           n17589, ZN => n15863);
   U13675 : AOI221_X1 port map( B1 => n17550, B2 => n17320, C1 => n17547, C2 =>
                           n16856, A => n15871, ZN => n15868);
   U13676 : OAI22_X1 port map( A1 => n16670, A2 => n17544, B1 => n17082, B2 => 
                           n17541, ZN => n15871);
   U13677 : AOI221_X1 port map( B1 => n17598, B2 => n17321, C1 => n17595, C2 =>
                           n16857, A => n15844, ZN => n15841);
   U13678 : OAI22_X1 port map( A1 => n16707, A2 => n17592, B1 => n17155, B2 => 
                           n17589, ZN => n15844);
   U13679 : AOI221_X1 port map( B1 => n17550, B2 => n17322, C1 => n17547, C2 =>
                           n16858, A => n15852, ZN => n15849);
   U13680 : OAI22_X1 port map( A1 => n16671, A2 => n17544, B1 => n17083, B2 => 
                           n17541, ZN => n15852);
   U13681 : AOI221_X1 port map( B1 => n17598, B2 => n17323, C1 => n17595, C2 =>
                           n16859, A => n15825, ZN => n15822);
   U13682 : OAI22_X1 port map( A1 => n16708, A2 => n17592, B1 => n17156, B2 => 
                           n17589, ZN => n15825);
   U13683 : AOI221_X1 port map( B1 => n17550, B2 => n17324, C1 => n17547, C2 =>
                           n16860, A => n15833, ZN => n15830);
   U13684 : OAI22_X1 port map( A1 => n16672, A2 => n17544, B1 => n17084, B2 => 
                           n17541, ZN => n15833);
   U13685 : AOI221_X1 port map( B1 => n17598, B2 => n17325, C1 => n17595, C2 =>
                           n16861, A => n15806, ZN => n15803);
   U13686 : OAI22_X1 port map( A1 => n16709, A2 => n17592, B1 => n17157, B2 => 
                           n17589, ZN => n15806);
   U13687 : AOI221_X1 port map( B1 => n17550, B2 => n17326, C1 => n17547, C2 =>
                           n16862, A => n15814, ZN => n15811);
   U13688 : OAI22_X1 port map( A1 => n16673, A2 => n17544, B1 => n17085, B2 => 
                           n17541, ZN => n15814);
   U13689 : AOI221_X1 port map( B1 => n17598, B2 => n17327, C1 => n17595, C2 =>
                           n16863, A => n15787, ZN => n15784);
   U13690 : OAI22_X1 port map( A1 => n16710, A2 => n17592, B1 => n17158, B2 => 
                           n17589, ZN => n15787);
   U13691 : AOI221_X1 port map( B1 => n17550, B2 => n17328, C1 => n17547, C2 =>
                           n16864, A => n15795, ZN => n15792);
   U13692 : OAI22_X1 port map( A1 => n16674, A2 => n17544, B1 => n17086, B2 => 
                           n17541, ZN => n15795);
   U13693 : AOI221_X1 port map( B1 => n17598, B2 => n17329, C1 => n17595, C2 =>
                           n16865, A => n15768, ZN => n15765);
   U13694 : OAI22_X1 port map( A1 => n16711, A2 => n17592, B1 => n17159, B2 => 
                           n17589, ZN => n15768);
   U13695 : AOI221_X1 port map( B1 => n17550, B2 => n17330, C1 => n17547, C2 =>
                           n16866, A => n15776, ZN => n15773);
   U13696 : OAI22_X1 port map( A1 => n16675, A2 => n17544, B1 => n17087, B2 => 
                           n17541, ZN => n15776);
   U13697 : AOI221_X1 port map( B1 => n17598, B2 => n17331, C1 => n17595, C2 =>
                           n16867, A => n15749, ZN => n15746);
   U13698 : OAI22_X1 port map( A1 => n16712, A2 => n17592, B1 => n17160, B2 => 
                           n17589, ZN => n15749);
   U13699 : AOI221_X1 port map( B1 => n17550, B2 => n17332, C1 => n17547, C2 =>
                           n16868, A => n15757, ZN => n15754);
   U13700 : OAI22_X1 port map( A1 => n16676, A2 => n17544, B1 => n17088, B2 => 
                           n17541, ZN => n15757);
   U13701 : AOI221_X1 port map( B1 => n17599, B2 => n17333, C1 => n17596, C2 =>
                           n16869, A => n15730, ZN => n15727);
   U13702 : OAI22_X1 port map( A1 => n16597, A2 => n17593, B1 => n17161, B2 => 
                           n17590, ZN => n15730);
   U13703 : AOI221_X1 port map( B1 => n17551, B2 => n17334, C1 => n17548, C2 =>
                           n16870, A => n15738, ZN => n15735);
   U13704 : OAI22_X1 port map( A1 => n16561, A2 => n17545, B1 => n17089, B2 => 
                           n17542, ZN => n15738);
   U13705 : AOI221_X1 port map( B1 => n17599, B2 => n17335, C1 => n17596, C2 =>
                           n16871, A => n15711, ZN => n15708);
   U13706 : OAI22_X1 port map( A1 => n16598, A2 => n17593, B1 => n17162, B2 => 
                           n17590, ZN => n15711);
   U13707 : AOI221_X1 port map( B1 => n17551, B2 => n17336, C1 => n17548, C2 =>
                           n16872, A => n15719, ZN => n15716);
   U13708 : OAI22_X1 port map( A1 => n16562, A2 => n17545, B1 => n17090, B2 => 
                           n17542, ZN => n15719);
   U13709 : AOI221_X1 port map( B1 => n17599, B2 => n17337, C1 => n17596, C2 =>
                           n16873, A => n15692, ZN => n15689);
   U13710 : OAI22_X1 port map( A1 => n16599, A2 => n17593, B1 => n17163, B2 => 
                           n17590, ZN => n15692);
   U13711 : AOI221_X1 port map( B1 => n17551, B2 => n17338, C1 => n17548, C2 =>
                           n16874, A => n15700, ZN => n15697);
   U13712 : OAI22_X1 port map( A1 => n16563, A2 => n17545, B1 => n17091, B2 => 
                           n17542, ZN => n15700);
   U13713 : AOI221_X1 port map( B1 => n17599, B2 => n17339, C1 => n17596, C2 =>
                           n16875, A => n15673, ZN => n15670);
   U13714 : OAI22_X1 port map( A1 => n16600, A2 => n17593, B1 => n17164, B2 => 
                           n17590, ZN => n15673);
   U13715 : AOI221_X1 port map( B1 => n17551, B2 => n17340, C1 => n17548, C2 =>
                           n16876, A => n15681, ZN => n15678);
   U13716 : OAI22_X1 port map( A1 => n16564, A2 => n17545, B1 => n17092, B2 => 
                           n17542, ZN => n15681);
   U13717 : AOI221_X1 port map( B1 => n17599, B2 => n17341, C1 => n17596, C2 =>
                           n16877, A => n15654, ZN => n15651);
   U13718 : OAI22_X1 port map( A1 => n16601, A2 => n17593, B1 => n17165, B2 => 
                           n17590, ZN => n15654);
   U13719 : AOI221_X1 port map( B1 => n17551, B2 => n17342, C1 => n17548, C2 =>
                           n16878, A => n15662, ZN => n15659);
   U13720 : OAI22_X1 port map( A1 => n16565, A2 => n17545, B1 => n17093, B2 => 
                           n17542, ZN => n15662);
   U13721 : AOI221_X1 port map( B1 => n17599, B2 => n17343, C1 => n17596, C2 =>
                           n16879, A => n15635, ZN => n15632);
   U13722 : OAI22_X1 port map( A1 => n16602, A2 => n17593, B1 => n17166, B2 => 
                           n17590, ZN => n15635);
   U13723 : AOI221_X1 port map( B1 => n17551, B2 => n17344, C1 => n17548, C2 =>
                           n16880, A => n15643, ZN => n15640);
   U13724 : OAI22_X1 port map( A1 => n16566, A2 => n17545, B1 => n17094, B2 => 
                           n17542, ZN => n15643);
   U13725 : AOI221_X1 port map( B1 => n17599, B2 => n17345, C1 => n17596, C2 =>
                           n16881, A => n15616, ZN => n15613);
   U13726 : OAI22_X1 port map( A1 => n16603, A2 => n17593, B1 => n17167, B2 => 
                           n17590, ZN => n15616);
   U13727 : AOI221_X1 port map( B1 => n17551, B2 => n17346, C1 => n17548, C2 =>
                           n16882, A => n15624, ZN => n15621);
   U13728 : OAI22_X1 port map( A1 => n16567, A2 => n17545, B1 => n17095, B2 => 
                           n17542, ZN => n15624);
   U13729 : AOI221_X1 port map( B1 => n17599, B2 => n17347, C1 => n17596, C2 =>
                           n16883, A => n15597, ZN => n15594);
   U13730 : OAI22_X1 port map( A1 => n16604, A2 => n17593, B1 => n17168, B2 => 
                           n17590, ZN => n15597);
   U13731 : AOI221_X1 port map( B1 => n17551, B2 => n17348, C1 => n17548, C2 =>
                           n16884, A => n15605, ZN => n15602);
   U13732 : OAI22_X1 port map( A1 => n16568, A2 => n17545, B1 => n17096, B2 => 
                           n17542, ZN => n15605);
   U13733 : AOI221_X1 port map( B1 => n17599, B2 => n17349, C1 => n17596, C2 =>
                           n16885, A => n15578, ZN => n15575);
   U13734 : OAI22_X1 port map( A1 => n16605, A2 => n17593, B1 => n17169, B2 => 
                           n17590, ZN => n15578);
   U13735 : AOI221_X1 port map( B1 => n17551, B2 => n17350, C1 => n17548, C2 =>
                           n16886, A => n15586, ZN => n15583);
   U13736 : OAI22_X1 port map( A1 => n16569, A2 => n17545, B1 => n17097, B2 => 
                           n17542, ZN => n15586);
   U13737 : AOI221_X1 port map( B1 => n17599, B2 => n17351, C1 => n17596, C2 =>
                           n16887, A => n15559, ZN => n15556);
   U13738 : OAI22_X1 port map( A1 => n16606, A2 => n17593, B1 => n17170, B2 => 
                           n17590, ZN => n15559);
   U13739 : AOI221_X1 port map( B1 => n17551, B2 => n17352, C1 => n17548, C2 =>
                           n16888, A => n15567, ZN => n15564);
   U13740 : OAI22_X1 port map( A1 => n16570, A2 => n17545, B1 => n17098, B2 => 
                           n17542, ZN => n15567);
   U13741 : AOI221_X1 port map( B1 => n17599, B2 => n17353, C1 => n17596, C2 =>
                           n16889, A => n15540, ZN => n15537);
   U13742 : OAI22_X1 port map( A1 => n16607, A2 => n17593, B1 => n17171, B2 => 
                           n17590, ZN => n15540);
   U13743 : AOI221_X1 port map( B1 => n17551, B2 => n17354, C1 => n17548, C2 =>
                           n16890, A => n15548, ZN => n15545);
   U13744 : OAI22_X1 port map( A1 => n16571, A2 => n17545, B1 => n17099, B2 => 
                           n17542, ZN => n15548);
   U13745 : AOI221_X1 port map( B1 => n17599, B2 => n17355, C1 => n17596, C2 =>
                           n16891, A => n15521, ZN => n15518);
   U13746 : OAI22_X1 port map( A1 => n16608, A2 => n17593, B1 => n17172, B2 => 
                           n17590, ZN => n15521);
   U13747 : AOI221_X1 port map( B1 => n17551, B2 => n17356, C1 => n17548, C2 =>
                           n16892, A => n15529, ZN => n15526);
   U13748 : OAI22_X1 port map( A1 => n16572, A2 => n17545, B1 => n17100, B2 => 
                           n17542, ZN => n15529);
   U13749 : AOI221_X1 port map( B1 => n17552, B2 => n17357, C1 => n17549, C2 =>
                           n16893, A => n15510, ZN => n15507);
   U13750 : OAI22_X1 port map( A1 => n16501, A2 => n17546, B1 => n16757, B2 => 
                           n17543, ZN => n15510);
   U13751 : AOI221_X1 port map( B1 => n17552, B2 => n17358, C1 => n17549, C2 =>
                           n16894, A => n15491, ZN => n15488);
   U13752 : OAI22_X1 port map( A1 => n16502, A2 => n17546, B1 => n16758, B2 => 
                           n17543, ZN => n15491);
   U13753 : AOI221_X1 port map( B1 => n17552, B2 => n17359, C1 => n17549, C2 =>
                           n16895, A => n15472, ZN => n15469);
   U13754 : OAI22_X1 port map( A1 => n16503, A2 => n17546, B1 => n16759, B2 => 
                           n17543, ZN => n15472);
   U13755 : AOI221_X1 port map( B1 => n17552, B2 => n17360, C1 => n17549, C2 =>
                           n16896, A => n15453, ZN => n15450);
   U13756 : OAI22_X1 port map( A1 => n16504, A2 => n17546, B1 => n16760, B2 => 
                           n17543, ZN => n15453);
   U13757 : AOI221_X1 port map( B1 => n17552, B2 => n17361, C1 => n17549, C2 =>
                           n16897, A => n15434, ZN => n15431);
   U13758 : OAI22_X1 port map( A1 => n16505, A2 => n17546, B1 => n16761, B2 => 
                           n17543, ZN => n15434);
   U13759 : AOI221_X1 port map( B1 => n17552, B2 => n17362, C1 => n17549, C2 =>
                           n16898, A => n15415, ZN => n15412);
   U13760 : OAI22_X1 port map( A1 => n16506, A2 => n17546, B1 => n16762, B2 => 
                           n17543, ZN => n15415);
   U13761 : AOI221_X1 port map( B1 => n17552, B2 => n17363, C1 => n17549, C2 =>
                           n16899, A => n15396, ZN => n15393);
   U13762 : OAI22_X1 port map( A1 => n16507, A2 => n17546, B1 => n16763, B2 => 
                           n17543, ZN => n15396);
   U13763 : AOI221_X1 port map( B1 => n17552, B2 => n17364, C1 => n17549, C2 =>
                           n16900, A => n15367, ZN => n15358);
   U13764 : OAI22_X1 port map( A1 => n16508, A2 => n17546, B1 => n16764, B2 => 
                           n17543, ZN => n15367);
   U13765 : AOI221_X1 port map( B1 => n17700, B2 => n17309, C1 => n17697, C2 =>
                           n16845, A => n15309, ZN => n15302);
   U13766 : OAI22_X1 port map( A1 => n16701, A2 => n17694, B1 => n17149, B2 => 
                           n17691, ZN => n15309);
   U13767 : AOI221_X1 port map( B1 => n17652, B2 => n17310, C1 => n17649, C2 =>
                           n16846, A => n15323, ZN => n15318);
   U13768 : OAI22_X1 port map( A1 => n16665, A2 => n17646, B1 => n17077, B2 => 
                           n17643, ZN => n15323);
   U13769 : AOI221_X1 port map( B1 => n17700, B2 => n17311, C1 => n17697, C2 =>
                           n16847, A => n15286, ZN => n15283);
   U13770 : OAI22_X1 port map( A1 => n16702, A2 => n17694, B1 => n17150, B2 => 
                           n17691, ZN => n15286);
   U13771 : AOI221_X1 port map( B1 => n17652, B2 => n17312, C1 => n17649, C2 =>
                           n16848, A => n15294, ZN => n15291);
   U13772 : OAI22_X1 port map( A1 => n16666, A2 => n17646, B1 => n17078, B2 => 
                           n17643, ZN => n15294);
   U13773 : AOI221_X1 port map( B1 => n17700, B2 => n17313, C1 => n17697, C2 =>
                           n16849, A => n15267, ZN => n15264);
   U13774 : OAI22_X1 port map( A1 => n16703, A2 => n17694, B1 => n17151, B2 => 
                           n17691, ZN => n15267);
   U13775 : AOI221_X1 port map( B1 => n17652, B2 => n17314, C1 => n17649, C2 =>
                           n16850, A => n15275, ZN => n15272);
   U13776 : OAI22_X1 port map( A1 => n16667, A2 => n17646, B1 => n17079, B2 => 
                           n17643, ZN => n15275);
   U13777 : AOI221_X1 port map( B1 => n17700, B2 => n17315, C1 => n17697, C2 =>
                           n16851, A => n15248, ZN => n15245);
   U13778 : OAI22_X1 port map( A1 => n16704, A2 => n17694, B1 => n17152, B2 => 
                           n17691, ZN => n15248);
   U13779 : AOI221_X1 port map( B1 => n17652, B2 => n17316, C1 => n17649, C2 =>
                           n16852, A => n15256, ZN => n15253);
   U13780 : OAI22_X1 port map( A1 => n16668, A2 => n17646, B1 => n17080, B2 => 
                           n17643, ZN => n15256);
   U13781 : AOI221_X1 port map( B1 => n17700, B2 => n17317, C1 => n17697, C2 =>
                           n16853, A => n15229, ZN => n15226);
   U13782 : OAI22_X1 port map( A1 => n16705, A2 => n17694, B1 => n17153, B2 => 
                           n17691, ZN => n15229);
   U13783 : AOI221_X1 port map( B1 => n17652, B2 => n17318, C1 => n17649, C2 =>
                           n16854, A => n15237, ZN => n15234);
   U13784 : OAI22_X1 port map( A1 => n16669, A2 => n17646, B1 => n17081, B2 => 
                           n17643, ZN => n15237);
   U13785 : AOI221_X1 port map( B1 => n17700, B2 => n17319, C1 => n17697, C2 =>
                           n16855, A => n15210, ZN => n15207);
   U13786 : OAI22_X1 port map( A1 => n16706, A2 => n17694, B1 => n17154, B2 => 
                           n17691, ZN => n15210);
   U13787 : AOI221_X1 port map( B1 => n17652, B2 => n17320, C1 => n17649, C2 =>
                           n16856, A => n15218, ZN => n15215);
   U13788 : OAI22_X1 port map( A1 => n16670, A2 => n17646, B1 => n17082, B2 => 
                           n17643, ZN => n15218);
   U13789 : AOI221_X1 port map( B1 => n17700, B2 => n17321, C1 => n17697, C2 =>
                           n16857, A => n15191, ZN => n15188);
   U13790 : OAI22_X1 port map( A1 => n16707, A2 => n17694, B1 => n17155, B2 => 
                           n17691, ZN => n15191);
   U13791 : AOI221_X1 port map( B1 => n17652, B2 => n17322, C1 => n17649, C2 =>
                           n16858, A => n15199, ZN => n15196);
   U13792 : OAI22_X1 port map( A1 => n16671, A2 => n17646, B1 => n17083, B2 => 
                           n17643, ZN => n15199);
   U13793 : AOI221_X1 port map( B1 => n17700, B2 => n17323, C1 => n17697, C2 =>
                           n16859, A => n15172, ZN => n15169);
   U13794 : OAI22_X1 port map( A1 => n16708, A2 => n17694, B1 => n17156, B2 => 
                           n17691, ZN => n15172);
   U13795 : AOI221_X1 port map( B1 => n17652, B2 => n17324, C1 => n17649, C2 =>
                           n16860, A => n15180, ZN => n15177);
   U13796 : OAI22_X1 port map( A1 => n16672, A2 => n17646, B1 => n17084, B2 => 
                           n17643, ZN => n15180);
   U13797 : AOI221_X1 port map( B1 => n17700, B2 => n17325, C1 => n17697, C2 =>
                           n16861, A => n15153, ZN => n15150);
   U13798 : OAI22_X1 port map( A1 => n16709, A2 => n17694, B1 => n17157, B2 => 
                           n17691, ZN => n15153);
   U13799 : AOI221_X1 port map( B1 => n17652, B2 => n17326, C1 => n17649, C2 =>
                           n16862, A => n15161, ZN => n15158);
   U13800 : OAI22_X1 port map( A1 => n16673, A2 => n17646, B1 => n17085, B2 => 
                           n17643, ZN => n15161);
   U13801 : AOI221_X1 port map( B1 => n17700, B2 => n17327, C1 => n17697, C2 =>
                           n16863, A => n15134, ZN => n15131);
   U13802 : OAI22_X1 port map( A1 => n16710, A2 => n17694, B1 => n17158, B2 => 
                           n17691, ZN => n15134);
   U13803 : AOI221_X1 port map( B1 => n17652, B2 => n17328, C1 => n17649, C2 =>
                           n16864, A => n15142, ZN => n15139);
   U13804 : OAI22_X1 port map( A1 => n16674, A2 => n17646, B1 => n17086, B2 => 
                           n17643, ZN => n15142);
   U13805 : AOI221_X1 port map( B1 => n17700, B2 => n17329, C1 => n17697, C2 =>
                           n16865, A => n15115, ZN => n15112);
   U13806 : OAI22_X1 port map( A1 => n16711, A2 => n17694, B1 => n17159, B2 => 
                           n17691, ZN => n15115);
   U13807 : AOI221_X1 port map( B1 => n17652, B2 => n17330, C1 => n17649, C2 =>
                           n16866, A => n15123, ZN => n15120);
   U13808 : OAI22_X1 port map( A1 => n16675, A2 => n17646, B1 => n17087, B2 => 
                           n17643, ZN => n15123);
   U13809 : AOI221_X1 port map( B1 => n17700, B2 => n17331, C1 => n17697, C2 =>
                           n16867, A => n15096, ZN => n15093);
   U13810 : OAI22_X1 port map( A1 => n16712, A2 => n17694, B1 => n17160, B2 => 
                           n17691, ZN => n15096);
   U13811 : AOI221_X1 port map( B1 => n17652, B2 => n17332, C1 => n17649, C2 =>
                           n16868, A => n15104, ZN => n15101);
   U13812 : OAI22_X1 port map( A1 => n16676, A2 => n17646, B1 => n17088, B2 => 
                           n17643, ZN => n15104);
   U13813 : AOI221_X1 port map( B1 => n17701, B2 => n17333, C1 => n17698, C2 =>
                           n16869, A => n15077, ZN => n15074);
   U13814 : OAI22_X1 port map( A1 => n16597, A2 => n17695, B1 => n17161, B2 => 
                           n17692, ZN => n15077);
   U13815 : AOI221_X1 port map( B1 => n17653, B2 => n17334, C1 => n17650, C2 =>
                           n16870, A => n15085, ZN => n15082);
   U13816 : OAI22_X1 port map( A1 => n16561, A2 => n17647, B1 => n17089, B2 => 
                           n17644, ZN => n15085);
   U13817 : AOI221_X1 port map( B1 => n17701, B2 => n17335, C1 => n17698, C2 =>
                           n16871, A => n15058, ZN => n15055);
   U13818 : OAI22_X1 port map( A1 => n16598, A2 => n17695, B1 => n17162, B2 => 
                           n17692, ZN => n15058);
   U13819 : AOI221_X1 port map( B1 => n17653, B2 => n17336, C1 => n17650, C2 =>
                           n16872, A => n15066, ZN => n15063);
   U13820 : OAI22_X1 port map( A1 => n16562, A2 => n17647, B1 => n17090, B2 => 
                           n17644, ZN => n15066);
   U13821 : AOI221_X1 port map( B1 => n17701, B2 => n17337, C1 => n17698, C2 =>
                           n16873, A => n15039, ZN => n15036);
   U13822 : OAI22_X1 port map( A1 => n16599, A2 => n17695, B1 => n17163, B2 => 
                           n17692, ZN => n15039);
   U13823 : AOI221_X1 port map( B1 => n17653, B2 => n17338, C1 => n17650, C2 =>
                           n16874, A => n15047, ZN => n15044);
   U13824 : OAI22_X1 port map( A1 => n16563, A2 => n17647, B1 => n17091, B2 => 
                           n17644, ZN => n15047);
   U13825 : AOI221_X1 port map( B1 => n17701, B2 => n17339, C1 => n17698, C2 =>
                           n16875, A => n15020, ZN => n15017);
   U13826 : OAI22_X1 port map( A1 => n16600, A2 => n17695, B1 => n17164, B2 => 
                           n17692, ZN => n15020);
   U13827 : AOI221_X1 port map( B1 => n17653, B2 => n17340, C1 => n17650, C2 =>
                           n16876, A => n15028, ZN => n15025);
   U13828 : OAI22_X1 port map( A1 => n16564, A2 => n17647, B1 => n17092, B2 => 
                           n17644, ZN => n15028);
   U13829 : AOI221_X1 port map( B1 => n17701, B2 => n17341, C1 => n17698, C2 =>
                           n16877, A => n15001, ZN => n14998);
   U13830 : OAI22_X1 port map( A1 => n16601, A2 => n17695, B1 => n17165, B2 => 
                           n17692, ZN => n15001);
   U13831 : AOI221_X1 port map( B1 => n17653, B2 => n17342, C1 => n17650, C2 =>
                           n16878, A => n15009, ZN => n15006);
   U13832 : OAI22_X1 port map( A1 => n16565, A2 => n17647, B1 => n17093, B2 => 
                           n17644, ZN => n15009);
   U13833 : AOI221_X1 port map( B1 => n17701, B2 => n17343, C1 => n17698, C2 =>
                           n16879, A => n14982, ZN => n14979);
   U13834 : OAI22_X1 port map( A1 => n16602, A2 => n17695, B1 => n17166, B2 => 
                           n17692, ZN => n14982);
   U13835 : AOI221_X1 port map( B1 => n17653, B2 => n17344, C1 => n17650, C2 =>
                           n16880, A => n14990, ZN => n14987);
   U13836 : OAI22_X1 port map( A1 => n16566, A2 => n17647, B1 => n17094, B2 => 
                           n17644, ZN => n14990);
   U13837 : AOI221_X1 port map( B1 => n17701, B2 => n17345, C1 => n17698, C2 =>
                           n16881, A => n14963, ZN => n14960);
   U13838 : OAI22_X1 port map( A1 => n16603, A2 => n17695, B1 => n17167, B2 => 
                           n17692, ZN => n14963);
   U13839 : AOI221_X1 port map( B1 => n17653, B2 => n17346, C1 => n17650, C2 =>
                           n16882, A => n14971, ZN => n14968);
   U13840 : OAI22_X1 port map( A1 => n16567, A2 => n17647, B1 => n17095, B2 => 
                           n17644, ZN => n14971);
   U13841 : AOI221_X1 port map( B1 => n17701, B2 => n17347, C1 => n17698, C2 =>
                           n16883, A => n14944, ZN => n14941);
   U13842 : OAI22_X1 port map( A1 => n16604, A2 => n17695, B1 => n17168, B2 => 
                           n17692, ZN => n14944);
   U13843 : AOI221_X1 port map( B1 => n17653, B2 => n17348, C1 => n17650, C2 =>
                           n16884, A => n14952, ZN => n14949);
   U13844 : OAI22_X1 port map( A1 => n16568, A2 => n17647, B1 => n17096, B2 => 
                           n17644, ZN => n14952);
   U13845 : AOI221_X1 port map( B1 => n17701, B2 => n17349, C1 => n17698, C2 =>
                           n16885, A => n14925, ZN => n14922);
   U13846 : OAI22_X1 port map( A1 => n16605, A2 => n17695, B1 => n17169, B2 => 
                           n17692, ZN => n14925);
   U13847 : AOI221_X1 port map( B1 => n17653, B2 => n17350, C1 => n17650, C2 =>
                           n16886, A => n14933, ZN => n14930);
   U13848 : OAI22_X1 port map( A1 => n16569, A2 => n17647, B1 => n17097, B2 => 
                           n17644, ZN => n14933);
   U13849 : AOI221_X1 port map( B1 => n17701, B2 => n17351, C1 => n17698, C2 =>
                           n16887, A => n14906, ZN => n14903);
   U13850 : OAI22_X1 port map( A1 => n16606, A2 => n17695, B1 => n17170, B2 => 
                           n17692, ZN => n14906);
   U13851 : AOI221_X1 port map( B1 => n17653, B2 => n17352, C1 => n17650, C2 =>
                           n16888, A => n14914, ZN => n14911);
   U13852 : OAI22_X1 port map( A1 => n16570, A2 => n17647, B1 => n17098, B2 => 
                           n17644, ZN => n14914);
   U13853 : AOI221_X1 port map( B1 => n17701, B2 => n17353, C1 => n17698, C2 =>
                           n16889, A => n14887, ZN => n14884);
   U13854 : OAI22_X1 port map( A1 => n16607, A2 => n17695, B1 => n17171, B2 => 
                           n17692, ZN => n14887);
   U13855 : AOI221_X1 port map( B1 => n17653, B2 => n17354, C1 => n17650, C2 =>
                           n16890, A => n14895, ZN => n14892);
   U13856 : OAI22_X1 port map( A1 => n16571, A2 => n17647, B1 => n17099, B2 => 
                           n17644, ZN => n14895);
   U13857 : AOI221_X1 port map( B1 => n17701, B2 => n17355, C1 => n17698, C2 =>
                           n16891, A => n14868, ZN => n14865);
   U13858 : OAI22_X1 port map( A1 => n16608, A2 => n17695, B1 => n17172, B2 => 
                           n17692, ZN => n14868);
   U13859 : AOI221_X1 port map( B1 => n17653, B2 => n17356, C1 => n17650, C2 =>
                           n16892, A => n14876, ZN => n14873);
   U13860 : OAI22_X1 port map( A1 => n16572, A2 => n17647, B1 => n17100, B2 => 
                           n17644, ZN => n14876);
   U13861 : AOI221_X1 port map( B1 => n17654, B2 => n17357, C1 => n17651, C2 =>
                           n16893, A => n14857, ZN => n14854);
   U13862 : OAI22_X1 port map( A1 => n16501, A2 => n17648, B1 => n16757, B2 => 
                           n17645, ZN => n14857);
   U13863 : AOI221_X1 port map( B1 => n17654, B2 => n17358, C1 => n17651, C2 =>
                           n16894, A => n14838, ZN => n14835);
   U13864 : OAI22_X1 port map( A1 => n16502, A2 => n17648, B1 => n16758, B2 => 
                           n17645, ZN => n14838);
   U13865 : AOI221_X1 port map( B1 => n17654, B2 => n17359, C1 => n17651, C2 =>
                           n16895, A => n14819, ZN => n14816);
   U13866 : OAI22_X1 port map( A1 => n16503, A2 => n17648, B1 => n16759, B2 => 
                           n17645, ZN => n14819);
   U13867 : AOI221_X1 port map( B1 => n17654, B2 => n17360, C1 => n17651, C2 =>
                           n16896, A => n14800, ZN => n14797);
   U13868 : OAI22_X1 port map( A1 => n16504, A2 => n17648, B1 => n16760, B2 => 
                           n17645, ZN => n14800);
   U13869 : AOI221_X1 port map( B1 => n17654, B2 => n17361, C1 => n17651, C2 =>
                           n16897, A => n14781, ZN => n14778);
   U13870 : OAI22_X1 port map( A1 => n16505, A2 => n17648, B1 => n16761, B2 => 
                           n17645, ZN => n14781);
   U13871 : AOI221_X1 port map( B1 => n17654, B2 => n17362, C1 => n17651, C2 =>
                           n16898, A => n14762, ZN => n14759);
   U13872 : OAI22_X1 port map( A1 => n16506, A2 => n17648, B1 => n16762, B2 => 
                           n17645, ZN => n14762);
   U13873 : AOI221_X1 port map( B1 => n17654, B2 => n17363, C1 => n17651, C2 =>
                           n16899, A => n14743, ZN => n14740);
   U13874 : OAI22_X1 port map( A1 => n16507, A2 => n17648, B1 => n16763, B2 => 
                           n17645, ZN => n14743);
   U13875 : AOI221_X1 port map( B1 => n17654, B2 => n17364, C1 => n17651, C2 =>
                           n16900, A => n14714, ZN => n14705);
   U13876 : OAI22_X1 port map( A1 => n16508, A2 => n17648, B1 => n16764, B2 => 
                           n17645, ZN => n14714);
   U13877 : AOI221_X1 port map( B1 => n17586, B2 => n17365, C1 => n17583, C2 =>
                           n16901, A => n15965, ZN => n15954);
   U13878 : OAI22_X1 port map( A1 => n16713, A2 => n17580, B1 => n17173, B2 => 
                           n17577, ZN => n15965);
   U13879 : AOI221_X1 port map( B1 => n17538, B2 => n17366, C1 => n17535, C2 =>
                           n16902, A => n15977, ZN => n15970);
   U13880 : OAI22_X1 port map( A1 => n16677, A2 => n17532, B1 => n17101, B2 => 
                           n17529, ZN => n15977);
   U13881 : AOI221_X1 port map( B1 => n17586, B2 => n17367, C1 => n17583, C2 =>
                           n16903, A => n15940, ZN => n15935);
   U13882 : OAI22_X1 port map( A1 => n16714, A2 => n17580, B1 => n17174, B2 => 
                           n17577, ZN => n15940);
   U13883 : AOI221_X1 port map( B1 => n17538, B2 => n17368, C1 => n17535, C2 =>
                           n16904, A => n15948, ZN => n15943);
   U13884 : OAI22_X1 port map( A1 => n16678, A2 => n17532, B1 => n17102, B2 => 
                           n17529, ZN => n15948);
   U13885 : AOI221_X1 port map( B1 => n17586, B2 => n17369, C1 => n17583, C2 =>
                           n16905, A => n15921, ZN => n15916);
   U13886 : OAI22_X1 port map( A1 => n16715, A2 => n17580, B1 => n17175, B2 => 
                           n17577, ZN => n15921);
   U13887 : AOI221_X1 port map( B1 => n17538, B2 => n17370, C1 => n17535, C2 =>
                           n16906, A => n15929, ZN => n15924);
   U13888 : OAI22_X1 port map( A1 => n16679, A2 => n17532, B1 => n17103, B2 => 
                           n17529, ZN => n15929);
   U13889 : AOI221_X1 port map( B1 => n17586, B2 => n17371, C1 => n17583, C2 =>
                           n16907, A => n15902, ZN => n15897);
   U13890 : OAI22_X1 port map( A1 => n16716, A2 => n17580, B1 => n17176, B2 => 
                           n17577, ZN => n15902);
   U13891 : AOI221_X1 port map( B1 => n17538, B2 => n17372, C1 => n17535, C2 =>
                           n16908, A => n15910, ZN => n15905);
   U13892 : OAI22_X1 port map( A1 => n16680, A2 => n17532, B1 => n17104, B2 => 
                           n17529, ZN => n15910);
   U13893 : AOI221_X1 port map( B1 => n17586, B2 => n17373, C1 => n17583, C2 =>
                           n16909, A => n15883, ZN => n15878);
   U13894 : OAI22_X1 port map( A1 => n16717, A2 => n17580, B1 => n17177, B2 => 
                           n17577, ZN => n15883);
   U13895 : AOI221_X1 port map( B1 => n17538, B2 => n17374, C1 => n17535, C2 =>
                           n16910, A => n15891, ZN => n15886);
   U13896 : OAI22_X1 port map( A1 => n16681, A2 => n17532, B1 => n17105, B2 => 
                           n17529, ZN => n15891);
   U13897 : AOI221_X1 port map( B1 => n17586, B2 => n17375, C1 => n17583, C2 =>
                           n16911, A => n15864, ZN => n15859);
   U13898 : OAI22_X1 port map( A1 => n16718, A2 => n17580, B1 => n17178, B2 => 
                           n17577, ZN => n15864);
   U13899 : AOI221_X1 port map( B1 => n17538, B2 => n17376, C1 => n17535, C2 =>
                           n16912, A => n15872, ZN => n15867);
   U13900 : OAI22_X1 port map( A1 => n16682, A2 => n17532, B1 => n17106, B2 => 
                           n17529, ZN => n15872);
   U13901 : AOI221_X1 port map( B1 => n17586, B2 => n17377, C1 => n17583, C2 =>
                           n16913, A => n15845, ZN => n15840);
   U13902 : OAI22_X1 port map( A1 => n16719, A2 => n17580, B1 => n17179, B2 => 
                           n17577, ZN => n15845);
   U13903 : AOI221_X1 port map( B1 => n17538, B2 => n17378, C1 => n17535, C2 =>
                           n16914, A => n15853, ZN => n15848);
   U13904 : OAI22_X1 port map( A1 => n16683, A2 => n17532, B1 => n17107, B2 => 
                           n17529, ZN => n15853);
   U13905 : AOI221_X1 port map( B1 => n17586, B2 => n17379, C1 => n17583, C2 =>
                           n16915, A => n15826, ZN => n15821);
   U13906 : OAI22_X1 port map( A1 => n16720, A2 => n17580, B1 => n17180, B2 => 
                           n17577, ZN => n15826);
   U13907 : AOI221_X1 port map( B1 => n17538, B2 => n17380, C1 => n17535, C2 =>
                           n16916, A => n15834, ZN => n15829);
   U13908 : OAI22_X1 port map( A1 => n16684, A2 => n17532, B1 => n17108, B2 => 
                           n17529, ZN => n15834);
   U13909 : AOI221_X1 port map( B1 => n17586, B2 => n17381, C1 => n17583, C2 =>
                           n16917, A => n15807, ZN => n15802);
   U13910 : OAI22_X1 port map( A1 => n16721, A2 => n17580, B1 => n17181, B2 => 
                           n17577, ZN => n15807);
   U13911 : AOI221_X1 port map( B1 => n17538, B2 => n17382, C1 => n17535, C2 =>
                           n16918, A => n15815, ZN => n15810);
   U13912 : OAI22_X1 port map( A1 => n16685, A2 => n17532, B1 => n17109, B2 => 
                           n17529, ZN => n15815);
   U13913 : AOI221_X1 port map( B1 => n17586, B2 => n17383, C1 => n17583, C2 =>
                           n16919, A => n15788, ZN => n15783);
   U13914 : OAI22_X1 port map( A1 => n16722, A2 => n17580, B1 => n17182, B2 => 
                           n17577, ZN => n15788);
   U13915 : AOI221_X1 port map( B1 => n17538, B2 => n17384, C1 => n17535, C2 =>
                           n16920, A => n15796, ZN => n15791);
   U13916 : OAI22_X1 port map( A1 => n16686, A2 => n17532, B1 => n17110, B2 => 
                           n17529, ZN => n15796);
   U13917 : AOI221_X1 port map( B1 => n17586, B2 => n17385, C1 => n17583, C2 =>
                           n16921, A => n15769, ZN => n15764);
   U13918 : OAI22_X1 port map( A1 => n16723, A2 => n17580, B1 => n17183, B2 => 
                           n17577, ZN => n15769);
   U13919 : AOI221_X1 port map( B1 => n17538, B2 => n17386, C1 => n17535, C2 =>
                           n16922, A => n15777, ZN => n15772);
   U13920 : OAI22_X1 port map( A1 => n16687, A2 => n17532, B1 => n17111, B2 => 
                           n17529, ZN => n15777);
   U13921 : AOI221_X1 port map( B1 => n17586, B2 => n17387, C1 => n17583, C2 =>
                           n16923, A => n15750, ZN => n15745);
   U13922 : OAI22_X1 port map( A1 => n16724, A2 => n17580, B1 => n17184, B2 => 
                           n17577, ZN => n15750);
   U13923 : AOI221_X1 port map( B1 => n17538, B2 => n17388, C1 => n17535, C2 =>
                           n16924, A => n15758, ZN => n15753);
   U13924 : OAI22_X1 port map( A1 => n16688, A2 => n17532, B1 => n17112, B2 => 
                           n17529, ZN => n15758);
   U13925 : AOI221_X1 port map( B1 => n17587, B2 => n17389, C1 => n17584, C2 =>
                           n16925, A => n15731, ZN => n15726);
   U13926 : OAI22_X1 port map( A1 => n16609, A2 => n17581, B1 => n17185, B2 => 
                           n17578, ZN => n15731);
   U13927 : AOI221_X1 port map( B1 => n17539, B2 => n17390, C1 => n17536, C2 =>
                           n16926, A => n15739, ZN => n15734);
   U13928 : OAI22_X1 port map( A1 => n16573, A2 => n17533, B1 => n17113, B2 => 
                           n17530, ZN => n15739);
   U13929 : AOI221_X1 port map( B1 => n17587, B2 => n17391, C1 => n17584, C2 =>
                           n16927, A => n15712, ZN => n15707);
   U13930 : OAI22_X1 port map( A1 => n16610, A2 => n17581, B1 => n17186, B2 => 
                           n17578, ZN => n15712);
   U13931 : AOI221_X1 port map( B1 => n17539, B2 => n17392, C1 => n17536, C2 =>
                           n16928, A => n15720, ZN => n15715);
   U13932 : OAI22_X1 port map( A1 => n16574, A2 => n17533, B1 => n17114, B2 => 
                           n17530, ZN => n15720);
   U13933 : AOI221_X1 port map( B1 => n17587, B2 => n17393, C1 => n17584, C2 =>
                           n16929, A => n15693, ZN => n15688);
   U13934 : OAI22_X1 port map( A1 => n16611, A2 => n17581, B1 => n17187, B2 => 
                           n17578, ZN => n15693);
   U13935 : AOI221_X1 port map( B1 => n17539, B2 => n17394, C1 => n17536, C2 =>
                           n16930, A => n15701, ZN => n15696);
   U13936 : OAI22_X1 port map( A1 => n16575, A2 => n17533, B1 => n17115, B2 => 
                           n17530, ZN => n15701);
   U13937 : AOI221_X1 port map( B1 => n17587, B2 => n17395, C1 => n17584, C2 =>
                           n16931, A => n15674, ZN => n15669);
   U13938 : OAI22_X1 port map( A1 => n16612, A2 => n17581, B1 => n17188, B2 => 
                           n17578, ZN => n15674);
   U13939 : AOI221_X1 port map( B1 => n17539, B2 => n17396, C1 => n17536, C2 =>
                           n16932, A => n15682, ZN => n15677);
   U13940 : OAI22_X1 port map( A1 => n16576, A2 => n17533, B1 => n17116, B2 => 
                           n17530, ZN => n15682);
   U13941 : AOI221_X1 port map( B1 => n17587, B2 => n17397, C1 => n17584, C2 =>
                           n16933, A => n15655, ZN => n15650);
   U13942 : OAI22_X1 port map( A1 => n16613, A2 => n17581, B1 => n17189, B2 => 
                           n17578, ZN => n15655);
   U13943 : AOI221_X1 port map( B1 => n17539, B2 => n17398, C1 => n17536, C2 =>
                           n16934, A => n15663, ZN => n15658);
   U13944 : OAI22_X1 port map( A1 => n16577, A2 => n17533, B1 => n17117, B2 => 
                           n17530, ZN => n15663);
   U13945 : AOI221_X1 port map( B1 => n17587, B2 => n17399, C1 => n17584, C2 =>
                           n16935, A => n15636, ZN => n15631);
   U13946 : OAI22_X1 port map( A1 => n16614, A2 => n17581, B1 => n17190, B2 => 
                           n17578, ZN => n15636);
   U13947 : AOI221_X1 port map( B1 => n17539, B2 => n17400, C1 => n17536, C2 =>
                           n16936, A => n15644, ZN => n15639);
   U13948 : OAI22_X1 port map( A1 => n16578, A2 => n17533, B1 => n17118, B2 => 
                           n17530, ZN => n15644);
   U13949 : AOI221_X1 port map( B1 => n17587, B2 => n17401, C1 => n17584, C2 =>
                           n16937, A => n15617, ZN => n15612);
   U13950 : OAI22_X1 port map( A1 => n16615, A2 => n17581, B1 => n17191, B2 => 
                           n17578, ZN => n15617);
   U13951 : AOI221_X1 port map( B1 => n17539, B2 => n17402, C1 => n17536, C2 =>
                           n16938, A => n15625, ZN => n15620);
   U13952 : OAI22_X1 port map( A1 => n16579, A2 => n17533, B1 => n17119, B2 => 
                           n17530, ZN => n15625);
   U13953 : AOI221_X1 port map( B1 => n17587, B2 => n17403, C1 => n17584, C2 =>
                           n16939, A => n15598, ZN => n15593);
   U13954 : OAI22_X1 port map( A1 => n16616, A2 => n17581, B1 => n17192, B2 => 
                           n17578, ZN => n15598);
   U13955 : AOI221_X1 port map( B1 => n17539, B2 => n17404, C1 => n17536, C2 =>
                           n16940, A => n15606, ZN => n15601);
   U13956 : OAI22_X1 port map( A1 => n16580, A2 => n17533, B1 => n17120, B2 => 
                           n17530, ZN => n15606);
   U13957 : AOI221_X1 port map( B1 => n17587, B2 => n17405, C1 => n17584, C2 =>
                           n16941, A => n15579, ZN => n15574);
   U13958 : OAI22_X1 port map( A1 => n16617, A2 => n17581, B1 => n17193, B2 => 
                           n17578, ZN => n15579);
   U13959 : AOI221_X1 port map( B1 => n17539, B2 => n17406, C1 => n17536, C2 =>
                           n16942, A => n15587, ZN => n15582);
   U13960 : OAI22_X1 port map( A1 => n16581, A2 => n17533, B1 => n17121, B2 => 
                           n17530, ZN => n15587);
   U13961 : AOI221_X1 port map( B1 => n17587, B2 => n17407, C1 => n17584, C2 =>
                           n16943, A => n15560, ZN => n15555);
   U13962 : OAI22_X1 port map( A1 => n16618, A2 => n17581, B1 => n17194, B2 => 
                           n17578, ZN => n15560);
   U13963 : AOI221_X1 port map( B1 => n17539, B2 => n17408, C1 => n17536, C2 =>
                           n16944, A => n15568, ZN => n15563);
   U13964 : OAI22_X1 port map( A1 => n16582, A2 => n17533, B1 => n17122, B2 => 
                           n17530, ZN => n15568);
   U13965 : AOI221_X1 port map( B1 => n17587, B2 => n17409, C1 => n17584, C2 =>
                           n16945, A => n15541, ZN => n15536);
   U13966 : OAI22_X1 port map( A1 => n16619, A2 => n17581, B1 => n17195, B2 => 
                           n17578, ZN => n15541);
   U13967 : AOI221_X1 port map( B1 => n17539, B2 => n17410, C1 => n17536, C2 =>
                           n16946, A => n15549, ZN => n15544);
   U13968 : OAI22_X1 port map( A1 => n16583, A2 => n17533, B1 => n17123, B2 => 
                           n17530, ZN => n15549);
   U13969 : AOI221_X1 port map( B1 => n17587, B2 => n17411, C1 => n17584, C2 =>
                           n16947, A => n15522, ZN => n15517);
   U13970 : OAI22_X1 port map( A1 => n16620, A2 => n17581, B1 => n17196, B2 => 
                           n17578, ZN => n15522);
   U13971 : AOI221_X1 port map( B1 => n17539, B2 => n17412, C1 => n17536, C2 =>
                           n16948, A => n15530, ZN => n15525);
   U13972 : OAI22_X1 port map( A1 => n16584, A2 => n17533, B1 => n17124, B2 => 
                           n17530, ZN => n15530);
   U13973 : AOI221_X1 port map( B1 => n17588, B2 => n17413, C1 => n17585, C2 =>
                           n16949, A => n15503, ZN => n15498);
   U13974 : OAI22_X1 port map( A1 => n16533, A2 => n17582, B1 => n16789, B2 => 
                           n17579, ZN => n15503);
   U13975 : AOI221_X1 port map( B1 => n17540, B2 => n17414, C1 => n17537, C2 =>
                           n16950, A => n15511, ZN => n15506);
   U13976 : OAI22_X1 port map( A1 => n16509, A2 => n17534, B1 => n16765, B2 => 
                           n17531, ZN => n15511);
   U13977 : AOI221_X1 port map( B1 => n17588, B2 => n17415, C1 => n17585, C2 =>
                           n16951, A => n15484, ZN => n15479);
   U13978 : OAI22_X1 port map( A1 => n16534, A2 => n17582, B1 => n16790, B2 => 
                           n17579, ZN => n15484);
   U13979 : AOI221_X1 port map( B1 => n17540, B2 => n17416, C1 => n17537, C2 =>
                           n16952, A => n15492, ZN => n15487);
   U13980 : OAI22_X1 port map( A1 => n16510, A2 => n17534, B1 => n16766, B2 => 
                           n17531, ZN => n15492);
   U13981 : AOI221_X1 port map( B1 => n17588, B2 => n17417, C1 => n17585, C2 =>
                           n16953, A => n15465, ZN => n15460);
   U13982 : OAI22_X1 port map( A1 => n16535, A2 => n17582, B1 => n16791, B2 => 
                           n17579, ZN => n15465);
   U13983 : AOI221_X1 port map( B1 => n17540, B2 => n17418, C1 => n17537, C2 =>
                           n16954, A => n15473, ZN => n15468);
   U13984 : OAI22_X1 port map( A1 => n16511, A2 => n17534, B1 => n16767, B2 => 
                           n17531, ZN => n15473);
   U13985 : AOI221_X1 port map( B1 => n17588, B2 => n17419, C1 => n17585, C2 =>
                           n16955, A => n15446, ZN => n15441);
   U13986 : OAI22_X1 port map( A1 => n16536, A2 => n17582, B1 => n16792, B2 => 
                           n17579, ZN => n15446);
   U13987 : AOI221_X1 port map( B1 => n17540, B2 => n17420, C1 => n17537, C2 =>
                           n16956, A => n15454, ZN => n15449);
   U13988 : OAI22_X1 port map( A1 => n16512, A2 => n17534, B1 => n16768, B2 => 
                           n17531, ZN => n15454);
   U13989 : AOI221_X1 port map( B1 => n17588, B2 => n17421, C1 => n17585, C2 =>
                           n16957, A => n15427, ZN => n15422);
   U13990 : OAI22_X1 port map( A1 => n16537, A2 => n17582, B1 => n16793, B2 => 
                           n17579, ZN => n15427);
   U13991 : AOI221_X1 port map( B1 => n17540, B2 => n17422, C1 => n17537, C2 =>
                           n16958, A => n15435, ZN => n15430);
   U13992 : OAI22_X1 port map( A1 => n16513, A2 => n17534, B1 => n16769, B2 => 
                           n17531, ZN => n15435);
   U13993 : AOI221_X1 port map( B1 => n17588, B2 => n17423, C1 => n17585, C2 =>
                           n16959, A => n15408, ZN => n15403);
   U13994 : OAI22_X1 port map( A1 => n16538, A2 => n17582, B1 => n16794, B2 => 
                           n17579, ZN => n15408);
   U13995 : AOI221_X1 port map( B1 => n17540, B2 => n17424, C1 => n17537, C2 =>
                           n16960, A => n15416, ZN => n15411);
   U13996 : OAI22_X1 port map( A1 => n16514, A2 => n17534, B1 => n16770, B2 => 
                           n17531, ZN => n15416);
   U13997 : AOI221_X1 port map( B1 => n17588, B2 => n17425, C1 => n17585, C2 =>
                           n16961, A => n15389, ZN => n15384);
   U13998 : OAI22_X1 port map( A1 => n16539, A2 => n17582, B1 => n16795, B2 => 
                           n17579, ZN => n15389);
   U13999 : AOI221_X1 port map( B1 => n17540, B2 => n17426, C1 => n17537, C2 =>
                           n16962, A => n15397, ZN => n15392);
   U14000 : OAI22_X1 port map( A1 => n16515, A2 => n17534, B1 => n16771, B2 => 
                           n17531, ZN => n15397);
   U14001 : AOI221_X1 port map( B1 => n17588, B2 => n17427, C1 => n17585, C2 =>
                           n16963, A => n15348, ZN => n15333);
   U14002 : OAI22_X1 port map( A1 => n16540, A2 => n17582, B1 => n16796, B2 => 
                           n17579, ZN => n15348);
   U14003 : AOI221_X1 port map( B1 => n17540, B2 => n17428, C1 => n17537, C2 =>
                           n16964, A => n15372, ZN => n15357);
   U14004 : OAI22_X1 port map( A1 => n16516, A2 => n17534, B1 => n16772, B2 => 
                           n17531, ZN => n15372);
   U14005 : AOI221_X1 port map( B1 => n17688, B2 => n17365, C1 => n17685, C2 =>
                           n16901, A => n15312, ZN => n15301);
   U14006 : OAI22_X1 port map( A1 => n16713, A2 => n17682, B1 => n17173, B2 => 
                           n17679, ZN => n15312);
   U14007 : AOI221_X1 port map( B1 => n17640, B2 => n17366, C1 => n17637, C2 =>
                           n16902, A => n15324, ZN => n15317);
   U14008 : OAI22_X1 port map( A1 => n16677, A2 => n17634, B1 => n17101, B2 => 
                           n17631, ZN => n15324);
   U14009 : AOI221_X1 port map( B1 => n17688, B2 => n17367, C1 => n17685, C2 =>
                           n16903, A => n15287, ZN => n15282);
   U14010 : OAI22_X1 port map( A1 => n16714, A2 => n17682, B1 => n17174, B2 => 
                           n17679, ZN => n15287);
   U14011 : AOI221_X1 port map( B1 => n17640, B2 => n17368, C1 => n17637, C2 =>
                           n16904, A => n15295, ZN => n15290);
   U14012 : OAI22_X1 port map( A1 => n16678, A2 => n17634, B1 => n17102, B2 => 
                           n17631, ZN => n15295);
   U14013 : AOI221_X1 port map( B1 => n17688, B2 => n17369, C1 => n17685, C2 =>
                           n16905, A => n15268, ZN => n15263);
   U14014 : OAI22_X1 port map( A1 => n16715, A2 => n17682, B1 => n17175, B2 => 
                           n17679, ZN => n15268);
   U14015 : AOI221_X1 port map( B1 => n17640, B2 => n17370, C1 => n17637, C2 =>
                           n16906, A => n15276, ZN => n15271);
   U14016 : OAI22_X1 port map( A1 => n16679, A2 => n17634, B1 => n17103, B2 => 
                           n17631, ZN => n15276);
   U14017 : AOI221_X1 port map( B1 => n17688, B2 => n17371, C1 => n17685, C2 =>
                           n16907, A => n15249, ZN => n15244);
   U14018 : OAI22_X1 port map( A1 => n16716, A2 => n17682, B1 => n17176, B2 => 
                           n17679, ZN => n15249);
   U14019 : AOI221_X1 port map( B1 => n17640, B2 => n17372, C1 => n17637, C2 =>
                           n16908, A => n15257, ZN => n15252);
   U14020 : OAI22_X1 port map( A1 => n16680, A2 => n17634, B1 => n17104, B2 => 
                           n17631, ZN => n15257);
   U14021 : AOI221_X1 port map( B1 => n17688, B2 => n17373, C1 => n17685, C2 =>
                           n16909, A => n15230, ZN => n15225);
   U14022 : OAI22_X1 port map( A1 => n16717, A2 => n17682, B1 => n17177, B2 => 
                           n17679, ZN => n15230);
   U14023 : AOI221_X1 port map( B1 => n17640, B2 => n17374, C1 => n17637, C2 =>
                           n16910, A => n15238, ZN => n15233);
   U14024 : OAI22_X1 port map( A1 => n16681, A2 => n17634, B1 => n17105, B2 => 
                           n17631, ZN => n15238);
   U14025 : AOI221_X1 port map( B1 => n17688, B2 => n17375, C1 => n17685, C2 =>
                           n16911, A => n15211, ZN => n15206);
   U14026 : OAI22_X1 port map( A1 => n16718, A2 => n17682, B1 => n17178, B2 => 
                           n17679, ZN => n15211);
   U14027 : AOI221_X1 port map( B1 => n17640, B2 => n17376, C1 => n17637, C2 =>
                           n16912, A => n15219, ZN => n15214);
   U14028 : OAI22_X1 port map( A1 => n16682, A2 => n17634, B1 => n17106, B2 => 
                           n17631, ZN => n15219);
   U14029 : AOI221_X1 port map( B1 => n17688, B2 => n17377, C1 => n17685, C2 =>
                           n16913, A => n15192, ZN => n15187);
   U14030 : OAI22_X1 port map( A1 => n16719, A2 => n17682, B1 => n17179, B2 => 
                           n17679, ZN => n15192);
   U14031 : AOI221_X1 port map( B1 => n17640, B2 => n17378, C1 => n17637, C2 =>
                           n16914, A => n15200, ZN => n15195);
   U14032 : OAI22_X1 port map( A1 => n16683, A2 => n17634, B1 => n17107, B2 => 
                           n17631, ZN => n15200);
   U14033 : AOI221_X1 port map( B1 => n17688, B2 => n17379, C1 => n17685, C2 =>
                           n16915, A => n15173, ZN => n15168);
   U14034 : OAI22_X1 port map( A1 => n16720, A2 => n17682, B1 => n17180, B2 => 
                           n17679, ZN => n15173);
   U14035 : AOI221_X1 port map( B1 => n17640, B2 => n17380, C1 => n17637, C2 =>
                           n16916, A => n15181, ZN => n15176);
   U14036 : OAI22_X1 port map( A1 => n16684, A2 => n17634, B1 => n17108, B2 => 
                           n17631, ZN => n15181);
   U14037 : AOI221_X1 port map( B1 => n17688, B2 => n17381, C1 => n17685, C2 =>
                           n16917, A => n15154, ZN => n15149);
   U14038 : OAI22_X1 port map( A1 => n16721, A2 => n17682, B1 => n17181, B2 => 
                           n17679, ZN => n15154);
   U14039 : AOI221_X1 port map( B1 => n17640, B2 => n17382, C1 => n17637, C2 =>
                           n16918, A => n15162, ZN => n15157);
   U14040 : OAI22_X1 port map( A1 => n16685, A2 => n17634, B1 => n17109, B2 => 
                           n17631, ZN => n15162);
   U14041 : AOI221_X1 port map( B1 => n17688, B2 => n17383, C1 => n17685, C2 =>
                           n16919, A => n15135, ZN => n15130);
   U14042 : OAI22_X1 port map( A1 => n16722, A2 => n17682, B1 => n17182, B2 => 
                           n17679, ZN => n15135);
   U14043 : AOI221_X1 port map( B1 => n17640, B2 => n17384, C1 => n17637, C2 =>
                           n16920, A => n15143, ZN => n15138);
   U14044 : OAI22_X1 port map( A1 => n16686, A2 => n17634, B1 => n17110, B2 => 
                           n17631, ZN => n15143);
   U14045 : AOI221_X1 port map( B1 => n17688, B2 => n17385, C1 => n17685, C2 =>
                           n16921, A => n15116, ZN => n15111);
   U14046 : OAI22_X1 port map( A1 => n16723, A2 => n17682, B1 => n17183, B2 => 
                           n17679, ZN => n15116);
   U14047 : AOI221_X1 port map( B1 => n17640, B2 => n17386, C1 => n17637, C2 =>
                           n16922, A => n15124, ZN => n15119);
   U14048 : OAI22_X1 port map( A1 => n16687, A2 => n17634, B1 => n17111, B2 => 
                           n17631, ZN => n15124);
   U14049 : AOI221_X1 port map( B1 => n17688, B2 => n17387, C1 => n17685, C2 =>
                           n16923, A => n15097, ZN => n15092);
   U14050 : OAI22_X1 port map( A1 => n16724, A2 => n17682, B1 => n17184, B2 => 
                           n17679, ZN => n15097);
   U14051 : AOI221_X1 port map( B1 => n17640, B2 => n17388, C1 => n17637, C2 =>
                           n16924, A => n15105, ZN => n15100);
   U14052 : OAI22_X1 port map( A1 => n16688, A2 => n17634, B1 => n17112, B2 => 
                           n17631, ZN => n15105);
   U14053 : AOI221_X1 port map( B1 => n17689, B2 => n17389, C1 => n17686, C2 =>
                           n16925, A => n15078, ZN => n15073);
   U14054 : OAI22_X1 port map( A1 => n16609, A2 => n17683, B1 => n17185, B2 => 
                           n17680, ZN => n15078);
   U14055 : AOI221_X1 port map( B1 => n17641, B2 => n17390, C1 => n17638, C2 =>
                           n16926, A => n15086, ZN => n15081);
   U14056 : OAI22_X1 port map( A1 => n16573, A2 => n17635, B1 => n17113, B2 => 
                           n17632, ZN => n15086);
   U14057 : AOI221_X1 port map( B1 => n17689, B2 => n17391, C1 => n17686, C2 =>
                           n16927, A => n15059, ZN => n15054);
   U14058 : OAI22_X1 port map( A1 => n16610, A2 => n17683, B1 => n17186, B2 => 
                           n17680, ZN => n15059);
   U14059 : AOI221_X1 port map( B1 => n17641, B2 => n17392, C1 => n17638, C2 =>
                           n16928, A => n15067, ZN => n15062);
   U14060 : OAI22_X1 port map( A1 => n16574, A2 => n17635, B1 => n17114, B2 => 
                           n17632, ZN => n15067);
   U14061 : AOI221_X1 port map( B1 => n17689, B2 => n17393, C1 => n17686, C2 =>
                           n16929, A => n15040, ZN => n15035);
   U14062 : OAI22_X1 port map( A1 => n16611, A2 => n17683, B1 => n17187, B2 => 
                           n17680, ZN => n15040);
   U14063 : AOI221_X1 port map( B1 => n17641, B2 => n17394, C1 => n17638, C2 =>
                           n16930, A => n15048, ZN => n15043);
   U14064 : OAI22_X1 port map( A1 => n16575, A2 => n17635, B1 => n17115, B2 => 
                           n17632, ZN => n15048);
   U14065 : AOI221_X1 port map( B1 => n17689, B2 => n17395, C1 => n17686, C2 =>
                           n16931, A => n15021, ZN => n15016);
   U14066 : OAI22_X1 port map( A1 => n16612, A2 => n17683, B1 => n17188, B2 => 
                           n17680, ZN => n15021);
   U14067 : AOI221_X1 port map( B1 => n17641, B2 => n17396, C1 => n17638, C2 =>
                           n16932, A => n15029, ZN => n15024);
   U14068 : OAI22_X1 port map( A1 => n16576, A2 => n17635, B1 => n17116, B2 => 
                           n17632, ZN => n15029);
   U14069 : AOI221_X1 port map( B1 => n17689, B2 => n17397, C1 => n17686, C2 =>
                           n16933, A => n15002, ZN => n14997);
   U14070 : OAI22_X1 port map( A1 => n16613, A2 => n17683, B1 => n17189, B2 => 
                           n17680, ZN => n15002);
   U14071 : AOI221_X1 port map( B1 => n17641, B2 => n17398, C1 => n17638, C2 =>
                           n16934, A => n15010, ZN => n15005);
   U14072 : OAI22_X1 port map( A1 => n16577, A2 => n17635, B1 => n17117, B2 => 
                           n17632, ZN => n15010);
   U14073 : AOI221_X1 port map( B1 => n17689, B2 => n17399, C1 => n17686, C2 =>
                           n16935, A => n14983, ZN => n14978);
   U14074 : OAI22_X1 port map( A1 => n16614, A2 => n17683, B1 => n17190, B2 => 
                           n17680, ZN => n14983);
   U14075 : AOI221_X1 port map( B1 => n17641, B2 => n17400, C1 => n17638, C2 =>
                           n16936, A => n14991, ZN => n14986);
   U14076 : OAI22_X1 port map( A1 => n16578, A2 => n17635, B1 => n17118, B2 => 
                           n17632, ZN => n14991);
   U14077 : AOI221_X1 port map( B1 => n17689, B2 => n17401, C1 => n17686, C2 =>
                           n16937, A => n14964, ZN => n14959);
   U14078 : OAI22_X1 port map( A1 => n16615, A2 => n17683, B1 => n17191, B2 => 
                           n17680, ZN => n14964);
   U14079 : AOI221_X1 port map( B1 => n17641, B2 => n17402, C1 => n17638, C2 =>
                           n16938, A => n14972, ZN => n14967);
   U14080 : OAI22_X1 port map( A1 => n16579, A2 => n17635, B1 => n17119, B2 => 
                           n17632, ZN => n14972);
   U14081 : AOI221_X1 port map( B1 => n17689, B2 => n17403, C1 => n17686, C2 =>
                           n16939, A => n14945, ZN => n14940);
   U14082 : OAI22_X1 port map( A1 => n16616, A2 => n17683, B1 => n17192, B2 => 
                           n17680, ZN => n14945);
   U14083 : AOI221_X1 port map( B1 => n17641, B2 => n17404, C1 => n17638, C2 =>
                           n16940, A => n14953, ZN => n14948);
   U14084 : OAI22_X1 port map( A1 => n16580, A2 => n17635, B1 => n17120, B2 => 
                           n17632, ZN => n14953);
   U14085 : AOI221_X1 port map( B1 => n17689, B2 => n17405, C1 => n17686, C2 =>
                           n16941, A => n14926, ZN => n14921);
   U14086 : OAI22_X1 port map( A1 => n16617, A2 => n17683, B1 => n17193, B2 => 
                           n17680, ZN => n14926);
   U14087 : AOI221_X1 port map( B1 => n17641, B2 => n17406, C1 => n17638, C2 =>
                           n16942, A => n14934, ZN => n14929);
   U14088 : OAI22_X1 port map( A1 => n16581, A2 => n17635, B1 => n17121, B2 => 
                           n17632, ZN => n14934);
   U14089 : AOI221_X1 port map( B1 => n17689, B2 => n17407, C1 => n17686, C2 =>
                           n16943, A => n14907, ZN => n14902);
   U14090 : OAI22_X1 port map( A1 => n16618, A2 => n17683, B1 => n17194, B2 => 
                           n17680, ZN => n14907);
   U14091 : AOI221_X1 port map( B1 => n17641, B2 => n17408, C1 => n17638, C2 =>
                           n16944, A => n14915, ZN => n14910);
   U14092 : OAI22_X1 port map( A1 => n16582, A2 => n17635, B1 => n17122, B2 => 
                           n17632, ZN => n14915);
   U14093 : AOI221_X1 port map( B1 => n17689, B2 => n17409, C1 => n17686, C2 =>
                           n16945, A => n14888, ZN => n14883);
   U14094 : OAI22_X1 port map( A1 => n16619, A2 => n17683, B1 => n17195, B2 => 
                           n17680, ZN => n14888);
   U14095 : AOI221_X1 port map( B1 => n17641, B2 => n17410, C1 => n17638, C2 =>
                           n16946, A => n14896, ZN => n14891);
   U14096 : OAI22_X1 port map( A1 => n16583, A2 => n17635, B1 => n17123, B2 => 
                           n17632, ZN => n14896);
   U14097 : AOI221_X1 port map( B1 => n17689, B2 => n17411, C1 => n17686, C2 =>
                           n16947, A => n14869, ZN => n14864);
   U14098 : OAI22_X1 port map( A1 => n16620, A2 => n17683, B1 => n17196, B2 => 
                           n17680, ZN => n14869);
   U14099 : AOI221_X1 port map( B1 => n17641, B2 => n17412, C1 => n17638, C2 =>
                           n16948, A => n14877, ZN => n14872);
   U14100 : OAI22_X1 port map( A1 => n16584, A2 => n17635, B1 => n17124, B2 => 
                           n17632, ZN => n14877);
   U14101 : AOI221_X1 port map( B1 => n17690, B2 => n17413, C1 => n17687, C2 =>
                           n16949, A => n14850, ZN => n14845);
   U14102 : OAI22_X1 port map( A1 => n16533, A2 => n17684, B1 => n16789, B2 => 
                           n17681, ZN => n14850);
   U14103 : AOI221_X1 port map( B1 => n17642, B2 => n17414, C1 => n17639, C2 =>
                           n16950, A => n14858, ZN => n14853);
   U14104 : OAI22_X1 port map( A1 => n16509, A2 => n17636, B1 => n16765, B2 => 
                           n17633, ZN => n14858);
   U14105 : AOI221_X1 port map( B1 => n17690, B2 => n17415, C1 => n17687, C2 =>
                           n16951, A => n14831, ZN => n14826);
   U14106 : OAI22_X1 port map( A1 => n16534, A2 => n17684, B1 => n16790, B2 => 
                           n17681, ZN => n14831);
   U14107 : AOI221_X1 port map( B1 => n17642, B2 => n17416, C1 => n17639, C2 =>
                           n16952, A => n14839, ZN => n14834);
   U14108 : OAI22_X1 port map( A1 => n16510, A2 => n17636, B1 => n16766, B2 => 
                           n17633, ZN => n14839);
   U14109 : AOI221_X1 port map( B1 => n17690, B2 => n17417, C1 => n17687, C2 =>
                           n16953, A => n14812, ZN => n14807);
   U14110 : OAI22_X1 port map( A1 => n16535, A2 => n17684, B1 => n16791, B2 => 
                           n17681, ZN => n14812);
   U14111 : AOI221_X1 port map( B1 => n17642, B2 => n17418, C1 => n17639, C2 =>
                           n16954, A => n14820, ZN => n14815);
   U14112 : OAI22_X1 port map( A1 => n16511, A2 => n17636, B1 => n16767, B2 => 
                           n17633, ZN => n14820);
   U14113 : AOI221_X1 port map( B1 => n17690, B2 => n17419, C1 => n17687, C2 =>
                           n16955, A => n14793, ZN => n14788);
   U14114 : OAI22_X1 port map( A1 => n16536, A2 => n17684, B1 => n16792, B2 => 
                           n17681, ZN => n14793);
   U14115 : AOI221_X1 port map( B1 => n17642, B2 => n17420, C1 => n17639, C2 =>
                           n16956, A => n14801, ZN => n14796);
   U14116 : OAI22_X1 port map( A1 => n16512, A2 => n17636, B1 => n16768, B2 => 
                           n17633, ZN => n14801);
   U14117 : AOI221_X1 port map( B1 => n17690, B2 => n17421, C1 => n17687, C2 =>
                           n16957, A => n14774, ZN => n14769);
   U14118 : OAI22_X1 port map( A1 => n16537, A2 => n17684, B1 => n16793, B2 => 
                           n17681, ZN => n14774);
   U14119 : AOI221_X1 port map( B1 => n17642, B2 => n17422, C1 => n17639, C2 =>
                           n16958, A => n14782, ZN => n14777);
   U14120 : OAI22_X1 port map( A1 => n16513, A2 => n17636, B1 => n16769, B2 => 
                           n17633, ZN => n14782);
   U14121 : AOI221_X1 port map( B1 => n17690, B2 => n17423, C1 => n17687, C2 =>
                           n16959, A => n14755, ZN => n14750);
   U14122 : OAI22_X1 port map( A1 => n16538, A2 => n17684, B1 => n16794, B2 => 
                           n17681, ZN => n14755);
   U14123 : AOI221_X1 port map( B1 => n17642, B2 => n17424, C1 => n17639, C2 =>
                           n16960, A => n14763, ZN => n14758);
   U14124 : OAI22_X1 port map( A1 => n16514, A2 => n17636, B1 => n16770, B2 => 
                           n17633, ZN => n14763);
   U14125 : AOI221_X1 port map( B1 => n17690, B2 => n17425, C1 => n17687, C2 =>
                           n16961, A => n14736, ZN => n14731);
   U14126 : OAI22_X1 port map( A1 => n16539, A2 => n17684, B1 => n16795, B2 => 
                           n17681, ZN => n14736);
   U14127 : AOI221_X1 port map( B1 => n17642, B2 => n17426, C1 => n17639, C2 =>
                           n16962, A => n14744, ZN => n14739);
   U14128 : OAI22_X1 port map( A1 => n16515, A2 => n17636, B1 => n16771, B2 => 
                           n17633, ZN => n14744);
   U14129 : AOI221_X1 port map( B1 => n17690, B2 => n17427, C1 => n17687, C2 =>
                           n16963, A => n14695, ZN => n14680);
   U14130 : OAI22_X1 port map( A1 => n16540, A2 => n17684, B1 => n16796, B2 => 
                           n17681, ZN => n14695);
   U14131 : AOI221_X1 port map( B1 => n17642, B2 => n17428, C1 => n17639, C2 =>
                           n16964, A => n14719, ZN => n14704);
   U14132 : OAI22_X1 port map( A1 => n16516, A2 => n17636, B1 => n16772, B2 => 
                           n17633, ZN => n14719);
   U14133 : AOI221_X1 port map( B1 => n17574, B2 => n17245, C1 => n17571, C2 =>
                           n16965, A => n15968, ZN => n15953);
   U14134 : OAI22_X1 port map( A1 => n16725, A2 => n17568, B1 => n17197, B2 => 
                           n17565, ZN => n15968);
   U14135 : AOI221_X1 port map( B1 => n17526, B2 => n17429, C1 => n17523, C2 =>
                           n16966, A => n15980, ZN => n15969);
   U14136 : OAI22_X1 port map( A1 => n16689, A2 => n17520, B1 => n17125, B2 => 
                           n17517, ZN => n15980);
   U14137 : AOI221_X1 port map( B1 => n17574, B2 => n17246, C1 => n17571, C2 =>
                           n16967, A => n15941, ZN => n15934);
   U14138 : OAI22_X1 port map( A1 => n16726, A2 => n17568, B1 => n17198, B2 => 
                           n17565, ZN => n15941);
   U14139 : AOI221_X1 port map( B1 => n17526, B2 => n17430, C1 => n17523, C2 =>
                           n16968, A => n15949, ZN => n15942);
   U14140 : OAI22_X1 port map( A1 => n16690, A2 => n17520, B1 => n17126, B2 => 
                           n17517, ZN => n15949);
   U14141 : AOI221_X1 port map( B1 => n17574, B2 => n17247, C1 => n17571, C2 =>
                           n16969, A => n15922, ZN => n15915);
   U14142 : OAI22_X1 port map( A1 => n16727, A2 => n17568, B1 => n17199, B2 => 
                           n17565, ZN => n15922);
   U14143 : AOI221_X1 port map( B1 => n17526, B2 => n17431, C1 => n17523, C2 =>
                           n16970, A => n15930, ZN => n15923);
   U14144 : OAI22_X1 port map( A1 => n16691, A2 => n17520, B1 => n17127, B2 => 
                           n17517, ZN => n15930);
   U14145 : AOI221_X1 port map( B1 => n17574, B2 => n17248, C1 => n17571, C2 =>
                           n16971, A => n15903, ZN => n15896);
   U14146 : OAI22_X1 port map( A1 => n16728, A2 => n17568, B1 => n17200, B2 => 
                           n17565, ZN => n15903);
   U14147 : AOI221_X1 port map( B1 => n17526, B2 => n17432, C1 => n17523, C2 =>
                           n16972, A => n15911, ZN => n15904);
   U14148 : OAI22_X1 port map( A1 => n16692, A2 => n17520, B1 => n17128, B2 => 
                           n17517, ZN => n15911);
   U14149 : AOI221_X1 port map( B1 => n17574, B2 => n17249, C1 => n17571, C2 =>
                           n16973, A => n15884, ZN => n15877);
   U14150 : OAI22_X1 port map( A1 => n16729, A2 => n17568, B1 => n17201, B2 => 
                           n17565, ZN => n15884);
   U14151 : AOI221_X1 port map( B1 => n17526, B2 => n17433, C1 => n17523, C2 =>
                           n16974, A => n15892, ZN => n15885);
   U14152 : OAI22_X1 port map( A1 => n16693, A2 => n17520, B1 => n17129, B2 => 
                           n17517, ZN => n15892);
   U14153 : AOI221_X1 port map( B1 => n17574, B2 => n17250, C1 => n17571, C2 =>
                           n16975, A => n15865, ZN => n15858);
   U14154 : OAI22_X1 port map( A1 => n16730, A2 => n17568, B1 => n17202, B2 => 
                           n17565, ZN => n15865);
   U14155 : AOI221_X1 port map( B1 => n17526, B2 => n17434, C1 => n17523, C2 =>
                           n16976, A => n15873, ZN => n15866);
   U14156 : OAI22_X1 port map( A1 => n16694, A2 => n17520, B1 => n17130, B2 => 
                           n17517, ZN => n15873);
   U14157 : AOI221_X1 port map( B1 => n17574, B2 => n17251, C1 => n17571, C2 =>
                           n16977, A => n15846, ZN => n15839);
   U14158 : OAI22_X1 port map( A1 => n16731, A2 => n17568, B1 => n17203, B2 => 
                           n17565, ZN => n15846);
   U14159 : AOI221_X1 port map( B1 => n17526, B2 => n17435, C1 => n17523, C2 =>
                           n16978, A => n15854, ZN => n15847);
   U14160 : OAI22_X1 port map( A1 => n16695, A2 => n17520, B1 => n17131, B2 => 
                           n17517, ZN => n15854);
   U14161 : AOI221_X1 port map( B1 => n17574, B2 => n17252, C1 => n17571, C2 =>
                           n16979, A => n15827, ZN => n15820);
   U14162 : OAI22_X1 port map( A1 => n16732, A2 => n17568, B1 => n17204, B2 => 
                           n17565, ZN => n15827);
   U14163 : AOI221_X1 port map( B1 => n17526, B2 => n17436, C1 => n17523, C2 =>
                           n16980, A => n15835, ZN => n15828);
   U14164 : OAI22_X1 port map( A1 => n16696, A2 => n17520, B1 => n17132, B2 => 
                           n17517, ZN => n15835);
   U14165 : AOI221_X1 port map( B1 => n17574, B2 => n17253, C1 => n17571, C2 =>
                           n16981, A => n15808, ZN => n15801);
   U14166 : OAI22_X1 port map( A1 => n16733, A2 => n17568, B1 => n17205, B2 => 
                           n17565, ZN => n15808);
   U14167 : AOI221_X1 port map( B1 => n17526, B2 => n17437, C1 => n17523, C2 =>
                           n16982, A => n15816, ZN => n15809);
   U14168 : OAI22_X1 port map( A1 => n16697, A2 => n17520, B1 => n17133, B2 => 
                           n17517, ZN => n15816);
   U14169 : AOI221_X1 port map( B1 => n17574, B2 => n17254, C1 => n17571, C2 =>
                           n16983, A => n15789, ZN => n15782);
   U14170 : OAI22_X1 port map( A1 => n16734, A2 => n17568, B1 => n17206, B2 => 
                           n17565, ZN => n15789);
   U14171 : AOI221_X1 port map( B1 => n17526, B2 => n17438, C1 => n17523, C2 =>
                           n16984, A => n15797, ZN => n15790);
   U14172 : OAI22_X1 port map( A1 => n16698, A2 => n17520, B1 => n17134, B2 => 
                           n17517, ZN => n15797);
   U14173 : AOI221_X1 port map( B1 => n17574, B2 => n17255, C1 => n17571, C2 =>
                           n16985, A => n15770, ZN => n15763);
   U14174 : OAI22_X1 port map( A1 => n16735, A2 => n17568, B1 => n17207, B2 => 
                           n17565, ZN => n15770);
   U14175 : AOI221_X1 port map( B1 => n17526, B2 => n17439, C1 => n17523, C2 =>
                           n16986, A => n15778, ZN => n15771);
   U14176 : OAI22_X1 port map( A1 => n16699, A2 => n17520, B1 => n17135, B2 => 
                           n17517, ZN => n15778);
   U14177 : AOI221_X1 port map( B1 => n17574, B2 => n17256, C1 => n17571, C2 =>
                           n16987, A => n15751, ZN => n15744);
   U14178 : OAI22_X1 port map( A1 => n16736, A2 => n17568, B1 => n17208, B2 => 
                           n17565, ZN => n15751);
   U14179 : AOI221_X1 port map( B1 => n17526, B2 => n17440, C1 => n17523, C2 =>
                           n16988, A => n15759, ZN => n15752);
   U14180 : OAI22_X1 port map( A1 => n16700, A2 => n17520, B1 => n17136, B2 => 
                           n17517, ZN => n15759);
   U14181 : AOI221_X1 port map( B1 => n17575, B2 => n17257, C1 => n17572, C2 =>
                           n16989, A => n15732, ZN => n15725);
   U14182 : OAI22_X1 port map( A1 => n16621, A2 => n17569, B1 => n17209, B2 => 
                           n17566, ZN => n15732);
   U14183 : AOI221_X1 port map( B1 => n17527, B2 => n17441, C1 => n17524, C2 =>
                           n16990, A => n15740, ZN => n15733);
   U14184 : OAI22_X1 port map( A1 => n16585, A2 => n17521, B1 => n17137, B2 => 
                           n17518, ZN => n15740);
   U14185 : AOI221_X1 port map( B1 => n17575, B2 => n17258, C1 => n17572, C2 =>
                           n16991, A => n15713, ZN => n15706);
   U14186 : OAI22_X1 port map( A1 => n16622, A2 => n17569, B1 => n17210, B2 => 
                           n17566, ZN => n15713);
   U14187 : AOI221_X1 port map( B1 => n17527, B2 => n17442, C1 => n17524, C2 =>
                           n16992, A => n15721, ZN => n15714);
   U14188 : OAI22_X1 port map( A1 => n16586, A2 => n17521, B1 => n17138, B2 => 
                           n17518, ZN => n15721);
   U14189 : AOI221_X1 port map( B1 => n17575, B2 => n17259, C1 => n17572, C2 =>
                           n16993, A => n15694, ZN => n15687);
   U14190 : OAI22_X1 port map( A1 => n16623, A2 => n17569, B1 => n17211, B2 => 
                           n17566, ZN => n15694);
   U14191 : AOI221_X1 port map( B1 => n17527, B2 => n17443, C1 => n17524, C2 =>
                           n16994, A => n15702, ZN => n15695);
   U14192 : OAI22_X1 port map( A1 => n16587, A2 => n17521, B1 => n17139, B2 => 
                           n17518, ZN => n15702);
   U14193 : AOI221_X1 port map( B1 => n17575, B2 => n17260, C1 => n17572, C2 =>
                           n16995, A => n15675, ZN => n15668);
   U14194 : OAI22_X1 port map( A1 => n16624, A2 => n17569, B1 => n17212, B2 => 
                           n17566, ZN => n15675);
   U14195 : AOI221_X1 port map( B1 => n17527, B2 => n17444, C1 => n17524, C2 =>
                           n16996, A => n15683, ZN => n15676);
   U14196 : OAI22_X1 port map( A1 => n16588, A2 => n17521, B1 => n17140, B2 => 
                           n17518, ZN => n15683);
   U14197 : AOI221_X1 port map( B1 => n17575, B2 => n17261, C1 => n17572, C2 =>
                           n16997, A => n15656, ZN => n15649);
   U14198 : OAI22_X1 port map( A1 => n16625, A2 => n17569, B1 => n17213, B2 => 
                           n17566, ZN => n15656);
   U14199 : AOI221_X1 port map( B1 => n17527, B2 => n17445, C1 => n17524, C2 =>
                           n16998, A => n15664, ZN => n15657);
   U14200 : OAI22_X1 port map( A1 => n16589, A2 => n17521, B1 => n17141, B2 => 
                           n17518, ZN => n15664);
   U14201 : AOI221_X1 port map( B1 => n17575, B2 => n17262, C1 => n17572, C2 =>
                           n16999, A => n15637, ZN => n15630);
   U14202 : OAI22_X1 port map( A1 => n16626, A2 => n17569, B1 => n17214, B2 => 
                           n17566, ZN => n15637);
   U14203 : AOI221_X1 port map( B1 => n17527, B2 => n17446, C1 => n17524, C2 =>
                           n17000, A => n15645, ZN => n15638);
   U14204 : OAI22_X1 port map( A1 => n16590, A2 => n17521, B1 => n17142, B2 => 
                           n17518, ZN => n15645);
   U14205 : AOI221_X1 port map( B1 => n17575, B2 => n17263, C1 => n17572, C2 =>
                           n17001, A => n15618, ZN => n15611);
   U14206 : OAI22_X1 port map( A1 => n16627, A2 => n17569, B1 => n17215, B2 => 
                           n17566, ZN => n15618);
   U14207 : AOI221_X1 port map( B1 => n17527, B2 => n17447, C1 => n17524, C2 =>
                           n17002, A => n15626, ZN => n15619);
   U14208 : OAI22_X1 port map( A1 => n16591, A2 => n17521, B1 => n17143, B2 => 
                           n17518, ZN => n15626);
   U14209 : AOI221_X1 port map( B1 => n17575, B2 => n17264, C1 => n17572, C2 =>
                           n17003, A => n15599, ZN => n15592);
   U14210 : OAI22_X1 port map( A1 => n16628, A2 => n17569, B1 => n17216, B2 => 
                           n17566, ZN => n15599);
   U14211 : AOI221_X1 port map( B1 => n17527, B2 => n17448, C1 => n17524, C2 =>
                           n17004, A => n15607, ZN => n15600);
   U14212 : OAI22_X1 port map( A1 => n16592, A2 => n17521, B1 => n17144, B2 => 
                           n17518, ZN => n15607);
   U14213 : AOI221_X1 port map( B1 => n17575, B2 => n17265, C1 => n17572, C2 =>
                           n17005, A => n15580, ZN => n15573);
   U14214 : OAI22_X1 port map( A1 => n16629, A2 => n17569, B1 => n17217, B2 => 
                           n17566, ZN => n15580);
   U14215 : AOI221_X1 port map( B1 => n17527, B2 => n17449, C1 => n17524, C2 =>
                           n17006, A => n15588, ZN => n15581);
   U14216 : OAI22_X1 port map( A1 => n16593, A2 => n17521, B1 => n17145, B2 => 
                           n17518, ZN => n15588);
   U14217 : AOI221_X1 port map( B1 => n17575, B2 => n17266, C1 => n17572, C2 =>
                           n17007, A => n15561, ZN => n15554);
   U14218 : OAI22_X1 port map( A1 => n16630, A2 => n17569, B1 => n17218, B2 => 
                           n17566, ZN => n15561);
   U14219 : AOI221_X1 port map( B1 => n17527, B2 => n17450, C1 => n17524, C2 =>
                           n17008, A => n15569, ZN => n15562);
   U14220 : OAI22_X1 port map( A1 => n16594, A2 => n17521, B1 => n17146, B2 => 
                           n17518, ZN => n15569);
   U14221 : AOI221_X1 port map( B1 => n17575, B2 => n17267, C1 => n17572, C2 =>
                           n17009, A => n15542, ZN => n15535);
   U14222 : OAI22_X1 port map( A1 => n16631, A2 => n17569, B1 => n17219, B2 => 
                           n17566, ZN => n15542);
   U14223 : AOI221_X1 port map( B1 => n17527, B2 => n17451, C1 => n17524, C2 =>
                           n17010, A => n15550, ZN => n15543);
   U14224 : OAI22_X1 port map( A1 => n16595, A2 => n17521, B1 => n17147, B2 => 
                           n17518, ZN => n15550);
   U14225 : AOI221_X1 port map( B1 => n17575, B2 => n17268, C1 => n17572, C2 =>
                           n17011, A => n15523, ZN => n15516);
   U14226 : OAI22_X1 port map( A1 => n16632, A2 => n17569, B1 => n17220, B2 => 
                           n17566, ZN => n15523);
   U14227 : AOI221_X1 port map( B1 => n17527, B2 => n17452, C1 => n17524, C2 =>
                           n17012, A => n15531, ZN => n15524);
   U14228 : OAI22_X1 port map( A1 => n16596, A2 => n17521, B1 => n17148, B2 => 
                           n17518, ZN => n15531);
   U14229 : AOI221_X1 port map( B1 => n17576, B2 => n17269, C1 => n17573, C2 =>
                           n17013, A => n15504, ZN => n15497);
   U14230 : OAI22_X1 port map( A1 => n16541, A2 => n17570, B1 => n16797, B2 => 
                           n17567, ZN => n15504);
   U14231 : AOI221_X1 port map( B1 => n17528, B2 => n17453, C1 => n17525, C2 =>
                           n17014, A => n15512, ZN => n15505);
   U14232 : OAI22_X1 port map( A1 => n16517, A2 => n17522, B1 => n16773, B2 => 
                           n17519, ZN => n15512);
   U14233 : AOI221_X1 port map( B1 => n17576, B2 => n17270, C1 => n17573, C2 =>
                           n17015, A => n15485, ZN => n15478);
   U14234 : OAI22_X1 port map( A1 => n16542, A2 => n17570, B1 => n16798, B2 => 
                           n17567, ZN => n15485);
   U14235 : AOI221_X1 port map( B1 => n17528, B2 => n17454, C1 => n17525, C2 =>
                           n17016, A => n15493, ZN => n15486);
   U14236 : OAI22_X1 port map( A1 => n16518, A2 => n17522, B1 => n16774, B2 => 
                           n17519, ZN => n15493);
   U14237 : AOI221_X1 port map( B1 => n17576, B2 => n17271, C1 => n17573, C2 =>
                           n17017, A => n15466, ZN => n15459);
   U14238 : OAI22_X1 port map( A1 => n16543, A2 => n17570, B1 => n16799, B2 => 
                           n17567, ZN => n15466);
   U14239 : AOI221_X1 port map( B1 => n17528, B2 => n17455, C1 => n17525, C2 =>
                           n17018, A => n15474, ZN => n15467);
   U14240 : OAI22_X1 port map( A1 => n16519, A2 => n17522, B1 => n16775, B2 => 
                           n17519, ZN => n15474);
   U14241 : AOI221_X1 port map( B1 => n17576, B2 => n17272, C1 => n17573, C2 =>
                           n17019, A => n15447, ZN => n15440);
   U14242 : OAI22_X1 port map( A1 => n16544, A2 => n17570, B1 => n16800, B2 => 
                           n17567, ZN => n15447);
   U14243 : AOI221_X1 port map( B1 => n17528, B2 => n17456, C1 => n17525, C2 =>
                           n17020, A => n15455, ZN => n15448);
   U14244 : OAI22_X1 port map( A1 => n16520, A2 => n17522, B1 => n16776, B2 => 
                           n17519, ZN => n15455);
   U14245 : AOI221_X1 port map( B1 => n17576, B2 => n17273, C1 => n17573, C2 =>
                           n17021, A => n15428, ZN => n15421);
   U14246 : OAI22_X1 port map( A1 => n16545, A2 => n17570, B1 => n16801, B2 => 
                           n17567, ZN => n15428);
   U14247 : AOI221_X1 port map( B1 => n17528, B2 => n17457, C1 => n17525, C2 =>
                           n17022, A => n15436, ZN => n15429);
   U14248 : OAI22_X1 port map( A1 => n16521, A2 => n17522, B1 => n16777, B2 => 
                           n17519, ZN => n15436);
   U14249 : AOI221_X1 port map( B1 => n17576, B2 => n17274, C1 => n17573, C2 =>
                           n17023, A => n15409, ZN => n15402);
   U14250 : OAI22_X1 port map( A1 => n16546, A2 => n17570, B1 => n16802, B2 => 
                           n17567, ZN => n15409);
   U14251 : AOI221_X1 port map( B1 => n17528, B2 => n17458, C1 => n17525, C2 =>
                           n17024, A => n15417, ZN => n15410);
   U14252 : OAI22_X1 port map( A1 => n16522, A2 => n17522, B1 => n16778, B2 => 
                           n17519, ZN => n15417);
   U14253 : AOI221_X1 port map( B1 => n17576, B2 => n17275, C1 => n17573, C2 =>
                           n17025, A => n15390, ZN => n15383);
   U14254 : OAI22_X1 port map( A1 => n16547, A2 => n17570, B1 => n16803, B2 => 
                           n17567, ZN => n15390);
   U14255 : AOI221_X1 port map( B1 => n17528, B2 => n17459, C1 => n17525, C2 =>
                           n17026, A => n15398, ZN => n15391);
   U14256 : OAI22_X1 port map( A1 => n16523, A2 => n17522, B1 => n16779, B2 => 
                           n17519, ZN => n15398);
   U14257 : AOI221_X1 port map( B1 => n17576, B2 => n17276, C1 => n17573, C2 =>
                           n17027, A => n15353, ZN => n15332);
   U14258 : OAI22_X1 port map( A1 => n16548, A2 => n17570, B1 => n16804, B2 => 
                           n17567, ZN => n15353);
   U14259 : AOI221_X1 port map( B1 => n17528, B2 => n17460, C1 => n17525, C2 =>
                           n17028, A => n15377, ZN => n15356);
   U14260 : OAI22_X1 port map( A1 => n16524, A2 => n17522, B1 => n16780, B2 => 
                           n17519, ZN => n15377);
   U14261 : AOI221_X1 port map( B1 => n17676, B2 => n17245, C1 => n17673, C2 =>
                           n16965, A => n15315, ZN => n15300);
   U14262 : OAI22_X1 port map( A1 => n16725, A2 => n17670, B1 => n17197, B2 => 
                           n17667, ZN => n15315);
   U14263 : AOI221_X1 port map( B1 => n17628, B2 => n17429, C1 => n17625, C2 =>
                           n16966, A => n15327, ZN => n15316);
   U14264 : OAI22_X1 port map( A1 => n16689, A2 => n17622, B1 => n17125, B2 => 
                           n17619, ZN => n15327);
   U14265 : AOI221_X1 port map( B1 => n17676, B2 => n17246, C1 => n17673, C2 =>
                           n16967, A => n15288, ZN => n15281);
   U14266 : OAI22_X1 port map( A1 => n16726, A2 => n17670, B1 => n17198, B2 => 
                           n17667, ZN => n15288);
   U14267 : AOI221_X1 port map( B1 => n17628, B2 => n17430, C1 => n17625, C2 =>
                           n16968, A => n15296, ZN => n15289);
   U14268 : OAI22_X1 port map( A1 => n16690, A2 => n17622, B1 => n17126, B2 => 
                           n17619, ZN => n15296);
   U14269 : AOI221_X1 port map( B1 => n17676, B2 => n17247, C1 => n17673, C2 =>
                           n16969, A => n15269, ZN => n15262);
   U14270 : OAI22_X1 port map( A1 => n16727, A2 => n17670, B1 => n17199, B2 => 
                           n17667, ZN => n15269);
   U14271 : AOI221_X1 port map( B1 => n17628, B2 => n17431, C1 => n17625, C2 =>
                           n16970, A => n15277, ZN => n15270);
   U14272 : OAI22_X1 port map( A1 => n16691, A2 => n17622, B1 => n17127, B2 => 
                           n17619, ZN => n15277);
   U14273 : AOI221_X1 port map( B1 => n17676, B2 => n17248, C1 => n17673, C2 =>
                           n16971, A => n15250, ZN => n15243);
   U14274 : OAI22_X1 port map( A1 => n16728, A2 => n17670, B1 => n17200, B2 => 
                           n17667, ZN => n15250);
   U14275 : AOI221_X1 port map( B1 => n17628, B2 => n17432, C1 => n17625, C2 =>
                           n16972, A => n15258, ZN => n15251);
   U14276 : OAI22_X1 port map( A1 => n16692, A2 => n17622, B1 => n17128, B2 => 
                           n17619, ZN => n15258);
   U14277 : AOI221_X1 port map( B1 => n17676, B2 => n17249, C1 => n17673, C2 =>
                           n16973, A => n15231, ZN => n15224);
   U14278 : OAI22_X1 port map( A1 => n16729, A2 => n17670, B1 => n17201, B2 => 
                           n17667, ZN => n15231);
   U14279 : AOI221_X1 port map( B1 => n17628, B2 => n17433, C1 => n17625, C2 =>
                           n16974, A => n15239, ZN => n15232);
   U14280 : OAI22_X1 port map( A1 => n16693, A2 => n17622, B1 => n17129, B2 => 
                           n17619, ZN => n15239);
   U14281 : AOI221_X1 port map( B1 => n17676, B2 => n17250, C1 => n17673, C2 =>
                           n16975, A => n15212, ZN => n15205);
   U14282 : OAI22_X1 port map( A1 => n16730, A2 => n17670, B1 => n17202, B2 => 
                           n17667, ZN => n15212);
   U14283 : AOI221_X1 port map( B1 => n17628, B2 => n17434, C1 => n17625, C2 =>
                           n16976, A => n15220, ZN => n15213);
   U14284 : OAI22_X1 port map( A1 => n16694, A2 => n17622, B1 => n17130, B2 => 
                           n17619, ZN => n15220);
   U14285 : AOI221_X1 port map( B1 => n17676, B2 => n17251, C1 => n17673, C2 =>
                           n16977, A => n15193, ZN => n15186);
   U14286 : OAI22_X1 port map( A1 => n16731, A2 => n17670, B1 => n17203, B2 => 
                           n17667, ZN => n15193);
   U14287 : AOI221_X1 port map( B1 => n17628, B2 => n17435, C1 => n17625, C2 =>
                           n16978, A => n15201, ZN => n15194);
   U14288 : OAI22_X1 port map( A1 => n16695, A2 => n17622, B1 => n17131, B2 => 
                           n17619, ZN => n15201);
   U14289 : AOI221_X1 port map( B1 => n17676, B2 => n17252, C1 => n17673, C2 =>
                           n16979, A => n15174, ZN => n15167);
   U14290 : OAI22_X1 port map( A1 => n16732, A2 => n17670, B1 => n17204, B2 => 
                           n17667, ZN => n15174);
   U14291 : AOI221_X1 port map( B1 => n17628, B2 => n17436, C1 => n17625, C2 =>
                           n16980, A => n15182, ZN => n15175);
   U14292 : OAI22_X1 port map( A1 => n16696, A2 => n17622, B1 => n17132, B2 => 
                           n17619, ZN => n15182);
   U14293 : AOI221_X1 port map( B1 => n17676, B2 => n17253, C1 => n17673, C2 =>
                           n16981, A => n15155, ZN => n15148);
   U14294 : OAI22_X1 port map( A1 => n16733, A2 => n17670, B1 => n17205, B2 => 
                           n17667, ZN => n15155);
   U14295 : AOI221_X1 port map( B1 => n17628, B2 => n17437, C1 => n17625, C2 =>
                           n16982, A => n15163, ZN => n15156);
   U14296 : OAI22_X1 port map( A1 => n16697, A2 => n17622, B1 => n17133, B2 => 
                           n17619, ZN => n15163);
   U14297 : AOI221_X1 port map( B1 => n17676, B2 => n17254, C1 => n17673, C2 =>
                           n16983, A => n15136, ZN => n15129);
   U14298 : OAI22_X1 port map( A1 => n16734, A2 => n17670, B1 => n17206, B2 => 
                           n17667, ZN => n15136);
   U14299 : AOI221_X1 port map( B1 => n17628, B2 => n17438, C1 => n17625, C2 =>
                           n16984, A => n15144, ZN => n15137);
   U14300 : OAI22_X1 port map( A1 => n16698, A2 => n17622, B1 => n17134, B2 => 
                           n17619, ZN => n15144);
   U14301 : AOI221_X1 port map( B1 => n17676, B2 => n17255, C1 => n17673, C2 =>
                           n16985, A => n15117, ZN => n15110);
   U14302 : OAI22_X1 port map( A1 => n16735, A2 => n17670, B1 => n17207, B2 => 
                           n17667, ZN => n15117);
   U14303 : AOI221_X1 port map( B1 => n17628, B2 => n17439, C1 => n17625, C2 =>
                           n16986, A => n15125, ZN => n15118);
   U14304 : OAI22_X1 port map( A1 => n16699, A2 => n17622, B1 => n17135, B2 => 
                           n17619, ZN => n15125);
   U14305 : AOI221_X1 port map( B1 => n17676, B2 => n17256, C1 => n17673, C2 =>
                           n16987, A => n15098, ZN => n15091);
   U14306 : OAI22_X1 port map( A1 => n16736, A2 => n17670, B1 => n17208, B2 => 
                           n17667, ZN => n15098);
   U14307 : AOI221_X1 port map( B1 => n17628, B2 => n17440, C1 => n17625, C2 =>
                           n16988, A => n15106, ZN => n15099);
   U14308 : OAI22_X1 port map( A1 => n16700, A2 => n17622, B1 => n17136, B2 => 
                           n17619, ZN => n15106);
   U14309 : AOI221_X1 port map( B1 => n17677, B2 => n17257, C1 => n17674, C2 =>
                           n16989, A => n15079, ZN => n15072);
   U14310 : OAI22_X1 port map( A1 => n16621, A2 => n17671, B1 => n17209, B2 => 
                           n17668, ZN => n15079);
   U14311 : AOI221_X1 port map( B1 => n17629, B2 => n17441, C1 => n17626, C2 =>
                           n16990, A => n15087, ZN => n15080);
   U14312 : OAI22_X1 port map( A1 => n16585, A2 => n17623, B1 => n17137, B2 => 
                           n17620, ZN => n15087);
   U14313 : AOI221_X1 port map( B1 => n17677, B2 => n17258, C1 => n17674, C2 =>
                           n16991, A => n15060, ZN => n15053);
   U14314 : OAI22_X1 port map( A1 => n16622, A2 => n17671, B1 => n17210, B2 => 
                           n17668, ZN => n15060);
   U14315 : AOI221_X1 port map( B1 => n17629, B2 => n17442, C1 => n17626, C2 =>
                           n16992, A => n15068, ZN => n15061);
   U14316 : OAI22_X1 port map( A1 => n16586, A2 => n17623, B1 => n17138, B2 => 
                           n17620, ZN => n15068);
   U14317 : AOI221_X1 port map( B1 => n17677, B2 => n17259, C1 => n17674, C2 =>
                           n16993, A => n15041, ZN => n15034);
   U14318 : OAI22_X1 port map( A1 => n16623, A2 => n17671, B1 => n17211, B2 => 
                           n17668, ZN => n15041);
   U14319 : AOI221_X1 port map( B1 => n17629, B2 => n17443, C1 => n17626, C2 =>
                           n16994, A => n15049, ZN => n15042);
   U14320 : OAI22_X1 port map( A1 => n16587, A2 => n17623, B1 => n17139, B2 => 
                           n17620, ZN => n15049);
   U14321 : AOI221_X1 port map( B1 => n17677, B2 => n17260, C1 => n17674, C2 =>
                           n16995, A => n15022, ZN => n15015);
   U14322 : OAI22_X1 port map( A1 => n16624, A2 => n17671, B1 => n17212, B2 => 
                           n17668, ZN => n15022);
   U14323 : AOI221_X1 port map( B1 => n17629, B2 => n17444, C1 => n17626, C2 =>
                           n16996, A => n15030, ZN => n15023);
   U14324 : OAI22_X1 port map( A1 => n16588, A2 => n17623, B1 => n17140, B2 => 
                           n17620, ZN => n15030);
   U14325 : AOI221_X1 port map( B1 => n17677, B2 => n17261, C1 => n17674, C2 =>
                           n16997, A => n15003, ZN => n14996);
   U14326 : OAI22_X1 port map( A1 => n16625, A2 => n17671, B1 => n17213, B2 => 
                           n17668, ZN => n15003);
   U14327 : AOI221_X1 port map( B1 => n17629, B2 => n17445, C1 => n17626, C2 =>
                           n16998, A => n15011, ZN => n15004);
   U14328 : OAI22_X1 port map( A1 => n16589, A2 => n17623, B1 => n17141, B2 => 
                           n17620, ZN => n15011);
   U14329 : AOI221_X1 port map( B1 => n17677, B2 => n17262, C1 => n17674, C2 =>
                           n16999, A => n14984, ZN => n14977);
   U14330 : OAI22_X1 port map( A1 => n16626, A2 => n17671, B1 => n17214, B2 => 
                           n17668, ZN => n14984);
   U14331 : AOI221_X1 port map( B1 => n17629, B2 => n17446, C1 => n17626, C2 =>
                           n17000, A => n14992, ZN => n14985);
   U14332 : OAI22_X1 port map( A1 => n16590, A2 => n17623, B1 => n17142, B2 => 
                           n17620, ZN => n14992);
   U14333 : AOI221_X1 port map( B1 => n17677, B2 => n17263, C1 => n17674, C2 =>
                           n17001, A => n14965, ZN => n14958);
   U14334 : OAI22_X1 port map( A1 => n16627, A2 => n17671, B1 => n17215, B2 => 
                           n17668, ZN => n14965);
   U14335 : AOI221_X1 port map( B1 => n17629, B2 => n17447, C1 => n17626, C2 =>
                           n17002, A => n14973, ZN => n14966);
   U14336 : OAI22_X1 port map( A1 => n16591, A2 => n17623, B1 => n17143, B2 => 
                           n17620, ZN => n14973);
   U14337 : AOI221_X1 port map( B1 => n17677, B2 => n17264, C1 => n17674, C2 =>
                           n17003, A => n14946, ZN => n14939);
   U14338 : OAI22_X1 port map( A1 => n16628, A2 => n17671, B1 => n17216, B2 => 
                           n17668, ZN => n14946);
   U14339 : AOI221_X1 port map( B1 => n17629, B2 => n17448, C1 => n17626, C2 =>
                           n17004, A => n14954, ZN => n14947);
   U14340 : OAI22_X1 port map( A1 => n16592, A2 => n17623, B1 => n17144, B2 => 
                           n17620, ZN => n14954);
   U14341 : AOI221_X1 port map( B1 => n17677, B2 => n17265, C1 => n17674, C2 =>
                           n17005, A => n14927, ZN => n14920);
   U14342 : OAI22_X1 port map( A1 => n16629, A2 => n17671, B1 => n17217, B2 => 
                           n17668, ZN => n14927);
   U14343 : AOI221_X1 port map( B1 => n17629, B2 => n17449, C1 => n17626, C2 =>
                           n17006, A => n14935, ZN => n14928);
   U14344 : OAI22_X1 port map( A1 => n16593, A2 => n17623, B1 => n17145, B2 => 
                           n17620, ZN => n14935);
   U14345 : AOI221_X1 port map( B1 => n17677, B2 => n17266, C1 => n17674, C2 =>
                           n17007, A => n14908, ZN => n14901);
   U14346 : OAI22_X1 port map( A1 => n16630, A2 => n17671, B1 => n17218, B2 => 
                           n17668, ZN => n14908);
   U14347 : AOI221_X1 port map( B1 => n17629, B2 => n17450, C1 => n17626, C2 =>
                           n17008, A => n14916, ZN => n14909);
   U14348 : OAI22_X1 port map( A1 => n16594, A2 => n17623, B1 => n17146, B2 => 
                           n17620, ZN => n14916);
   U14349 : AOI221_X1 port map( B1 => n17677, B2 => n17267, C1 => n17674, C2 =>
                           n17009, A => n14889, ZN => n14882);
   U14350 : OAI22_X1 port map( A1 => n16631, A2 => n17671, B1 => n17219, B2 => 
                           n17668, ZN => n14889);
   U14351 : AOI221_X1 port map( B1 => n17629, B2 => n17451, C1 => n17626, C2 =>
                           n17010, A => n14897, ZN => n14890);
   U14352 : OAI22_X1 port map( A1 => n16595, A2 => n17623, B1 => n17147, B2 => 
                           n17620, ZN => n14897);
   U14353 : AOI221_X1 port map( B1 => n17677, B2 => n17268, C1 => n17674, C2 =>
                           n17011, A => n14870, ZN => n14863);
   U14354 : OAI22_X1 port map( A1 => n16632, A2 => n17671, B1 => n17220, B2 => 
                           n17668, ZN => n14870);
   U14355 : AOI221_X1 port map( B1 => n17629, B2 => n17452, C1 => n17626, C2 =>
                           n17012, A => n14878, ZN => n14871);
   U14356 : OAI22_X1 port map( A1 => n16596, A2 => n17623, B1 => n17148, B2 => 
                           n17620, ZN => n14878);
   U14357 : AOI221_X1 port map( B1 => n17678, B2 => n17269, C1 => n17675, C2 =>
                           n17013, A => n14851, ZN => n14844);
   U14358 : OAI22_X1 port map( A1 => n16541, A2 => n17672, B1 => n16797, B2 => 
                           n17669, ZN => n14851);
   U14359 : AOI221_X1 port map( B1 => n17630, B2 => n17453, C1 => n17627, C2 =>
                           n17014, A => n14859, ZN => n14852);
   U14360 : OAI22_X1 port map( A1 => n16517, A2 => n17624, B1 => n16773, B2 => 
                           n17621, ZN => n14859);
   U14361 : AOI221_X1 port map( B1 => n17678, B2 => n17270, C1 => n17675, C2 =>
                           n17015, A => n14832, ZN => n14825);
   U14362 : OAI22_X1 port map( A1 => n16542, A2 => n17672, B1 => n16798, B2 => 
                           n17669, ZN => n14832);
   U14363 : AOI221_X1 port map( B1 => n17630, B2 => n17454, C1 => n17627, C2 =>
                           n17016, A => n14840, ZN => n14833);
   U14364 : OAI22_X1 port map( A1 => n16518, A2 => n17624, B1 => n16774, B2 => 
                           n17621, ZN => n14840);
   U14365 : AOI221_X1 port map( B1 => n17678, B2 => n17271, C1 => n17675, C2 =>
                           n17017, A => n14813, ZN => n14806);
   U14366 : OAI22_X1 port map( A1 => n16543, A2 => n17672, B1 => n16799, B2 => 
                           n17669, ZN => n14813);
   U14367 : AOI221_X1 port map( B1 => n17630, B2 => n17455, C1 => n17627, C2 =>
                           n17018, A => n14821, ZN => n14814);
   U14368 : OAI22_X1 port map( A1 => n16519, A2 => n17624, B1 => n16775, B2 => 
                           n17621, ZN => n14821);
   U14369 : AOI221_X1 port map( B1 => n17678, B2 => n17272, C1 => n17675, C2 =>
                           n17019, A => n14794, ZN => n14787);
   U14370 : OAI22_X1 port map( A1 => n16544, A2 => n17672, B1 => n16800, B2 => 
                           n17669, ZN => n14794);
   U14371 : AOI221_X1 port map( B1 => n17630, B2 => n17456, C1 => n17627, C2 =>
                           n17020, A => n14802, ZN => n14795);
   U14372 : OAI22_X1 port map( A1 => n16520, A2 => n17624, B1 => n16776, B2 => 
                           n17621, ZN => n14802);
   U14373 : AOI221_X1 port map( B1 => n17678, B2 => n17273, C1 => n17675, C2 =>
                           n17021, A => n14775, ZN => n14768);
   U14374 : OAI22_X1 port map( A1 => n16545, A2 => n17672, B1 => n16801, B2 => 
                           n17669, ZN => n14775);
   U14375 : AOI221_X1 port map( B1 => n17630, B2 => n17457, C1 => n17627, C2 =>
                           n17022, A => n14783, ZN => n14776);
   U14376 : OAI22_X1 port map( A1 => n16521, A2 => n17624, B1 => n16777, B2 => 
                           n17621, ZN => n14783);
   U14377 : AOI221_X1 port map( B1 => n17678, B2 => n17274, C1 => n17675, C2 =>
                           n17023, A => n14756, ZN => n14749);
   U14378 : OAI22_X1 port map( A1 => n16546, A2 => n17672, B1 => n16802, B2 => 
                           n17669, ZN => n14756);
   U14379 : AOI221_X1 port map( B1 => n17630, B2 => n17458, C1 => n17627, C2 =>
                           n17024, A => n14764, ZN => n14757);
   U14380 : OAI22_X1 port map( A1 => n16522, A2 => n17624, B1 => n16778, B2 => 
                           n17621, ZN => n14764);
   U14381 : AOI221_X1 port map( B1 => n17678, B2 => n17275, C1 => n17675, C2 =>
                           n17025, A => n14737, ZN => n14730);
   U14382 : OAI22_X1 port map( A1 => n16547, A2 => n17672, B1 => n16803, B2 => 
                           n17669, ZN => n14737);
   U14383 : AOI221_X1 port map( B1 => n17630, B2 => n17459, C1 => n17627, C2 =>
                           n17026, A => n14745, ZN => n14738);
   U14384 : OAI22_X1 port map( A1 => n16523, A2 => n17624, B1 => n16779, B2 => 
                           n17621, ZN => n14745);
   U14385 : AOI221_X1 port map( B1 => n17678, B2 => n17276, C1 => n17675, C2 =>
                           n17027, A => n14700, ZN => n14679);
   U14386 : OAI22_X1 port map( A1 => n16548, A2 => n17672, B1 => n16804, B2 => 
                           n17669, ZN => n14700);
   U14387 : AOI221_X1 port map( B1 => n17630, B2 => n17460, C1 => n17627, C2 =>
                           n17028, A => n14724, ZN => n14703);
   U14388 : OAI22_X1 port map( A1 => n16524, A2 => n17624, B1 => n16780, B2 => 
                           n17621, ZN => n14724);
   U14389 : AOI221_X1 port map( B1 => n17600, B2 => n17461, C1 => n17597, C2 =>
                           n17029, A => n15502, ZN => n15499);
   U14390 : OAI22_X1 port map( A1 => n16525, A2 => n17594, B1 => n16781, B2 => 
                           n17591, ZN => n15502);
   U14391 : AOI221_X1 port map( B1 => n17600, B2 => n17462, C1 => n17597, C2 =>
                           n17030, A => n15483, ZN => n15480);
   U14392 : OAI22_X1 port map( A1 => n16526, A2 => n17594, B1 => n16782, B2 => 
                           n17591, ZN => n15483);
   U14393 : AOI221_X1 port map( B1 => n17600, B2 => n17463, C1 => n17597, C2 =>
                           n17031, A => n15464, ZN => n15461);
   U14394 : OAI22_X1 port map( A1 => n16527, A2 => n17594, B1 => n16783, B2 => 
                           n17591, ZN => n15464);
   U14395 : AOI221_X1 port map( B1 => n17600, B2 => n17464, C1 => n17597, C2 =>
                           n17032, A => n15445, ZN => n15442);
   U14396 : OAI22_X1 port map( A1 => n16528, A2 => n17594, B1 => n16784, B2 => 
                           n17591, ZN => n15445);
   U14397 : AOI221_X1 port map( B1 => n17600, B2 => n17465, C1 => n17597, C2 =>
                           n17033, A => n15426, ZN => n15423);
   U14398 : OAI22_X1 port map( A1 => n16529, A2 => n17594, B1 => n16785, B2 => 
                           n17591, ZN => n15426);
   U14399 : AOI221_X1 port map( B1 => n17600, B2 => n17466, C1 => n17597, C2 =>
                           n17034, A => n15407, ZN => n15404);
   U14400 : OAI22_X1 port map( A1 => n16530, A2 => n17594, B1 => n16786, B2 => 
                           n17591, ZN => n15407);
   U14401 : AOI221_X1 port map( B1 => n17600, B2 => n17467, C1 => n17597, C2 =>
                           n17035, A => n15388, ZN => n15385);
   U14402 : OAI22_X1 port map( A1 => n16531, A2 => n17594, B1 => n16787, B2 => 
                           n17591, ZN => n15388);
   U14403 : AOI221_X1 port map( B1 => n17600, B2 => n17468, C1 => n17597, C2 =>
                           n17036, A => n15343, ZN => n15334);
   U14404 : OAI22_X1 port map( A1 => n16532, A2 => n17594, B1 => n16788, B2 => 
                           n17591, ZN => n15343);
   U14405 : AOI221_X1 port map( B1 => n17702, B2 => n17461, C1 => n17699, C2 =>
                           n17029, A => n14849, ZN => n14846);
   U14406 : OAI22_X1 port map( A1 => n16525, A2 => n17696, B1 => n16781, B2 => 
                           n17693, ZN => n14849);
   U14407 : AOI221_X1 port map( B1 => n17702, B2 => n17462, C1 => n17699, C2 =>
                           n17030, A => n14830, ZN => n14827);
   U14408 : OAI22_X1 port map( A1 => n16526, A2 => n17696, B1 => n16782, B2 => 
                           n17693, ZN => n14830);
   U14409 : AOI221_X1 port map( B1 => n17702, B2 => n17463, C1 => n17699, C2 =>
                           n17031, A => n14811, ZN => n14808);
   U14410 : OAI22_X1 port map( A1 => n16527, A2 => n17696, B1 => n16783, B2 => 
                           n17693, ZN => n14811);
   U14411 : AOI221_X1 port map( B1 => n17702, B2 => n17464, C1 => n17699, C2 =>
                           n17032, A => n14792, ZN => n14789);
   U14412 : OAI22_X1 port map( A1 => n16528, A2 => n17696, B1 => n16784, B2 => 
                           n17693, ZN => n14792);
   U14413 : AOI221_X1 port map( B1 => n17702, B2 => n17465, C1 => n17699, C2 =>
                           n17033, A => n14773, ZN => n14770);
   U14414 : OAI22_X1 port map( A1 => n16529, A2 => n17696, B1 => n16785, B2 => 
                           n17693, ZN => n14773);
   U14415 : AOI221_X1 port map( B1 => n17702, B2 => n17466, C1 => n17699, C2 =>
                           n17034, A => n14754, ZN => n14751);
   U14416 : OAI22_X1 port map( A1 => n16530, A2 => n17696, B1 => n16786, B2 => 
                           n17693, ZN => n14754);
   U14417 : AOI221_X1 port map( B1 => n17702, B2 => n17467, C1 => n17699, C2 =>
                           n17035, A => n14735, ZN => n14732);
   U14418 : OAI22_X1 port map( A1 => n16531, A2 => n17696, B1 => n16787, B2 => 
                           n17693, ZN => n14735);
   U14419 : AOI221_X1 port map( B1 => n17702, B2 => n17468, C1 => n17699, C2 =>
                           n17036, A => n14690, ZN => n14681);
   U14420 : OAI22_X1 port map( A1 => n16532, A2 => n17696, B1 => n16788, B2 => 
                           n17693, ZN => n14690);
   U14421 : OAI22_X1 port map( A1 => n18102, A2 => n18076, B1 => n14598, B2 => 
                           n16493, ZN => n3609);
   U14422 : OAI22_X1 port map( A1 => n18103, A2 => n18079, B1 => n14598, B2 => 
                           n16494, ZN => n3610);
   U14423 : OAI22_X1 port map( A1 => n18103, A2 => n18082, B1 => n14598, B2 => 
                           n16495, ZN => n3611);
   U14424 : OAI22_X1 port map( A1 => n18103, A2 => n18085, B1 => n14598, B2 => 
                           n16496, ZN => n3612);
   U14425 : OAI22_X1 port map( A1 => n18103, A2 => n18088, B1 => n14598, B2 => 
                           n16497, ZN => n3613);
   U14426 : OAI22_X1 port map( A1 => n18103, A2 => n18091, B1 => n14598, B2 => 
                           n16498, ZN => n3614);
   U14427 : OAI22_X1 port map( A1 => n18104, A2 => n18094, B1 => n14598, B2 => 
                           n16499, ZN => n3615);
   U14428 : OAI22_X1 port map( A1 => n18104, A2 => n18106, B1 => n14598, B2 => 
                           n16500, ZN => n3616);
   U14429 : OAI22_X1 port map( A1 => n17943, A2 => n18076, B1 => n14645, B2 => 
                           n16501, ZN => n3385);
   U14430 : OAI22_X1 port map( A1 => n17944, A2 => n18079, B1 => n14645, B2 => 
                           n16502, ZN => n3386);
   U14431 : OAI22_X1 port map( A1 => n17944, A2 => n18082, B1 => n14645, B2 => 
                           n16503, ZN => n3387);
   U14432 : OAI22_X1 port map( A1 => n17944, A2 => n18085, B1 => n14645, B2 => 
                           n16504, ZN => n3388);
   U14433 : OAI22_X1 port map( A1 => n17944, A2 => n18088, B1 => n14645, B2 => 
                           n16505, ZN => n3389);
   U14434 : OAI22_X1 port map( A1 => n17944, A2 => n18091, B1 => n14645, B2 => 
                           n16506, ZN => n3390);
   U14435 : OAI22_X1 port map( A1 => n17945, A2 => n18094, B1 => n14645, B2 => 
                           n16507, ZN => n3391);
   U14436 : OAI22_X1 port map( A1 => n17945, A2 => n18106, B1 => n14645, B2 => 
                           n16508, ZN => n3392);
   U14437 : OAI22_X1 port map( A1 => n17907, A2 => n18076, B1 => n14652, B2 => 
                           n16509, ZN => n3257);
   U14438 : OAI22_X1 port map( A1 => n17908, A2 => n18079, B1 => n14652, B2 => 
                           n16510, ZN => n3258);
   U14439 : OAI22_X1 port map( A1 => n17908, A2 => n18082, B1 => n14652, B2 => 
                           n16511, ZN => n3259);
   U14440 : OAI22_X1 port map( A1 => n17908, A2 => n18085, B1 => n14652, B2 => 
                           n16512, ZN => n3260);
   U14441 : OAI22_X1 port map( A1 => n17908, A2 => n18088, B1 => n14652, B2 => 
                           n16513, ZN => n3261);
   U14442 : OAI22_X1 port map( A1 => n17908, A2 => n18091, B1 => n14652, B2 => 
                           n16514, ZN => n3262);
   U14443 : OAI22_X1 port map( A1 => n17909, A2 => n18094, B1 => n14652, B2 => 
                           n16515, ZN => n3263);
   U14444 : OAI22_X1 port map( A1 => n17909, A2 => n18106, B1 => n14652, B2 => 
                           n16516, ZN => n3264);
   U14445 : OAI22_X1 port map( A1 => n17871, A2 => n18077, B1 => n14656, B2 => 
                           n16517, ZN => n3129);
   U14446 : OAI22_X1 port map( A1 => n17872, A2 => n18080, B1 => n14656, B2 => 
                           n16518, ZN => n3130);
   U14447 : OAI22_X1 port map( A1 => n17872, A2 => n18083, B1 => n14656, B2 => 
                           n16519, ZN => n3131);
   U14448 : OAI22_X1 port map( A1 => n17872, A2 => n18086, B1 => n14656, B2 => 
                           n16520, ZN => n3132);
   U14449 : OAI22_X1 port map( A1 => n17872, A2 => n18089, B1 => n14656, B2 => 
                           n16521, ZN => n3133);
   U14450 : OAI22_X1 port map( A1 => n17872, A2 => n18092, B1 => n14656, B2 => 
                           n16522, ZN => n3134);
   U14451 : OAI22_X1 port map( A1 => n17873, A2 => n18095, B1 => n14656, B2 => 
                           n16523, ZN => n3135);
   U14452 : OAI22_X1 port map( A1 => n17873, A2 => n18107, B1 => n14656, B2 => 
                           n16524, ZN => n3136);
   U14453 : OAI22_X1 port map( A1 => n17799, A2 => n18077, B1 => n14665, B2 => 
                           n16525, ZN => n2873);
   U14454 : OAI22_X1 port map( A1 => n17800, A2 => n18080, B1 => n14665, B2 => 
                           n16526, ZN => n2874);
   U14455 : OAI22_X1 port map( A1 => n17800, A2 => n18083, B1 => n14665, B2 => 
                           n16527, ZN => n2875);
   U14456 : OAI22_X1 port map( A1 => n17800, A2 => n18086, B1 => n14665, B2 => 
                           n16528, ZN => n2876);
   U14457 : OAI22_X1 port map( A1 => n17800, A2 => n18089, B1 => n14665, B2 => 
                           n16529, ZN => n2877);
   U14458 : OAI22_X1 port map( A1 => n17800, A2 => n18092, B1 => n14665, B2 => 
                           n16530, ZN => n2878);
   U14459 : OAI22_X1 port map( A1 => n17801, A2 => n18095, B1 => n14665, B2 => 
                           n16531, ZN => n2879);
   U14460 : OAI22_X1 port map( A1 => n17801, A2 => n18107, B1 => n14665, B2 => 
                           n16532, ZN => n2880);
   U14461 : OAI22_X1 port map( A1 => n17781, A2 => n18078, B1 => n14668, B2 => 
                           n16533, ZN => n2809);
   U14462 : OAI22_X1 port map( A1 => n17782, A2 => n18081, B1 => n14668, B2 => 
                           n16534, ZN => n2810);
   U14463 : OAI22_X1 port map( A1 => n17782, A2 => n18084, B1 => n14668, B2 => 
                           n16535, ZN => n2811);
   U14464 : OAI22_X1 port map( A1 => n17782, A2 => n18087, B1 => n14668, B2 => 
                           n16536, ZN => n2812);
   U14465 : OAI22_X1 port map( A1 => n17782, A2 => n18090, B1 => n14668, B2 => 
                           n16537, ZN => n2813);
   U14466 : OAI22_X1 port map( A1 => n17782, A2 => n18093, B1 => n14668, B2 => 
                           n16538, ZN => n2814);
   U14467 : OAI22_X1 port map( A1 => n17783, A2 => n18096, B1 => n14668, B2 => 
                           n16539, ZN => n2815);
   U14468 : OAI22_X1 port map( A1 => n17783, A2 => n18108, B1 => n14668, B2 => 
                           n16540, ZN => n2816);
   U14469 : OAI22_X1 port map( A1 => n17745, A2 => n18078, B1 => n14672, B2 => 
                           n16541, ZN => n2681);
   U14470 : OAI22_X1 port map( A1 => n17746, A2 => n18081, B1 => n14672, B2 => 
                           n16542, ZN => n2682);
   U14471 : OAI22_X1 port map( A1 => n17746, A2 => n18084, B1 => n14672, B2 => 
                           n16543, ZN => n2683);
   U14472 : OAI22_X1 port map( A1 => n17746, A2 => n18087, B1 => n14672, B2 => 
                           n16544, ZN => n2684);
   U14473 : OAI22_X1 port map( A1 => n17746, A2 => n18090, B1 => n14672, B2 => 
                           n16545, ZN => n2685);
   U14474 : OAI22_X1 port map( A1 => n17746, A2 => n18093, B1 => n14672, B2 => 
                           n16546, ZN => n2686);
   U14475 : OAI22_X1 port map( A1 => n17747, A2 => n18096, B1 => n14672, B2 => 
                           n16547, ZN => n2687);
   U14476 : OAI22_X1 port map( A1 => n17747, A2 => n18108, B1 => n14672, B2 => 
                           n16548, ZN => n2688);
   U14477 : OAI22_X1 port map( A1 => n17997, A2 => n18076, B1 => n14633, B2 => 
                           n16749, ZN => n3577);
   U14478 : OAI22_X1 port map( A1 => n17998, A2 => n18079, B1 => n14633, B2 => 
                           n16750, ZN => n3578);
   U14479 : OAI22_X1 port map( A1 => n17998, A2 => n18082, B1 => n14633, B2 => 
                           n16751, ZN => n3579);
   U14480 : OAI22_X1 port map( A1 => n17998, A2 => n18085, B1 => n14633, B2 => 
                           n16752, ZN => n3580);
   U14481 : OAI22_X1 port map( A1 => n17998, A2 => n18088, B1 => n14633, B2 => 
                           n16753, ZN => n3581);
   U14482 : OAI22_X1 port map( A1 => n17998, A2 => n18091, B1 => n14633, B2 => 
                           n16754, ZN => n3582);
   U14483 : OAI22_X1 port map( A1 => n17999, A2 => n18094, B1 => n14633, B2 => 
                           n16755, ZN => n3583);
   U14484 : OAI22_X1 port map( A1 => n17999, A2 => n18106, B1 => n14633, B2 => 
                           n16756, ZN => n3584);
   U14485 : OAI22_X1 port map( A1 => n17952, A2 => n18076, B1 => n14643, B2 => 
                           n16757, ZN => n3417);
   U14486 : OAI22_X1 port map( A1 => n17953, A2 => n18079, B1 => n14643, B2 => 
                           n16758, ZN => n3418);
   U14487 : OAI22_X1 port map( A1 => n17953, A2 => n18082, B1 => n14643, B2 => 
                           n16759, ZN => n3419);
   U14488 : OAI22_X1 port map( A1 => n17953, A2 => n18085, B1 => n14643, B2 => 
                           n16760, ZN => n3420);
   U14489 : OAI22_X1 port map( A1 => n17953, A2 => n18088, B1 => n14643, B2 => 
                           n16761, ZN => n3421);
   U14490 : OAI22_X1 port map( A1 => n17953, A2 => n18091, B1 => n14643, B2 => 
                           n16762, ZN => n3422);
   U14491 : OAI22_X1 port map( A1 => n17954, A2 => n18094, B1 => n14643, B2 => 
                           n16763, ZN => n3423);
   U14492 : OAI22_X1 port map( A1 => n17954, A2 => n18106, B1 => n14643, B2 => 
                           n16764, ZN => n3424);
   U14493 : OAI22_X1 port map( A1 => n17916, A2 => n18076, B1 => n14651, B2 => 
                           n16765, ZN => n3289);
   U14494 : OAI22_X1 port map( A1 => n17917, A2 => n18079, B1 => n14651, B2 => 
                           n16766, ZN => n3290);
   U14495 : OAI22_X1 port map( A1 => n17917, A2 => n18082, B1 => n14651, B2 => 
                           n16767, ZN => n3291);
   U14496 : OAI22_X1 port map( A1 => n17917, A2 => n18085, B1 => n14651, B2 => 
                           n16768, ZN => n3292);
   U14497 : OAI22_X1 port map( A1 => n17917, A2 => n18088, B1 => n14651, B2 => 
                           n16769, ZN => n3293);
   U14498 : OAI22_X1 port map( A1 => n17917, A2 => n18091, B1 => n14651, B2 => 
                           n16770, ZN => n3294);
   U14499 : OAI22_X1 port map( A1 => n17918, A2 => n18094, B1 => n14651, B2 => 
                           n16771, ZN => n3295);
   U14500 : OAI22_X1 port map( A1 => n17918, A2 => n18106, B1 => n14651, B2 => 
                           n16772, ZN => n3296);
   U14501 : OAI22_X1 port map( A1 => n17880, A2 => n18077, B1 => n14655, B2 => 
                           n16773, ZN => n3161);
   U14502 : OAI22_X1 port map( A1 => n17881, A2 => n18080, B1 => n14655, B2 => 
                           n16774, ZN => n3162);
   U14503 : OAI22_X1 port map( A1 => n17881, A2 => n18083, B1 => n14655, B2 => 
                           n16775, ZN => n3163);
   U14504 : OAI22_X1 port map( A1 => n17881, A2 => n18086, B1 => n14655, B2 => 
                           n16776, ZN => n3164);
   U14505 : OAI22_X1 port map( A1 => n17881, A2 => n18089, B1 => n14655, B2 => 
                           n16777, ZN => n3165);
   U14506 : OAI22_X1 port map( A1 => n17881, A2 => n18092, B1 => n14655, B2 => 
                           n16778, ZN => n3166);
   U14507 : OAI22_X1 port map( A1 => n17882, A2 => n18095, B1 => n14655, B2 => 
                           n16779, ZN => n3167);
   U14508 : OAI22_X1 port map( A1 => n17882, A2 => n18107, B1 => n14655, B2 => 
                           n16780, ZN => n3168);
   U14509 : OAI22_X1 port map( A1 => n17808, A2 => n18077, B1 => n14664, B2 => 
                           n16781, ZN => n2905);
   U14510 : OAI22_X1 port map( A1 => n17809, A2 => n18080, B1 => n14664, B2 => 
                           n16782, ZN => n2906);
   U14511 : OAI22_X1 port map( A1 => n17809, A2 => n18083, B1 => n14664, B2 => 
                           n16783, ZN => n2907);
   U14512 : OAI22_X1 port map( A1 => n17809, A2 => n18086, B1 => n14664, B2 => 
                           n16784, ZN => n2908);
   U14513 : OAI22_X1 port map( A1 => n17809, A2 => n18089, B1 => n14664, B2 => 
                           n16785, ZN => n2909);
   U14514 : OAI22_X1 port map( A1 => n17809, A2 => n18092, B1 => n14664, B2 => 
                           n16786, ZN => n2910);
   U14515 : OAI22_X1 port map( A1 => n17810, A2 => n18095, B1 => n14664, B2 => 
                           n16787, ZN => n2911);
   U14516 : OAI22_X1 port map( A1 => n17810, A2 => n18107, B1 => n14664, B2 => 
                           n16788, ZN => n2912);
   U14517 : OAI22_X1 port map( A1 => n17790, A2 => n18078, B1 => n14666, B2 => 
                           n16789, ZN => n2841);
   U14518 : OAI22_X1 port map( A1 => n17791, A2 => n18081, B1 => n14666, B2 => 
                           n16790, ZN => n2842);
   U14519 : OAI22_X1 port map( A1 => n17791, A2 => n18084, B1 => n14666, B2 => 
                           n16791, ZN => n2843);
   U14520 : OAI22_X1 port map( A1 => n17791, A2 => n18087, B1 => n14666, B2 => 
                           n16792, ZN => n2844);
   U14521 : OAI22_X1 port map( A1 => n17791, A2 => n18090, B1 => n14666, B2 => 
                           n16793, ZN => n2845);
   U14522 : OAI22_X1 port map( A1 => n17791, A2 => n18093, B1 => n14666, B2 => 
                           n16794, ZN => n2846);
   U14523 : OAI22_X1 port map( A1 => n17792, A2 => n18096, B1 => n14666, B2 => 
                           n16795, ZN => n2847);
   U14524 : OAI22_X1 port map( A1 => n17792, A2 => n18108, B1 => n14666, B2 => 
                           n16796, ZN => n2848);
   U14525 : OAI22_X1 port map( A1 => n17754, A2 => n18078, B1 => n14671, B2 => 
                           n16797, ZN => n2713);
   U14526 : OAI22_X1 port map( A1 => n17755, A2 => n18081, B1 => n14671, B2 => 
                           n16798, ZN => n2714);
   U14527 : OAI22_X1 port map( A1 => n17755, A2 => n18084, B1 => n14671, B2 => 
                           n16799, ZN => n2715);
   U14528 : OAI22_X1 port map( A1 => n17755, A2 => n18087, B1 => n14671, B2 => 
                           n16800, ZN => n2716);
   U14529 : OAI22_X1 port map( A1 => n17755, A2 => n18090, B1 => n14671, B2 => 
                           n16801, ZN => n2717);
   U14530 : OAI22_X1 port map( A1 => n17755, A2 => n18093, B1 => n14671, B2 => 
                           n16802, ZN => n2718);
   U14531 : OAI22_X1 port map( A1 => n17756, A2 => n18096, B1 => n14671, B2 => 
                           n16803, ZN => n2719);
   U14532 : OAI22_X1 port map( A1 => n17756, A2 => n18108, B1 => n14671, B2 => 
                           n16804, ZN => n2720);
   U14533 : OAI22_X1 port map( A1 => n17864, A2 => n18107, B1 => n14657, B2 => 
                           n16812, ZN => n3104);
   U14534 : OAI22_X1 port map( A1 => n17862, A2 => n18077, B1 => n14657, B2 => 
                           n16805, ZN => n3097);
   U14535 : OAI22_X1 port map( A1 => n17863, A2 => n18080, B1 => n14657, B2 => 
                           n16806, ZN => n3098);
   U14536 : OAI22_X1 port map( A1 => n17863, A2 => n18083, B1 => n14657, B2 => 
                           n16807, ZN => n3099);
   U14537 : OAI22_X1 port map( A1 => n17863, A2 => n18086, B1 => n14657, B2 => 
                           n16808, ZN => n3100);
   U14538 : OAI22_X1 port map( A1 => n17863, A2 => n18089, B1 => n14657, B2 => 
                           n16809, ZN => n3101);
   U14539 : OAI22_X1 port map( A1 => n17863, A2 => n18092, B1 => n14657, B2 => 
                           n16810, ZN => n3102);
   U14540 : OAI22_X1 port map( A1 => n17864, A2 => n18095, B1 => n14657, B2 => 
                           n16811, ZN => n3103);
   U14541 : OAI22_X1 port map( A1 => n17853, A2 => n18077, B1 => n14659, B2 => 
                           n16645, ZN => n3065);
   U14542 : OAI22_X1 port map( A1 => n17854, A2 => n18080, B1 => n14659, B2 => 
                           n16646, ZN => n3066);
   U14543 : OAI22_X1 port map( A1 => n17854, A2 => n18083, B1 => n14659, B2 => 
                           n16647, ZN => n3067);
   U14544 : OAI22_X1 port map( A1 => n17854, A2 => n18086, B1 => n14659, B2 => 
                           n16648, ZN => n3068);
   U14545 : OAI22_X1 port map( A1 => n17854, A2 => n18089, B1 => n14659, B2 => 
                           n16649, ZN => n3069);
   U14546 : OAI22_X1 port map( A1 => n17854, A2 => n18092, B1 => n14659, B2 => 
                           n16650, ZN => n3070);
   U14547 : OAI22_X1 port map( A1 => n17855, A2 => n18095, B1 => n14659, B2 => 
                           n16651, ZN => n3071);
   U14548 : OAI22_X1 port map( A1 => n17855, A2 => n18107, B1 => n14659, B2 => 
                           n16652, ZN => n3072);
   U14549 : OAI22_X1 port map( A1 => n18098, A2 => n18004, B1 => n18097, B2 => 
                           n16653, ZN => n3585);
   U14550 : OAI22_X1 port map( A1 => n18098, A2 => n18007, B1 => n18097, B2 => 
                           n16654, ZN => n3586);
   U14551 : OAI22_X1 port map( A1 => n18098, A2 => n18010, B1 => n18097, B2 => 
                           n16655, ZN => n3587);
   U14552 : OAI22_X1 port map( A1 => n18098, A2 => n18013, B1 => n18097, B2 => 
                           n16656, ZN => n3588);
   U14553 : OAI22_X1 port map( A1 => n18098, A2 => n18016, B1 => n18097, B2 => 
                           n16657, ZN => n3589);
   U14554 : OAI22_X1 port map( A1 => n18099, A2 => n18019, B1 => n18097, B2 => 
                           n16658, ZN => n3590);
   U14555 : OAI22_X1 port map( A1 => n18099, A2 => n18022, B1 => n18097, B2 => 
                           n16659, ZN => n3591);
   U14556 : OAI22_X1 port map( A1 => n18099, A2 => n18025, B1 => n18097, B2 => 
                           n16660, ZN => n3592);
   U14557 : OAI22_X1 port map( A1 => n18099, A2 => n18028, B1 => n18097, B2 => 
                           n16661, ZN => n3593);
   U14558 : OAI22_X1 port map( A1 => n18099, A2 => n18031, B1 => n18097, B2 => 
                           n16662, ZN => n3594);
   U14559 : OAI22_X1 port map( A1 => n18100, A2 => n18034, B1 => n18097, B2 => 
                           n16663, ZN => n3595);
   U14560 : OAI22_X1 port map( A1 => n18100, A2 => n18037, B1 => n18097, B2 => 
                           n16664, ZN => n3596);
   U14561 : OAI22_X1 port map( A1 => n18100, A2 => n18040, B1 => n14598, B2 => 
                           n16549, ZN => n3597);
   U14562 : OAI22_X1 port map( A1 => n18100, A2 => n18043, B1 => n14598, B2 => 
                           n16550, ZN => n3598);
   U14563 : OAI22_X1 port map( A1 => n18100, A2 => n18046, B1 => n14598, B2 => 
                           n16551, ZN => n3599);
   U14564 : OAI22_X1 port map( A1 => n18101, A2 => n18049, B1 => n18097, B2 => 
                           n16552, ZN => n3600);
   U14565 : OAI22_X1 port map( A1 => n18101, A2 => n18052, B1 => n18097, B2 => 
                           n16553, ZN => n3601);
   U14566 : OAI22_X1 port map( A1 => n18101, A2 => n18055, B1 => n18097, B2 => 
                           n16554, ZN => n3602);
   U14567 : OAI22_X1 port map( A1 => n18101, A2 => n18058, B1 => n18097, B2 => 
                           n16555, ZN => n3603);
   U14568 : OAI22_X1 port map( A1 => n18101, A2 => n18061, B1 => n18097, B2 => 
                           n16556, ZN => n3604);
   U14569 : OAI22_X1 port map( A1 => n18102, A2 => n18064, B1 => n18097, B2 => 
                           n16557, ZN => n3605);
   U14570 : OAI22_X1 port map( A1 => n18102, A2 => n18067, B1 => n18097, B2 => 
                           n16558, ZN => n3606);
   U14571 : OAI22_X1 port map( A1 => n18102, A2 => n18070, B1 => n18097, B2 => 
                           n16559, ZN => n3607);
   U14572 : OAI22_X1 port map( A1 => n18102, A2 => n18073, B1 => n18097, B2 => 
                           n16560, ZN => n3608);
   U14573 : OAI22_X1 port map( A1 => n17939, A2 => n18004, B1 => n17938, B2 => 
                           n16665, ZN => n3361);
   U14574 : OAI22_X1 port map( A1 => n17939, A2 => n18007, B1 => n17938, B2 => 
                           n16666, ZN => n3362);
   U14575 : OAI22_X1 port map( A1 => n17939, A2 => n18010, B1 => n17938, B2 => 
                           n16667, ZN => n3363);
   U14576 : OAI22_X1 port map( A1 => n17939, A2 => n18013, B1 => n17938, B2 => 
                           n16668, ZN => n3364);
   U14577 : OAI22_X1 port map( A1 => n17939, A2 => n18016, B1 => n17938, B2 => 
                           n16669, ZN => n3365);
   U14578 : OAI22_X1 port map( A1 => n17940, A2 => n18019, B1 => n17938, B2 => 
                           n16670, ZN => n3366);
   U14579 : OAI22_X1 port map( A1 => n17940, A2 => n18022, B1 => n17938, B2 => 
                           n16671, ZN => n3367);
   U14580 : OAI22_X1 port map( A1 => n17940, A2 => n18025, B1 => n17938, B2 => 
                           n16672, ZN => n3368);
   U14581 : OAI22_X1 port map( A1 => n17940, A2 => n18028, B1 => n17938, B2 => 
                           n16673, ZN => n3369);
   U14582 : OAI22_X1 port map( A1 => n17940, A2 => n18031, B1 => n17938, B2 => 
                           n16674, ZN => n3370);
   U14583 : OAI22_X1 port map( A1 => n17941, A2 => n18034, B1 => n17938, B2 => 
                           n16675, ZN => n3371);
   U14584 : OAI22_X1 port map( A1 => n17941, A2 => n18037, B1 => n17938, B2 => 
                           n16676, ZN => n3372);
   U14585 : OAI22_X1 port map( A1 => n17941, A2 => n18040, B1 => n14645, B2 => 
                           n16561, ZN => n3373);
   U14586 : OAI22_X1 port map( A1 => n17941, A2 => n18043, B1 => n14645, B2 => 
                           n16562, ZN => n3374);
   U14587 : OAI22_X1 port map( A1 => n17941, A2 => n18046, B1 => n14645, B2 => 
                           n16563, ZN => n3375);
   U14588 : OAI22_X1 port map( A1 => n17942, A2 => n18049, B1 => n17938, B2 => 
                           n16564, ZN => n3376);
   U14589 : OAI22_X1 port map( A1 => n17942, A2 => n18052, B1 => n17938, B2 => 
                           n16565, ZN => n3377);
   U14590 : OAI22_X1 port map( A1 => n17942, A2 => n18055, B1 => n17938, B2 => 
                           n16566, ZN => n3378);
   U14591 : OAI22_X1 port map( A1 => n17942, A2 => n18058, B1 => n17938, B2 => 
                           n16567, ZN => n3379);
   U14592 : OAI22_X1 port map( A1 => n17942, A2 => n18061, B1 => n17938, B2 => 
                           n16568, ZN => n3380);
   U14593 : OAI22_X1 port map( A1 => n17943, A2 => n18064, B1 => n17938, B2 => 
                           n16569, ZN => n3381);
   U14594 : OAI22_X1 port map( A1 => n17943, A2 => n18067, B1 => n17938, B2 => 
                           n16570, ZN => n3382);
   U14595 : OAI22_X1 port map( A1 => n17943, A2 => n18070, B1 => n17938, B2 => 
                           n16571, ZN => n3383);
   U14596 : OAI22_X1 port map( A1 => n17943, A2 => n18073, B1 => n17938, B2 => 
                           n16572, ZN => n3384);
   U14597 : OAI22_X1 port map( A1 => n17903, A2 => n18004, B1 => n17902, B2 => 
                           n16677, ZN => n3233);
   U14598 : OAI22_X1 port map( A1 => n17903, A2 => n18007, B1 => n17902, B2 => 
                           n16678, ZN => n3234);
   U14599 : OAI22_X1 port map( A1 => n17903, A2 => n18010, B1 => n17902, B2 => 
                           n16679, ZN => n3235);
   U14600 : OAI22_X1 port map( A1 => n17903, A2 => n18013, B1 => n17902, B2 => 
                           n16680, ZN => n3236);
   U14601 : OAI22_X1 port map( A1 => n17903, A2 => n18016, B1 => n17902, B2 => 
                           n16681, ZN => n3237);
   U14602 : OAI22_X1 port map( A1 => n17904, A2 => n18019, B1 => n17902, B2 => 
                           n16682, ZN => n3238);
   U14603 : OAI22_X1 port map( A1 => n17904, A2 => n18022, B1 => n17902, B2 => 
                           n16683, ZN => n3239);
   U14604 : OAI22_X1 port map( A1 => n17904, A2 => n18025, B1 => n17902, B2 => 
                           n16684, ZN => n3240);
   U14605 : OAI22_X1 port map( A1 => n17904, A2 => n18028, B1 => n17902, B2 => 
                           n16685, ZN => n3241);
   U14606 : OAI22_X1 port map( A1 => n17904, A2 => n18031, B1 => n17902, B2 => 
                           n16686, ZN => n3242);
   U14607 : OAI22_X1 port map( A1 => n17905, A2 => n18034, B1 => n17902, B2 => 
                           n16687, ZN => n3243);
   U14608 : OAI22_X1 port map( A1 => n17905, A2 => n18037, B1 => n17902, B2 => 
                           n16688, ZN => n3244);
   U14609 : OAI22_X1 port map( A1 => n17905, A2 => n18040, B1 => n14652, B2 => 
                           n16573, ZN => n3245);
   U14610 : OAI22_X1 port map( A1 => n17905, A2 => n18043, B1 => n14652, B2 => 
                           n16574, ZN => n3246);
   U14611 : OAI22_X1 port map( A1 => n17905, A2 => n18046, B1 => n14652, B2 => 
                           n16575, ZN => n3247);
   U14612 : OAI22_X1 port map( A1 => n17906, A2 => n18049, B1 => n17902, B2 => 
                           n16576, ZN => n3248);
   U14613 : OAI22_X1 port map( A1 => n17906, A2 => n18052, B1 => n17902, B2 => 
                           n16577, ZN => n3249);
   U14614 : OAI22_X1 port map( A1 => n17906, A2 => n18055, B1 => n17902, B2 => 
                           n16578, ZN => n3250);
   U14615 : OAI22_X1 port map( A1 => n17906, A2 => n18058, B1 => n17902, B2 => 
                           n16579, ZN => n3251);
   U14616 : OAI22_X1 port map( A1 => n17906, A2 => n18061, B1 => n17902, B2 => 
                           n16580, ZN => n3252);
   U14617 : OAI22_X1 port map( A1 => n17907, A2 => n18064, B1 => n17902, B2 => 
                           n16581, ZN => n3253);
   U14618 : OAI22_X1 port map( A1 => n17907, A2 => n18067, B1 => n17902, B2 => 
                           n16582, ZN => n3254);
   U14619 : OAI22_X1 port map( A1 => n17907, A2 => n18070, B1 => n17902, B2 => 
                           n16583, ZN => n3255);
   U14620 : OAI22_X1 port map( A1 => n17907, A2 => n18073, B1 => n17902, B2 => 
                           n16584, ZN => n3256);
   U14621 : OAI22_X1 port map( A1 => n17867, A2 => n18005, B1 => n17866, B2 => 
                           n16689, ZN => n3105);
   U14622 : OAI22_X1 port map( A1 => n17867, A2 => n18008, B1 => n17866, B2 => 
                           n16690, ZN => n3106);
   U14623 : OAI22_X1 port map( A1 => n17867, A2 => n18011, B1 => n17866, B2 => 
                           n16691, ZN => n3107);
   U14624 : OAI22_X1 port map( A1 => n17867, A2 => n18014, B1 => n17866, B2 => 
                           n16692, ZN => n3108);
   U14625 : OAI22_X1 port map( A1 => n17867, A2 => n18017, B1 => n17866, B2 => 
                           n16693, ZN => n3109);
   U14626 : OAI22_X1 port map( A1 => n17868, A2 => n18020, B1 => n17866, B2 => 
                           n16694, ZN => n3110);
   U14627 : OAI22_X1 port map( A1 => n17868, A2 => n18023, B1 => n17866, B2 => 
                           n16695, ZN => n3111);
   U14628 : OAI22_X1 port map( A1 => n17868, A2 => n18026, B1 => n17866, B2 => 
                           n16696, ZN => n3112);
   U14629 : OAI22_X1 port map( A1 => n17868, A2 => n18029, B1 => n17866, B2 => 
                           n16697, ZN => n3113);
   U14630 : OAI22_X1 port map( A1 => n17868, A2 => n18032, B1 => n17866, B2 => 
                           n16698, ZN => n3114);
   U14631 : OAI22_X1 port map( A1 => n17869, A2 => n18035, B1 => n17866, B2 => 
                           n16699, ZN => n3115);
   U14632 : OAI22_X1 port map( A1 => n17869, A2 => n18038, B1 => n17866, B2 => 
                           n16700, ZN => n3116);
   U14633 : OAI22_X1 port map( A1 => n17869, A2 => n18041, B1 => n14656, B2 => 
                           n16585, ZN => n3117);
   U14634 : OAI22_X1 port map( A1 => n17869, A2 => n18044, B1 => n14656, B2 => 
                           n16586, ZN => n3118);
   U14635 : OAI22_X1 port map( A1 => n17869, A2 => n18047, B1 => n14656, B2 => 
                           n16587, ZN => n3119);
   U14636 : OAI22_X1 port map( A1 => n17870, A2 => n18050, B1 => n17866, B2 => 
                           n16588, ZN => n3120);
   U14637 : OAI22_X1 port map( A1 => n17870, A2 => n18053, B1 => n17866, B2 => 
                           n16589, ZN => n3121);
   U14638 : OAI22_X1 port map( A1 => n17870, A2 => n18056, B1 => n17866, B2 => 
                           n16590, ZN => n3122);
   U14639 : OAI22_X1 port map( A1 => n17870, A2 => n18059, B1 => n17866, B2 => 
                           n16591, ZN => n3123);
   U14640 : OAI22_X1 port map( A1 => n17870, A2 => n18062, B1 => n17866, B2 => 
                           n16592, ZN => n3124);
   U14641 : OAI22_X1 port map( A1 => n17871, A2 => n18065, B1 => n17866, B2 => 
                           n16593, ZN => n3125);
   U14642 : OAI22_X1 port map( A1 => n17871, A2 => n18068, B1 => n17866, B2 => 
                           n16594, ZN => n3126);
   U14643 : OAI22_X1 port map( A1 => n17871, A2 => n18071, B1 => n17866, B2 => 
                           n16595, ZN => n3127);
   U14644 : OAI22_X1 port map( A1 => n17871, A2 => n18074, B1 => n17866, B2 => 
                           n16596, ZN => n3128);
   U14645 : OAI22_X1 port map( A1 => n17795, A2 => n18005, B1 => n17794, B2 => 
                           n16701, ZN => n2849);
   U14646 : OAI22_X1 port map( A1 => n17795, A2 => n18008, B1 => n17794, B2 => 
                           n16702, ZN => n2850);
   U14647 : OAI22_X1 port map( A1 => n17795, A2 => n18011, B1 => n17794, B2 => 
                           n16703, ZN => n2851);
   U14648 : OAI22_X1 port map( A1 => n17795, A2 => n18014, B1 => n17794, B2 => 
                           n16704, ZN => n2852);
   U14649 : OAI22_X1 port map( A1 => n17795, A2 => n18017, B1 => n17794, B2 => 
                           n16705, ZN => n2853);
   U14650 : OAI22_X1 port map( A1 => n17796, A2 => n18020, B1 => n17794, B2 => 
                           n16706, ZN => n2854);
   U14651 : OAI22_X1 port map( A1 => n17796, A2 => n18023, B1 => n17794, B2 => 
                           n16707, ZN => n2855);
   U14652 : OAI22_X1 port map( A1 => n17796, A2 => n18026, B1 => n17794, B2 => 
                           n16708, ZN => n2856);
   U14653 : OAI22_X1 port map( A1 => n17796, A2 => n18029, B1 => n17794, B2 => 
                           n16709, ZN => n2857);
   U14654 : OAI22_X1 port map( A1 => n17796, A2 => n18032, B1 => n17794, B2 => 
                           n16710, ZN => n2858);
   U14655 : OAI22_X1 port map( A1 => n17797, A2 => n18035, B1 => n17794, B2 => 
                           n16711, ZN => n2859);
   U14656 : OAI22_X1 port map( A1 => n17797, A2 => n18038, B1 => n17794, B2 => 
                           n16712, ZN => n2860);
   U14657 : OAI22_X1 port map( A1 => n17797, A2 => n18041, B1 => n14665, B2 => 
                           n16597, ZN => n2861);
   U14658 : OAI22_X1 port map( A1 => n17797, A2 => n18044, B1 => n14665, B2 => 
                           n16598, ZN => n2862);
   U14659 : OAI22_X1 port map( A1 => n17797, A2 => n18047, B1 => n14665, B2 => 
                           n16599, ZN => n2863);
   U14660 : OAI22_X1 port map( A1 => n17798, A2 => n18050, B1 => n17794, B2 => 
                           n16600, ZN => n2864);
   U14661 : OAI22_X1 port map( A1 => n17798, A2 => n18053, B1 => n17794, B2 => 
                           n16601, ZN => n2865);
   U14662 : OAI22_X1 port map( A1 => n17798, A2 => n18056, B1 => n17794, B2 => 
                           n16602, ZN => n2866);
   U14663 : OAI22_X1 port map( A1 => n17798, A2 => n18059, B1 => n17794, B2 => 
                           n16603, ZN => n2867);
   U14664 : OAI22_X1 port map( A1 => n17798, A2 => n18062, B1 => n17794, B2 => 
                           n16604, ZN => n2868);
   U14665 : OAI22_X1 port map( A1 => n17799, A2 => n18065, B1 => n17794, B2 => 
                           n16605, ZN => n2869);
   U14666 : OAI22_X1 port map( A1 => n17799, A2 => n18068, B1 => n17794, B2 => 
                           n16606, ZN => n2870);
   U14667 : OAI22_X1 port map( A1 => n17799, A2 => n18071, B1 => n17794, B2 => 
                           n16607, ZN => n2871);
   U14668 : OAI22_X1 port map( A1 => n17799, A2 => n18074, B1 => n17794, B2 => 
                           n16608, ZN => n2872);
   U14669 : OAI22_X1 port map( A1 => n17777, A2 => n18006, B1 => n17776, B2 => 
                           n16713, ZN => n2785);
   U14670 : OAI22_X1 port map( A1 => n17777, A2 => n18009, B1 => n17776, B2 => 
                           n16714, ZN => n2786);
   U14671 : OAI22_X1 port map( A1 => n17777, A2 => n18012, B1 => n17776, B2 => 
                           n16715, ZN => n2787);
   U14672 : OAI22_X1 port map( A1 => n17777, A2 => n18015, B1 => n17776, B2 => 
                           n16716, ZN => n2788);
   U14673 : OAI22_X1 port map( A1 => n17777, A2 => n18018, B1 => n17776, B2 => 
                           n16717, ZN => n2789);
   U14674 : OAI22_X1 port map( A1 => n17778, A2 => n18021, B1 => n17776, B2 => 
                           n16718, ZN => n2790);
   U14675 : OAI22_X1 port map( A1 => n17778, A2 => n18024, B1 => n17776, B2 => 
                           n16719, ZN => n2791);
   U14676 : OAI22_X1 port map( A1 => n17778, A2 => n18027, B1 => n17776, B2 => 
                           n16720, ZN => n2792);
   U14677 : OAI22_X1 port map( A1 => n17778, A2 => n18030, B1 => n17776, B2 => 
                           n16721, ZN => n2793);
   U14678 : OAI22_X1 port map( A1 => n17778, A2 => n18033, B1 => n17776, B2 => 
                           n16722, ZN => n2794);
   U14679 : OAI22_X1 port map( A1 => n17779, A2 => n18036, B1 => n17776, B2 => 
                           n16723, ZN => n2795);
   U14680 : OAI22_X1 port map( A1 => n17779, A2 => n18039, B1 => n17776, B2 => 
                           n16724, ZN => n2796);
   U14681 : OAI22_X1 port map( A1 => n17779, A2 => n18042, B1 => n14668, B2 => 
                           n16609, ZN => n2797);
   U14682 : OAI22_X1 port map( A1 => n17779, A2 => n18045, B1 => n14668, B2 => 
                           n16610, ZN => n2798);
   U14683 : OAI22_X1 port map( A1 => n17779, A2 => n18048, B1 => n14668, B2 => 
                           n16611, ZN => n2799);
   U14684 : OAI22_X1 port map( A1 => n17780, A2 => n18051, B1 => n17776, B2 => 
                           n16612, ZN => n2800);
   U14685 : OAI22_X1 port map( A1 => n17780, A2 => n18054, B1 => n17776, B2 => 
                           n16613, ZN => n2801);
   U14686 : OAI22_X1 port map( A1 => n17780, A2 => n18057, B1 => n17776, B2 => 
                           n16614, ZN => n2802);
   U14687 : OAI22_X1 port map( A1 => n17780, A2 => n18060, B1 => n17776, B2 => 
                           n16615, ZN => n2803);
   U14688 : OAI22_X1 port map( A1 => n17780, A2 => n18063, B1 => n17776, B2 => 
                           n16616, ZN => n2804);
   U14689 : OAI22_X1 port map( A1 => n17781, A2 => n18066, B1 => n17776, B2 => 
                           n16617, ZN => n2805);
   U14690 : OAI22_X1 port map( A1 => n17781, A2 => n18069, B1 => n17776, B2 => 
                           n16618, ZN => n2806);
   U14691 : OAI22_X1 port map( A1 => n17781, A2 => n18072, B1 => n17776, B2 => 
                           n16619, ZN => n2807);
   U14692 : OAI22_X1 port map( A1 => n17781, A2 => n18075, B1 => n17776, B2 => 
                           n16620, ZN => n2808);
   U14693 : OAI22_X1 port map( A1 => n17741, A2 => n18006, B1 => n17740, B2 => 
                           n16725, ZN => n2657);
   U14694 : OAI22_X1 port map( A1 => n17741, A2 => n18009, B1 => n17740, B2 => 
                           n16726, ZN => n2658);
   U14695 : OAI22_X1 port map( A1 => n17741, A2 => n18012, B1 => n17740, B2 => 
                           n16727, ZN => n2659);
   U14696 : OAI22_X1 port map( A1 => n17741, A2 => n18015, B1 => n17740, B2 => 
                           n16728, ZN => n2660);
   U14697 : OAI22_X1 port map( A1 => n17741, A2 => n18018, B1 => n17740, B2 => 
                           n16729, ZN => n2661);
   U14698 : OAI22_X1 port map( A1 => n17742, A2 => n18021, B1 => n17740, B2 => 
                           n16730, ZN => n2662);
   U14699 : OAI22_X1 port map( A1 => n17742, A2 => n18024, B1 => n17740, B2 => 
                           n16731, ZN => n2663);
   U14700 : OAI22_X1 port map( A1 => n17742, A2 => n18027, B1 => n17740, B2 => 
                           n16732, ZN => n2664);
   U14701 : OAI22_X1 port map( A1 => n17742, A2 => n18030, B1 => n17740, B2 => 
                           n16733, ZN => n2665);
   U14702 : OAI22_X1 port map( A1 => n17742, A2 => n18033, B1 => n17740, B2 => 
                           n16734, ZN => n2666);
   U14703 : OAI22_X1 port map( A1 => n17743, A2 => n18036, B1 => n17740, B2 => 
                           n16735, ZN => n2667);
   U14704 : OAI22_X1 port map( A1 => n17743, A2 => n18039, B1 => n17740, B2 => 
                           n16736, ZN => n2668);
   U14705 : OAI22_X1 port map( A1 => n17743, A2 => n18042, B1 => n14672, B2 => 
                           n16621, ZN => n2669);
   U14706 : OAI22_X1 port map( A1 => n17743, A2 => n18045, B1 => n14672, B2 => 
                           n16622, ZN => n2670);
   U14707 : OAI22_X1 port map( A1 => n17743, A2 => n18048, B1 => n14672, B2 => 
                           n16623, ZN => n2671);
   U14708 : OAI22_X1 port map( A1 => n17744, A2 => n18051, B1 => n17740, B2 => 
                           n16624, ZN => n2672);
   U14709 : OAI22_X1 port map( A1 => n17744, A2 => n18054, B1 => n17740, B2 => 
                           n16625, ZN => n2673);
   U14710 : OAI22_X1 port map( A1 => n17744, A2 => n18057, B1 => n17740, B2 => 
                           n16626, ZN => n2674);
   U14711 : OAI22_X1 port map( A1 => n17744, A2 => n18060, B1 => n17740, B2 => 
                           n16627, ZN => n2675);
   U14712 : OAI22_X1 port map( A1 => n17744, A2 => n18063, B1 => n17740, B2 => 
                           n16628, ZN => n2676);
   U14713 : OAI22_X1 port map( A1 => n17745, A2 => n18066, B1 => n17740, B2 => 
                           n16629, ZN => n2677);
   U14714 : OAI22_X1 port map( A1 => n17745, A2 => n18069, B1 => n17740, B2 => 
                           n16630, ZN => n2678);
   U14715 : OAI22_X1 port map( A1 => n17745, A2 => n18072, B1 => n17740, B2 => 
                           n16631, ZN => n2679);
   U14716 : OAI22_X1 port map( A1 => n17745, A2 => n18075, B1 => n17740, B2 => 
                           n16632, ZN => n2680);
   U14717 : OAI22_X1 port map( A1 => n17993, A2 => n18004, B1 => n17992, B2 => 
                           n17053, ZN => n3553);
   U14718 : OAI22_X1 port map( A1 => n17993, A2 => n18007, B1 => n17992, B2 => 
                           n17054, ZN => n3554);
   U14719 : OAI22_X1 port map( A1 => n17993, A2 => n18010, B1 => n17992, B2 => 
                           n17055, ZN => n3555);
   U14720 : OAI22_X1 port map( A1 => n17993, A2 => n18013, B1 => n17992, B2 => 
                           n17056, ZN => n3556);
   U14721 : OAI22_X1 port map( A1 => n17993, A2 => n18016, B1 => n17992, B2 => 
                           n17057, ZN => n3557);
   U14722 : OAI22_X1 port map( A1 => n17994, A2 => n18019, B1 => n17992, B2 => 
                           n17058, ZN => n3558);
   U14723 : OAI22_X1 port map( A1 => n17994, A2 => n18022, B1 => n17992, B2 => 
                           n17059, ZN => n3559);
   U14724 : OAI22_X1 port map( A1 => n17994, A2 => n18025, B1 => n17992, B2 => 
                           n17060, ZN => n3560);
   U14725 : OAI22_X1 port map( A1 => n17994, A2 => n18028, B1 => n17992, B2 => 
                           n17061, ZN => n3561);
   U14726 : OAI22_X1 port map( A1 => n17994, A2 => n18031, B1 => n17992, B2 => 
                           n17062, ZN => n3562);
   U14727 : OAI22_X1 port map( A1 => n17995, A2 => n18034, B1 => n17992, B2 => 
                           n17063, ZN => n3563);
   U14728 : OAI22_X1 port map( A1 => n17995, A2 => n18037, B1 => n17992, B2 => 
                           n17064, ZN => n3564);
   U14729 : OAI22_X1 port map( A1 => n17995, A2 => n18040, B1 => n14633, B2 => 
                           n17065, ZN => n3565);
   U14730 : OAI22_X1 port map( A1 => n17995, A2 => n18043, B1 => n14633, B2 => 
                           n17066, ZN => n3566);
   U14731 : OAI22_X1 port map( A1 => n17995, A2 => n18046, B1 => n14633, B2 => 
                           n17067, ZN => n3567);
   U14732 : OAI22_X1 port map( A1 => n17996, A2 => n18049, B1 => n17992, B2 => 
                           n17068, ZN => n3568);
   U14733 : OAI22_X1 port map( A1 => n17996, A2 => n18052, B1 => n17992, B2 => 
                           n17069, ZN => n3569);
   U14734 : OAI22_X1 port map( A1 => n17996, A2 => n18055, B1 => n17992, B2 => 
                           n17070, ZN => n3570);
   U14735 : OAI22_X1 port map( A1 => n17996, A2 => n18058, B1 => n17992, B2 => 
                           n17071, ZN => n3571);
   U14736 : OAI22_X1 port map( A1 => n17996, A2 => n18061, B1 => n17992, B2 => 
                           n17072, ZN => n3572);
   U14737 : OAI22_X1 port map( A1 => n17997, A2 => n18064, B1 => n17992, B2 => 
                           n17073, ZN => n3573);
   U14738 : OAI22_X1 port map( A1 => n17997, A2 => n18067, B1 => n17992, B2 => 
                           n17074, ZN => n3574);
   U14739 : OAI22_X1 port map( A1 => n17997, A2 => n18070, B1 => n17992, B2 => 
                           n17075, ZN => n3575);
   U14740 : OAI22_X1 port map( A1 => n17997, A2 => n18073, B1 => n17992, B2 => 
                           n17076, ZN => n3576);
   U14741 : OAI22_X1 port map( A1 => n17948, A2 => n18004, B1 => n17947, B2 => 
                           n17077, ZN => n3393);
   U14742 : OAI22_X1 port map( A1 => n17948, A2 => n18007, B1 => n17947, B2 => 
                           n17078, ZN => n3394);
   U14743 : OAI22_X1 port map( A1 => n17948, A2 => n18010, B1 => n17947, B2 => 
                           n17079, ZN => n3395);
   U14744 : OAI22_X1 port map( A1 => n17948, A2 => n18013, B1 => n17947, B2 => 
                           n17080, ZN => n3396);
   U14745 : OAI22_X1 port map( A1 => n17948, A2 => n18016, B1 => n17947, B2 => 
                           n17081, ZN => n3397);
   U14746 : OAI22_X1 port map( A1 => n17949, A2 => n18019, B1 => n17947, B2 => 
                           n17082, ZN => n3398);
   U14747 : OAI22_X1 port map( A1 => n17949, A2 => n18022, B1 => n17947, B2 => 
                           n17083, ZN => n3399);
   U14748 : OAI22_X1 port map( A1 => n17949, A2 => n18025, B1 => n17947, B2 => 
                           n17084, ZN => n3400);
   U14749 : OAI22_X1 port map( A1 => n17949, A2 => n18028, B1 => n17947, B2 => 
                           n17085, ZN => n3401);
   U14750 : OAI22_X1 port map( A1 => n17949, A2 => n18031, B1 => n17947, B2 => 
                           n17086, ZN => n3402);
   U14751 : OAI22_X1 port map( A1 => n17950, A2 => n18034, B1 => n17947, B2 => 
                           n17087, ZN => n3403);
   U14752 : OAI22_X1 port map( A1 => n17950, A2 => n18037, B1 => n17947, B2 => 
                           n17088, ZN => n3404);
   U14753 : OAI22_X1 port map( A1 => n17950, A2 => n18040, B1 => n14643, B2 => 
                           n17089, ZN => n3405);
   U14754 : OAI22_X1 port map( A1 => n17950, A2 => n18043, B1 => n14643, B2 => 
                           n17090, ZN => n3406);
   U14755 : OAI22_X1 port map( A1 => n17950, A2 => n18046, B1 => n14643, B2 => 
                           n17091, ZN => n3407);
   U14756 : OAI22_X1 port map( A1 => n17951, A2 => n18049, B1 => n17947, B2 => 
                           n17092, ZN => n3408);
   U14757 : OAI22_X1 port map( A1 => n17951, A2 => n18052, B1 => n17947, B2 => 
                           n17093, ZN => n3409);
   U14758 : OAI22_X1 port map( A1 => n17951, A2 => n18055, B1 => n17947, B2 => 
                           n17094, ZN => n3410);
   U14759 : OAI22_X1 port map( A1 => n17951, A2 => n18058, B1 => n17947, B2 => 
                           n17095, ZN => n3411);
   U14760 : OAI22_X1 port map( A1 => n17951, A2 => n18061, B1 => n17947, B2 => 
                           n17096, ZN => n3412);
   U14761 : OAI22_X1 port map( A1 => n17952, A2 => n18064, B1 => n17947, B2 => 
                           n17097, ZN => n3413);
   U14762 : OAI22_X1 port map( A1 => n17952, A2 => n18067, B1 => n17947, B2 => 
                           n17098, ZN => n3414);
   U14763 : OAI22_X1 port map( A1 => n17952, A2 => n18070, B1 => n17947, B2 => 
                           n17099, ZN => n3415);
   U14764 : OAI22_X1 port map( A1 => n17952, A2 => n18073, B1 => n17947, B2 => 
                           n17100, ZN => n3416);
   U14765 : OAI22_X1 port map( A1 => n17912, A2 => n18004, B1 => n17911, B2 => 
                           n17101, ZN => n3265);
   U14766 : OAI22_X1 port map( A1 => n17912, A2 => n18007, B1 => n17911, B2 => 
                           n17102, ZN => n3266);
   U14767 : OAI22_X1 port map( A1 => n17912, A2 => n18010, B1 => n17911, B2 => 
                           n17103, ZN => n3267);
   U14768 : OAI22_X1 port map( A1 => n17912, A2 => n18013, B1 => n17911, B2 => 
                           n17104, ZN => n3268);
   U14769 : OAI22_X1 port map( A1 => n17912, A2 => n18016, B1 => n17911, B2 => 
                           n17105, ZN => n3269);
   U14770 : OAI22_X1 port map( A1 => n17913, A2 => n18019, B1 => n17911, B2 => 
                           n17106, ZN => n3270);
   U14771 : OAI22_X1 port map( A1 => n17913, A2 => n18022, B1 => n17911, B2 => 
                           n17107, ZN => n3271);
   U14772 : OAI22_X1 port map( A1 => n17913, A2 => n18025, B1 => n17911, B2 => 
                           n17108, ZN => n3272);
   U14773 : OAI22_X1 port map( A1 => n17913, A2 => n18028, B1 => n17911, B2 => 
                           n17109, ZN => n3273);
   U14774 : OAI22_X1 port map( A1 => n17913, A2 => n18031, B1 => n17911, B2 => 
                           n17110, ZN => n3274);
   U14775 : OAI22_X1 port map( A1 => n17914, A2 => n18034, B1 => n17911, B2 => 
                           n17111, ZN => n3275);
   U14776 : OAI22_X1 port map( A1 => n17914, A2 => n18037, B1 => n17911, B2 => 
                           n17112, ZN => n3276);
   U14777 : OAI22_X1 port map( A1 => n17914, A2 => n18040, B1 => n14651, B2 => 
                           n17113, ZN => n3277);
   U14778 : OAI22_X1 port map( A1 => n17914, A2 => n18043, B1 => n14651, B2 => 
                           n17114, ZN => n3278);
   U14779 : OAI22_X1 port map( A1 => n17914, A2 => n18046, B1 => n14651, B2 => 
                           n17115, ZN => n3279);
   U14780 : OAI22_X1 port map( A1 => n17915, A2 => n18049, B1 => n17911, B2 => 
                           n17116, ZN => n3280);
   U14781 : OAI22_X1 port map( A1 => n17915, A2 => n18052, B1 => n17911, B2 => 
                           n17117, ZN => n3281);
   U14782 : OAI22_X1 port map( A1 => n17915, A2 => n18055, B1 => n17911, B2 => 
                           n17118, ZN => n3282);
   U14783 : OAI22_X1 port map( A1 => n17915, A2 => n18058, B1 => n17911, B2 => 
                           n17119, ZN => n3283);
   U14784 : OAI22_X1 port map( A1 => n17915, A2 => n18061, B1 => n17911, B2 => 
                           n17120, ZN => n3284);
   U14785 : OAI22_X1 port map( A1 => n17916, A2 => n18064, B1 => n17911, B2 => 
                           n17121, ZN => n3285);
   U14786 : OAI22_X1 port map( A1 => n17916, A2 => n18067, B1 => n17911, B2 => 
                           n17122, ZN => n3286);
   U14787 : OAI22_X1 port map( A1 => n17916, A2 => n18070, B1 => n17911, B2 => 
                           n17123, ZN => n3287);
   U14788 : OAI22_X1 port map( A1 => n17916, A2 => n18073, B1 => n17911, B2 => 
                           n17124, ZN => n3288);
   U14789 : OAI22_X1 port map( A1 => n17876, A2 => n18005, B1 => n17875, B2 => 
                           n17125, ZN => n3137);
   U14790 : OAI22_X1 port map( A1 => n17876, A2 => n18008, B1 => n17875, B2 => 
                           n17126, ZN => n3138);
   U14791 : OAI22_X1 port map( A1 => n17876, A2 => n18011, B1 => n17875, B2 => 
                           n17127, ZN => n3139);
   U14792 : OAI22_X1 port map( A1 => n17876, A2 => n18014, B1 => n17875, B2 => 
                           n17128, ZN => n3140);
   U14793 : OAI22_X1 port map( A1 => n17876, A2 => n18017, B1 => n17875, B2 => 
                           n17129, ZN => n3141);
   U14794 : OAI22_X1 port map( A1 => n17877, A2 => n18020, B1 => n17875, B2 => 
                           n17130, ZN => n3142);
   U14795 : OAI22_X1 port map( A1 => n17877, A2 => n18023, B1 => n17875, B2 => 
                           n17131, ZN => n3143);
   U14796 : OAI22_X1 port map( A1 => n17877, A2 => n18026, B1 => n17875, B2 => 
                           n17132, ZN => n3144);
   U14797 : OAI22_X1 port map( A1 => n17877, A2 => n18029, B1 => n17875, B2 => 
                           n17133, ZN => n3145);
   U14798 : OAI22_X1 port map( A1 => n17877, A2 => n18032, B1 => n17875, B2 => 
                           n17134, ZN => n3146);
   U14799 : OAI22_X1 port map( A1 => n17878, A2 => n18035, B1 => n17875, B2 => 
                           n17135, ZN => n3147);
   U14800 : OAI22_X1 port map( A1 => n17878, A2 => n18038, B1 => n17875, B2 => 
                           n17136, ZN => n3148);
   U14801 : OAI22_X1 port map( A1 => n17878, A2 => n18041, B1 => n14655, B2 => 
                           n17137, ZN => n3149);
   U14802 : OAI22_X1 port map( A1 => n17878, A2 => n18044, B1 => n14655, B2 => 
                           n17138, ZN => n3150);
   U14803 : OAI22_X1 port map( A1 => n17878, A2 => n18047, B1 => n14655, B2 => 
                           n17139, ZN => n3151);
   U14804 : OAI22_X1 port map( A1 => n17879, A2 => n18050, B1 => n17875, B2 => 
                           n17140, ZN => n3152);
   U14805 : OAI22_X1 port map( A1 => n17879, A2 => n18053, B1 => n17875, B2 => 
                           n17141, ZN => n3153);
   U14806 : OAI22_X1 port map( A1 => n17879, A2 => n18056, B1 => n17875, B2 => 
                           n17142, ZN => n3154);
   U14807 : OAI22_X1 port map( A1 => n17879, A2 => n18059, B1 => n17875, B2 => 
                           n17143, ZN => n3155);
   U14808 : OAI22_X1 port map( A1 => n17879, A2 => n18062, B1 => n17875, B2 => 
                           n17144, ZN => n3156);
   U14809 : OAI22_X1 port map( A1 => n17880, A2 => n18065, B1 => n17875, B2 => 
                           n17145, ZN => n3157);
   U14810 : OAI22_X1 port map( A1 => n17880, A2 => n18068, B1 => n17875, B2 => 
                           n17146, ZN => n3158);
   U14811 : OAI22_X1 port map( A1 => n17880, A2 => n18071, B1 => n17875, B2 => 
                           n17147, ZN => n3159);
   U14812 : OAI22_X1 port map( A1 => n17880, A2 => n18074, B1 => n17875, B2 => 
                           n17148, ZN => n3160);
   U14813 : OAI22_X1 port map( A1 => n17804, A2 => n18005, B1 => n17803, B2 => 
                           n17149, ZN => n2881);
   U14814 : OAI22_X1 port map( A1 => n17804, A2 => n18008, B1 => n17803, B2 => 
                           n17150, ZN => n2882);
   U14815 : OAI22_X1 port map( A1 => n17804, A2 => n18011, B1 => n17803, B2 => 
                           n17151, ZN => n2883);
   U14816 : OAI22_X1 port map( A1 => n17804, A2 => n18014, B1 => n17803, B2 => 
                           n17152, ZN => n2884);
   U14817 : OAI22_X1 port map( A1 => n17804, A2 => n18017, B1 => n17803, B2 => 
                           n17153, ZN => n2885);
   U14818 : OAI22_X1 port map( A1 => n17805, A2 => n18020, B1 => n17803, B2 => 
                           n17154, ZN => n2886);
   U14819 : OAI22_X1 port map( A1 => n17805, A2 => n18023, B1 => n17803, B2 => 
                           n17155, ZN => n2887);
   U14820 : OAI22_X1 port map( A1 => n17805, A2 => n18026, B1 => n17803, B2 => 
                           n17156, ZN => n2888);
   U14821 : OAI22_X1 port map( A1 => n17805, A2 => n18029, B1 => n17803, B2 => 
                           n17157, ZN => n2889);
   U14822 : OAI22_X1 port map( A1 => n17805, A2 => n18032, B1 => n17803, B2 => 
                           n17158, ZN => n2890);
   U14823 : OAI22_X1 port map( A1 => n17806, A2 => n18035, B1 => n17803, B2 => 
                           n17159, ZN => n2891);
   U14824 : OAI22_X1 port map( A1 => n17806, A2 => n18038, B1 => n17803, B2 => 
                           n17160, ZN => n2892);
   U14825 : OAI22_X1 port map( A1 => n17806, A2 => n18041, B1 => n14664, B2 => 
                           n17161, ZN => n2893);
   U14826 : OAI22_X1 port map( A1 => n17806, A2 => n18044, B1 => n14664, B2 => 
                           n17162, ZN => n2894);
   U14827 : OAI22_X1 port map( A1 => n17806, A2 => n18047, B1 => n14664, B2 => 
                           n17163, ZN => n2895);
   U14828 : OAI22_X1 port map( A1 => n17807, A2 => n18050, B1 => n17803, B2 => 
                           n17164, ZN => n2896);
   U14829 : OAI22_X1 port map( A1 => n17807, A2 => n18053, B1 => n17803, B2 => 
                           n17165, ZN => n2897);
   U14830 : OAI22_X1 port map( A1 => n17807, A2 => n18056, B1 => n17803, B2 => 
                           n17166, ZN => n2898);
   U14831 : OAI22_X1 port map( A1 => n17807, A2 => n18059, B1 => n17803, B2 => 
                           n17167, ZN => n2899);
   U14832 : OAI22_X1 port map( A1 => n17807, A2 => n18062, B1 => n17803, B2 => 
                           n17168, ZN => n2900);
   U14833 : OAI22_X1 port map( A1 => n17808, A2 => n18065, B1 => n17803, B2 => 
                           n17169, ZN => n2901);
   U14834 : OAI22_X1 port map( A1 => n17808, A2 => n18068, B1 => n17803, B2 => 
                           n17170, ZN => n2902);
   U14835 : OAI22_X1 port map( A1 => n17808, A2 => n18071, B1 => n17803, B2 => 
                           n17171, ZN => n2903);
   U14836 : OAI22_X1 port map( A1 => n17808, A2 => n18074, B1 => n17803, B2 => 
                           n17172, ZN => n2904);
   U14837 : OAI22_X1 port map( A1 => n17786, A2 => n18006, B1 => n17785, B2 => 
                           n17173, ZN => n2817);
   U14838 : OAI22_X1 port map( A1 => n17786, A2 => n18009, B1 => n17785, B2 => 
                           n17174, ZN => n2818);
   U14839 : OAI22_X1 port map( A1 => n17786, A2 => n18012, B1 => n17785, B2 => 
                           n17175, ZN => n2819);
   U14840 : OAI22_X1 port map( A1 => n17786, A2 => n18015, B1 => n17785, B2 => 
                           n17176, ZN => n2820);
   U14841 : OAI22_X1 port map( A1 => n17786, A2 => n18018, B1 => n17785, B2 => 
                           n17177, ZN => n2821);
   U14842 : OAI22_X1 port map( A1 => n17787, A2 => n18021, B1 => n17785, B2 => 
                           n17178, ZN => n2822);
   U14843 : OAI22_X1 port map( A1 => n17787, A2 => n18024, B1 => n17785, B2 => 
                           n17179, ZN => n2823);
   U14844 : OAI22_X1 port map( A1 => n17787, A2 => n18027, B1 => n17785, B2 => 
                           n17180, ZN => n2824);
   U14845 : OAI22_X1 port map( A1 => n17787, A2 => n18030, B1 => n17785, B2 => 
                           n17181, ZN => n2825);
   U14846 : OAI22_X1 port map( A1 => n17787, A2 => n18033, B1 => n17785, B2 => 
                           n17182, ZN => n2826);
   U14847 : OAI22_X1 port map( A1 => n17788, A2 => n18036, B1 => n17785, B2 => 
                           n17183, ZN => n2827);
   U14848 : OAI22_X1 port map( A1 => n17788, A2 => n18039, B1 => n17785, B2 => 
                           n17184, ZN => n2828);
   U14849 : OAI22_X1 port map( A1 => n17788, A2 => n18042, B1 => n14666, B2 => 
                           n17185, ZN => n2829);
   U14850 : OAI22_X1 port map( A1 => n17788, A2 => n18045, B1 => n14666, B2 => 
                           n17186, ZN => n2830);
   U14851 : OAI22_X1 port map( A1 => n17788, A2 => n18048, B1 => n14666, B2 => 
                           n17187, ZN => n2831);
   U14852 : OAI22_X1 port map( A1 => n17789, A2 => n18051, B1 => n17785, B2 => 
                           n17188, ZN => n2832);
   U14853 : OAI22_X1 port map( A1 => n17789, A2 => n18054, B1 => n17785, B2 => 
                           n17189, ZN => n2833);
   U14854 : OAI22_X1 port map( A1 => n17789, A2 => n18057, B1 => n17785, B2 => 
                           n17190, ZN => n2834);
   U14855 : OAI22_X1 port map( A1 => n17789, A2 => n18060, B1 => n17785, B2 => 
                           n17191, ZN => n2835);
   U14856 : OAI22_X1 port map( A1 => n17789, A2 => n18063, B1 => n17785, B2 => 
                           n17192, ZN => n2836);
   U14857 : OAI22_X1 port map( A1 => n17790, A2 => n18066, B1 => n17785, B2 => 
                           n17193, ZN => n2837);
   U14858 : OAI22_X1 port map( A1 => n17790, A2 => n18069, B1 => n17785, B2 => 
                           n17194, ZN => n2838);
   U14859 : OAI22_X1 port map( A1 => n17790, A2 => n18072, B1 => n17785, B2 => 
                           n17195, ZN => n2839);
   U14860 : OAI22_X1 port map( A1 => n17790, A2 => n18075, B1 => n17785, B2 => 
                           n17196, ZN => n2840);
   U14861 : OAI22_X1 port map( A1 => n17750, A2 => n18006, B1 => n17749, B2 => 
                           n17197, ZN => n2689);
   U14862 : OAI22_X1 port map( A1 => n17750, A2 => n18009, B1 => n17749, B2 => 
                           n17198, ZN => n2690);
   U14863 : OAI22_X1 port map( A1 => n17750, A2 => n18012, B1 => n17749, B2 => 
                           n17199, ZN => n2691);
   U14864 : OAI22_X1 port map( A1 => n17750, A2 => n18015, B1 => n17749, B2 => 
                           n17200, ZN => n2692);
   U14865 : OAI22_X1 port map( A1 => n17750, A2 => n18018, B1 => n17749, B2 => 
                           n17201, ZN => n2693);
   U14866 : OAI22_X1 port map( A1 => n17751, A2 => n18021, B1 => n17749, B2 => 
                           n17202, ZN => n2694);
   U14867 : OAI22_X1 port map( A1 => n17751, A2 => n18024, B1 => n17749, B2 => 
                           n17203, ZN => n2695);
   U14868 : OAI22_X1 port map( A1 => n17751, A2 => n18027, B1 => n17749, B2 => 
                           n17204, ZN => n2696);
   U14869 : OAI22_X1 port map( A1 => n17751, A2 => n18030, B1 => n17749, B2 => 
                           n17205, ZN => n2697);
   U14870 : OAI22_X1 port map( A1 => n17751, A2 => n18033, B1 => n17749, B2 => 
                           n17206, ZN => n2698);
   U14871 : OAI22_X1 port map( A1 => n17752, A2 => n18036, B1 => n17749, B2 => 
                           n17207, ZN => n2699);
   U14872 : OAI22_X1 port map( A1 => n17752, A2 => n18039, B1 => n17749, B2 => 
                           n17208, ZN => n2700);
   U14873 : OAI22_X1 port map( A1 => n17752, A2 => n18042, B1 => n14671, B2 => 
                           n17209, ZN => n2701);
   U14874 : OAI22_X1 port map( A1 => n17752, A2 => n18045, B1 => n14671, B2 => 
                           n17210, ZN => n2702);
   U14875 : OAI22_X1 port map( A1 => n17752, A2 => n18048, B1 => n14671, B2 => 
                           n17211, ZN => n2703);
   U14876 : OAI22_X1 port map( A1 => n17753, A2 => n18051, B1 => n17749, B2 => 
                           n17212, ZN => n2704);
   U14877 : OAI22_X1 port map( A1 => n17753, A2 => n18054, B1 => n17749, B2 => 
                           n17213, ZN => n2705);
   U14878 : OAI22_X1 port map( A1 => n17753, A2 => n18057, B1 => n17749, B2 => 
                           n17214, ZN => n2706);
   U14879 : OAI22_X1 port map( A1 => n17753, A2 => n18060, B1 => n17749, B2 => 
                           n17215, ZN => n2707);
   U14880 : OAI22_X1 port map( A1 => n17753, A2 => n18063, B1 => n17749, B2 => 
                           n17216, ZN => n2708);
   U14881 : OAI22_X1 port map( A1 => n17754, A2 => n18066, B1 => n17749, B2 => 
                           n17217, ZN => n2709);
   U14882 : OAI22_X1 port map( A1 => n17754, A2 => n18069, B1 => n17749, B2 => 
                           n17218, ZN => n2710);
   U14883 : OAI22_X1 port map( A1 => n17754, A2 => n18072, B1 => n17749, B2 => 
                           n17219, ZN => n2711);
   U14884 : OAI22_X1 port map( A1 => n17754, A2 => n18075, B1 => n17749, B2 => 
                           n17220, ZN => n2712);
   U14885 : OAI22_X1 port map( A1 => n17858, A2 => n18005, B1 => n17857, B2 => 
                           n17221, ZN => n3073);
   U14886 : OAI22_X1 port map( A1 => n17858, A2 => n18008, B1 => n17857, B2 => 
                           n17222, ZN => n3074);
   U14887 : OAI22_X1 port map( A1 => n17858, A2 => n18011, B1 => n17857, B2 => 
                           n17223, ZN => n3075);
   U14888 : OAI22_X1 port map( A1 => n17858, A2 => n18014, B1 => n17857, B2 => 
                           n17224, ZN => n3076);
   U14889 : OAI22_X1 port map( A1 => n17858, A2 => n18017, B1 => n17857, B2 => 
                           n17225, ZN => n3077);
   U14890 : OAI22_X1 port map( A1 => n17859, A2 => n18020, B1 => n17857, B2 => 
                           n17226, ZN => n3078);
   U14891 : OAI22_X1 port map( A1 => n17859, A2 => n18023, B1 => n17857, B2 => 
                           n17227, ZN => n3079);
   U14892 : OAI22_X1 port map( A1 => n17859, A2 => n18026, B1 => n17857, B2 => 
                           n17228, ZN => n3080);
   U14893 : OAI22_X1 port map( A1 => n17859, A2 => n18029, B1 => n17857, B2 => 
                           n17229, ZN => n3081);
   U14894 : OAI22_X1 port map( A1 => n17859, A2 => n18032, B1 => n17857, B2 => 
                           n17230, ZN => n3082);
   U14895 : OAI22_X1 port map( A1 => n17860, A2 => n18035, B1 => n17857, B2 => 
                           n17231, ZN => n3083);
   U14896 : OAI22_X1 port map( A1 => n17860, A2 => n18038, B1 => n17857, B2 => 
                           n17232, ZN => n3084);
   U14897 : OAI22_X1 port map( A1 => n17860, A2 => n18041, B1 => n14657, B2 => 
                           n17233, ZN => n3085);
   U14898 : OAI22_X1 port map( A1 => n17860, A2 => n18044, B1 => n14657, B2 => 
                           n17234, ZN => n3086);
   U14899 : OAI22_X1 port map( A1 => n17860, A2 => n18047, B1 => n14657, B2 => 
                           n17235, ZN => n3087);
   U14900 : OAI22_X1 port map( A1 => n17861, A2 => n18050, B1 => n17857, B2 => 
                           n17236, ZN => n3088);
   U14901 : OAI22_X1 port map( A1 => n17861, A2 => n18053, B1 => n17857, B2 => 
                           n17237, ZN => n3089);
   U14902 : OAI22_X1 port map( A1 => n17861, A2 => n18056, B1 => n17857, B2 => 
                           n17238, ZN => n3090);
   U14903 : OAI22_X1 port map( A1 => n17861, A2 => n18059, B1 => n17857, B2 => 
                           n17239, ZN => n3091);
   U14904 : OAI22_X1 port map( A1 => n17861, A2 => n18062, B1 => n17857, B2 => 
                           n17240, ZN => n3092);
   U14905 : OAI22_X1 port map( A1 => n17862, A2 => n18065, B1 => n17857, B2 => 
                           n17241, ZN => n3093);
   U14906 : OAI22_X1 port map( A1 => n17862, A2 => n18068, B1 => n17857, B2 => 
                           n17242, ZN => n3094);
   U14907 : OAI22_X1 port map( A1 => n17862, A2 => n18071, B1 => n17857, B2 => 
                           n17243, ZN => n3095);
   U14908 : OAI22_X1 port map( A1 => n17862, A2 => n18074, B1 => n17857, B2 => 
                           n17244, ZN => n3096);
   U14909 : OAI22_X1 port map( A1 => n17849, A2 => n18005, B1 => n17848, B2 => 
                           n16737, ZN => n3041);
   U14910 : OAI22_X1 port map( A1 => n17849, A2 => n18008, B1 => n17848, B2 => 
                           n16738, ZN => n3042);
   U14911 : OAI22_X1 port map( A1 => n17849, A2 => n18011, B1 => n17848, B2 => 
                           n16739, ZN => n3043);
   U14912 : OAI22_X1 port map( A1 => n17849, A2 => n18014, B1 => n17848, B2 => 
                           n16740, ZN => n3044);
   U14913 : OAI22_X1 port map( A1 => n17849, A2 => n18017, B1 => n17848, B2 => 
                           n16741, ZN => n3045);
   U14914 : OAI22_X1 port map( A1 => n17850, A2 => n18020, B1 => n17848, B2 => 
                           n16742, ZN => n3046);
   U14915 : OAI22_X1 port map( A1 => n17850, A2 => n18023, B1 => n17848, B2 => 
                           n16743, ZN => n3047);
   U14916 : OAI22_X1 port map( A1 => n17850, A2 => n18026, B1 => n17848, B2 => 
                           n16744, ZN => n3048);
   U14917 : OAI22_X1 port map( A1 => n17850, A2 => n18029, B1 => n17848, B2 => 
                           n16745, ZN => n3049);
   U14918 : OAI22_X1 port map( A1 => n17850, A2 => n18032, B1 => n17848, B2 => 
                           n16746, ZN => n3050);
   U14919 : OAI22_X1 port map( A1 => n17851, A2 => n18035, B1 => n17848, B2 => 
                           n16747, ZN => n3051);
   U14920 : OAI22_X1 port map( A1 => n17851, A2 => n18038, B1 => n17848, B2 => 
                           n16748, ZN => n3052);
   U14921 : OAI22_X1 port map( A1 => n17851, A2 => n18041, B1 => n14659, B2 => 
                           n16633, ZN => n3053);
   U14922 : OAI22_X1 port map( A1 => n17851, A2 => n18044, B1 => n14659, B2 => 
                           n16634, ZN => n3054);
   U14923 : OAI22_X1 port map( A1 => n17851, A2 => n18047, B1 => n14659, B2 => 
                           n16635, ZN => n3055);
   U14924 : OAI22_X1 port map( A1 => n17852, A2 => n18050, B1 => n17848, B2 => 
                           n16636, ZN => n3056);
   U14925 : OAI22_X1 port map( A1 => n17852, A2 => n18053, B1 => n17848, B2 => 
                           n16637, ZN => n3057);
   U14926 : OAI22_X1 port map( A1 => n17852, A2 => n18056, B1 => n17848, B2 => 
                           n16638, ZN => n3058);
   U14927 : OAI22_X1 port map( A1 => n17852, A2 => n18059, B1 => n17848, B2 => 
                           n16639, ZN => n3059);
   U14928 : OAI22_X1 port map( A1 => n17852, A2 => n18062, B1 => n17848, B2 => 
                           n16640, ZN => n3060);
   U14929 : OAI22_X1 port map( A1 => n17853, A2 => n18065, B1 => n17848, B2 => 
                           n16641, ZN => n3061);
   U14930 : OAI22_X1 port map( A1 => n17853, A2 => n18068, B1 => n17848, B2 => 
                           n16642, ZN => n3062);
   U14931 : OAI22_X1 port map( A1 => n17853, A2 => n18071, B1 => n17848, B2 => 
                           n16643, ZN => n3063);
   U14932 : OAI22_X1 port map( A1 => n17853, A2 => n18074, B1 => n17848, B2 => 
                           n16644, ZN => n3064);
   U14933 : NOR2_X1 port map( A1 => n13570, A2 => n13571, ZN => n15963);
   U14934 : NOR2_X1 port map( A1 => n13566, A2 => n13567, ZN => n15310);
   U14935 : BUF_X1 port map( A => n15328, Z => n17615);
   U14936 : BUF_X1 port map( A => n14675, Z => n17717);
   U14937 : BUF_X1 port map( A => n15328, Z => n17616);
   U14938 : BUF_X1 port map( A => n15328, Z => n17617);
   U14939 : BUF_X1 port map( A => n14675, Z => n17718);
   U14940 : BUF_X1 port map( A => n14675, Z => n17719);
   U14941 : BUF_X1 port map( A => n13559, Z => n18111);
   U14942 : BUF_X1 port map( A => n13559, Z => n18110);
   U14943 : BUF_X1 port map( A => n13559, Z => n18109);
   U14944 : BUF_X1 port map( A => n14629, Z => n18004);
   U14945 : BUF_X1 port map( A => n14628, Z => n18007);
   U14946 : BUF_X1 port map( A => n14627, Z => n18010);
   U14947 : BUF_X1 port map( A => n14626, Z => n18013);
   U14948 : BUF_X1 port map( A => n14625, Z => n18016);
   U14949 : BUF_X1 port map( A => n14624, Z => n18019);
   U14950 : BUF_X1 port map( A => n14623, Z => n18022);
   U14951 : BUF_X1 port map( A => n14622, Z => n18025);
   U14952 : BUF_X1 port map( A => n14629, Z => n18005);
   U14953 : BUF_X1 port map( A => n14628, Z => n18008);
   U14954 : BUF_X1 port map( A => n14627, Z => n18011);
   U14955 : BUF_X1 port map( A => n14626, Z => n18014);
   U14956 : BUF_X1 port map( A => n14625, Z => n18017);
   U14957 : BUF_X1 port map( A => n14624, Z => n18020);
   U14958 : BUF_X1 port map( A => n14623, Z => n18023);
   U14959 : BUF_X1 port map( A => n14622, Z => n18026);
   U14960 : BUF_X1 port map( A => n14621, Z => n18028);
   U14961 : BUF_X1 port map( A => n14620, Z => n18031);
   U14962 : BUF_X1 port map( A => n14619, Z => n18034);
   U14963 : BUF_X1 port map( A => n14618, Z => n18037);
   U14964 : BUF_X1 port map( A => n14617, Z => n18040);
   U14965 : BUF_X1 port map( A => n14616, Z => n18043);
   U14966 : BUF_X1 port map( A => n14615, Z => n18046);
   U14967 : BUF_X1 port map( A => n14614, Z => n18049);
   U14968 : BUF_X1 port map( A => n14613, Z => n18052);
   U14969 : BUF_X1 port map( A => n14612, Z => n18055);
   U14970 : BUF_X1 port map( A => n14611, Z => n18058);
   U14971 : BUF_X1 port map( A => n14610, Z => n18061);
   U14972 : BUF_X1 port map( A => n14609, Z => n18064);
   U14973 : BUF_X1 port map( A => n14608, Z => n18067);
   U14974 : BUF_X1 port map( A => n14607, Z => n18070);
   U14975 : BUF_X1 port map( A => n14606, Z => n18073);
   U14976 : BUF_X1 port map( A => n14605, Z => n18076);
   U14977 : BUF_X1 port map( A => n14604, Z => n18079);
   U14978 : BUF_X1 port map( A => n14603, Z => n18082);
   U14979 : BUF_X1 port map( A => n14602, Z => n18085);
   U14980 : BUF_X1 port map( A => n14601, Z => n18088);
   U14981 : BUF_X1 port map( A => n14600, Z => n18091);
   U14982 : BUF_X1 port map( A => n14599, Z => n18094);
   U14983 : BUF_X1 port map( A => n14597, Z => n18106);
   U14984 : BUF_X1 port map( A => n14621, Z => n18029);
   U14985 : BUF_X1 port map( A => n14620, Z => n18032);
   U14986 : BUF_X1 port map( A => n14619, Z => n18035);
   U14987 : BUF_X1 port map( A => n14618, Z => n18038);
   U14988 : BUF_X1 port map( A => n14617, Z => n18041);
   U14989 : BUF_X1 port map( A => n14616, Z => n18044);
   U14990 : BUF_X1 port map( A => n14615, Z => n18047);
   U14991 : BUF_X1 port map( A => n14614, Z => n18050);
   U14992 : BUF_X1 port map( A => n14613, Z => n18053);
   U14993 : BUF_X1 port map( A => n14612, Z => n18056);
   U14994 : BUF_X1 port map( A => n14611, Z => n18059);
   U14995 : BUF_X1 port map( A => n14610, Z => n18062);
   U14996 : BUF_X1 port map( A => n14609, Z => n18065);
   U14997 : BUF_X1 port map( A => n14608, Z => n18068);
   U14998 : BUF_X1 port map( A => n14607, Z => n18071);
   U14999 : BUF_X1 port map( A => n14606, Z => n18074);
   U15000 : BUF_X1 port map( A => n14605, Z => n18077);
   U15001 : BUF_X1 port map( A => n14604, Z => n18080);
   U15002 : BUF_X1 port map( A => n14603, Z => n18083);
   U15003 : BUF_X1 port map( A => n14602, Z => n18086);
   U15004 : BUF_X1 port map( A => n14601, Z => n18089);
   U15005 : BUF_X1 port map( A => n14600, Z => n18092);
   U15006 : BUF_X1 port map( A => n14599, Z => n18095);
   U15007 : BUF_X1 port map( A => n14597, Z => n18107);
   U15008 : BUF_X1 port map( A => n15328, Z => n17613);
   U15009 : BUF_X1 port map( A => n15328, Z => n17614);
   U15010 : BUF_X1 port map( A => n14675, Z => n17715);
   U15011 : BUF_X1 port map( A => n14675, Z => n17716);
   U15012 : BUF_X1 port map( A => n14632, Z => n18001);
   U15013 : BUF_X1 port map( A => n14632, Z => n18002);
   U15014 : BUF_X1 port map( A => n14629, Z => n18006);
   U15015 : BUF_X1 port map( A => n14628, Z => n18009);
   U15016 : BUF_X1 port map( A => n14627, Z => n18012);
   U15017 : BUF_X1 port map( A => n14626, Z => n18015);
   U15018 : BUF_X1 port map( A => n14625, Z => n18018);
   U15019 : BUF_X1 port map( A => n14624, Z => n18021);
   U15020 : BUF_X1 port map( A => n14623, Z => n18024);
   U15021 : BUF_X1 port map( A => n14622, Z => n18027);
   U15022 : BUF_X1 port map( A => n14621, Z => n18030);
   U15023 : BUF_X1 port map( A => n14620, Z => n18033);
   U15024 : BUF_X1 port map( A => n14619, Z => n18036);
   U15025 : BUF_X1 port map( A => n14618, Z => n18039);
   U15026 : BUF_X1 port map( A => n14617, Z => n18042);
   U15027 : BUF_X1 port map( A => n14616, Z => n18045);
   U15028 : BUF_X1 port map( A => n14615, Z => n18048);
   U15029 : BUF_X1 port map( A => n14614, Z => n18051);
   U15030 : BUF_X1 port map( A => n14613, Z => n18054);
   U15031 : BUF_X1 port map( A => n14612, Z => n18057);
   U15032 : BUF_X1 port map( A => n14611, Z => n18060);
   U15033 : BUF_X1 port map( A => n14610, Z => n18063);
   U15034 : BUF_X1 port map( A => n14609, Z => n18066);
   U15035 : BUF_X1 port map( A => n14608, Z => n18069);
   U15036 : BUF_X1 port map( A => n14607, Z => n18072);
   U15037 : BUF_X1 port map( A => n14606, Z => n18075);
   U15038 : BUF_X1 port map( A => n14605, Z => n18078);
   U15039 : BUF_X1 port map( A => n14604, Z => n18081);
   U15040 : BUF_X1 port map( A => n14603, Z => n18084);
   U15041 : BUF_X1 port map( A => n14602, Z => n18087);
   U15042 : BUF_X1 port map( A => n14601, Z => n18090);
   U15043 : BUF_X1 port map( A => n14600, Z => n18093);
   U15044 : BUF_X1 port map( A => n14599, Z => n18096);
   U15045 : BUF_X1 port map( A => n14597, Z => n18108);
   U15046 : BUF_X1 port map( A => n14632, Z => n18003);
   U15047 : NAND2_X1 port map( A1 => n15959, A2 => n15974, ZN => n15364);
   U15048 : NAND2_X1 port map( A1 => n15306, A2 => n15321, ZN => n14711);
   U15049 : NAND2_X1 port map( A1 => n15963, A2 => n15974, ZN => n15368);
   U15050 : NAND2_X1 port map( A1 => n15963, A2 => n15975, ZN => n15369);
   U15051 : NAND2_X1 port map( A1 => n15310, A2 => n15321, ZN => n14715);
   U15052 : NAND2_X1 port map( A1 => n15310, A2 => n15322, ZN => n14716);
   U15053 : NAND2_X1 port map( A1 => n15975, A2 => n15959, ZN => n15363);
   U15054 : NAND2_X1 port map( A1 => n15322, A2 => n15306, ZN => n14710);
   U15055 : NAND2_X1 port map( A1 => n15979, A2 => n15961, ZN => n15373);
   U15056 : NAND2_X1 port map( A1 => n15979, A2 => n15963, ZN => n15378);
   U15057 : NAND2_X1 port map( A1 => n15326, A2 => n15308, ZN => n14720);
   U15058 : NAND2_X1 port map( A1 => n15326, A2 => n15310, ZN => n14725);
   U15059 : NAND2_X1 port map( A1 => n15978, A2 => n15961, ZN => n15374);
   U15060 : NAND2_X1 port map( A1 => n15978, A2 => n15963, ZN => n15379);
   U15061 : NAND2_X1 port map( A1 => n15325, A2 => n15308, ZN => n14721);
   U15062 : NAND2_X1 port map( A1 => n15325, A2 => n15310, ZN => n14726);
   U15063 : NAND2_X1 port map( A1 => n15960, A2 => n15959, ZN => n15339);
   U15064 : NAND2_X1 port map( A1 => n15958, A2 => n15959, ZN => n15340);
   U15065 : NAND2_X1 port map( A1 => n15967, A2 => n15959, ZN => n15349);
   U15066 : NAND2_X1 port map( A1 => n15966, A2 => n15959, ZN => n15350);
   U15067 : NAND2_X1 port map( A1 => n15307, A2 => n15306, ZN => n14686);
   U15068 : NAND2_X1 port map( A1 => n15305, A2 => n15306, ZN => n14687);
   U15069 : NAND2_X1 port map( A1 => n15314, A2 => n15306, ZN => n14696);
   U15070 : NAND2_X1 port map( A1 => n15313, A2 => n15306, ZN => n14697);
   U15071 : NAND2_X1 port map( A1 => n15960, A2 => n15963, ZN => n15344);
   U15072 : NAND2_X1 port map( A1 => n15958, A2 => n15963, ZN => n15345);
   U15073 : NAND2_X1 port map( A1 => n15307, A2 => n15310, ZN => n14691);
   U15074 : NAND2_X1 port map( A1 => n15305, A2 => n15310, ZN => n14692);
   U15075 : NAND2_X1 port map( A1 => n15967, A2 => n15964, ZN => n15354);
   U15076 : NAND2_X1 port map( A1 => n15966, A2 => n15964, ZN => n15355);
   U15077 : NAND2_X1 port map( A1 => n15314, A2 => n15311, ZN => n14701);
   U15078 : NAND2_X1 port map( A1 => n15313, A2 => n15311, ZN => n14702);
   U15079 : AND2_X1 port map( A1 => n15961, A2 => n15975, ZN => n15360);
   U15080 : AND2_X1 port map( A1 => n15961, A2 => n15974, ZN => n15361);
   U15081 : AND2_X1 port map( A1 => n15964, A2 => n15974, ZN => n15365);
   U15082 : AND2_X1 port map( A1 => n15964, A2 => n15975, ZN => n15366);
   U15083 : AND2_X1 port map( A1 => n15308, A2 => n15322, ZN => n14707);
   U15084 : AND2_X1 port map( A1 => n15308, A2 => n15321, ZN => n14708);
   U15085 : AND2_X1 port map( A1 => n15311, A2 => n15321, ZN => n14712);
   U15086 : AND2_X1 port map( A1 => n15311, A2 => n15322, ZN => n14713);
   U15087 : AND2_X1 port map( A1 => n15979, A2 => n15959, ZN => n15370);
   U15088 : AND2_X1 port map( A1 => n15978, A2 => n15959, ZN => n15371);
   U15089 : AND2_X1 port map( A1 => n15326, A2 => n15306, ZN => n14717);
   U15090 : AND2_X1 port map( A1 => n15325, A2 => n15306, ZN => n14718);
   U15091 : AND2_X1 port map( A1 => n15967, A2 => n15963, ZN => n15351);
   U15092 : AND2_X1 port map( A1 => n15966, A2 => n15963, ZN => n15352);
   U15093 : AND2_X1 port map( A1 => n15314, A2 => n15310, ZN => n14698);
   U15094 : AND2_X1 port map( A1 => n15313, A2 => n15310, ZN => n14699);
   U15095 : AND2_X1 port map( A1 => n15979, A2 => n15964, ZN => n15375);
   U15096 : AND2_X1 port map( A1 => n15978, A2 => n15964, ZN => n15376);
   U15097 : AND2_X1 port map( A1 => n15326, A2 => n15311, ZN => n14722);
   U15098 : AND2_X1 port map( A1 => n15325, A2 => n15311, ZN => n14723);
   U15099 : AND2_X1 port map( A1 => n15960, A2 => n15961, ZN => n15336);
   U15100 : AND2_X1 port map( A1 => n15958, A2 => n15961, ZN => n15337);
   U15101 : AND2_X1 port map( A1 => n15960, A2 => n15964, ZN => n15341);
   U15102 : AND2_X1 port map( A1 => n15958, A2 => n15964, ZN => n15342);
   U15103 : AND2_X1 port map( A1 => n15967, A2 => n15961, ZN => n15346);
   U15104 : AND2_X1 port map( A1 => n15966, A2 => n15961, ZN => n15347);
   U15105 : AND2_X1 port map( A1 => n15307, A2 => n15308, ZN => n14683);
   U15106 : AND2_X1 port map( A1 => n15305, A2 => n15308, ZN => n14684);
   U15107 : AND2_X1 port map( A1 => n15307, A2 => n15311, ZN => n14688);
   U15108 : AND2_X1 port map( A1 => n15305, A2 => n15311, ZN => n14689);
   U15109 : AND2_X1 port map( A1 => n15314, A2 => n15308, ZN => n14693);
   U15110 : AND2_X1 port map( A1 => n15313, A2 => n15308, ZN => n14694);
   U15111 : BUF_X1 port map( A => n14674, Z => n17721);
   U15112 : OAI21_X1 port map( B1 => n14646, B2 => n14667, A => n18001, ZN => 
                           n14674);
   U15113 : INV_X1 port map( A => n14661, ZN => n17838);
   U15114 : OAI21_X1 port map( B1 => n14638, B2 => n14658, A => n18002, ZN => 
                           n14661);
   U15115 : INV_X1 port map( A => n14660, ZN => n17847);
   U15116 : OAI21_X1 port map( B1 => n14636, B2 => n14658, A => n18002, ZN => 
                           n14660);
   U15117 : INV_X1 port map( A => n14652, ZN => n17910);
   U15118 : OAI21_X1 port map( B1 => n14638, B2 => n14649, A => n18002, ZN => 
                           n14652);
   U15119 : INV_X1 port map( A => n14656, ZN => n17874);
   U15120 : OAI21_X1 port map( B1 => n14646, B2 => n14649, A => n18002, ZN => 
                           n14656);
   U15121 : INV_X1 port map( A => n14665, ZN => n17802);
   U15122 : OAI21_X1 port map( B1 => n14646, B2 => n14658, A => n18001, ZN => 
                           n14665);
   U15123 : INV_X1 port map( A => n14668, ZN => n17784);
   U15124 : OAI21_X1 port map( B1 => n14634, B2 => n14667, A => n18001, ZN => 
                           n14668);
   U15125 : INV_X1 port map( A => n14672, ZN => n17748);
   U15126 : OAI21_X1 port map( B1 => n14642, B2 => n14667, A => n18001, ZN => 
                           n14672);
   U15127 : INV_X1 port map( A => n14651, ZN => n17919);
   U15128 : OAI21_X1 port map( B1 => n14636, B2 => n14649, A => n18002, ZN => 
                           n14651);
   U15129 : INV_X1 port map( A => n14655, ZN => n17883);
   U15130 : OAI21_X1 port map( B1 => n14644, B2 => n14649, A => n18002, ZN => 
                           n14655);
   U15131 : INV_X1 port map( A => n14664, ZN => n17811);
   U15132 : OAI21_X1 port map( B1 => n14644, B2 => n14658, A => n18001, ZN => 
                           n14664);
   U15133 : INV_X1 port map( A => n14666, ZN => n17793);
   U15134 : OAI21_X1 port map( B1 => n14631, B2 => n14667, A => n18001, ZN => 
                           n14666);
   U15135 : INV_X1 port map( A => n14671, ZN => n17757);
   U15136 : OAI21_X1 port map( B1 => n14640, B2 => n14667, A => n18001, ZN => 
                           n14671);
   U15137 : INV_X1 port map( A => n14648, ZN => n17937);
   U15138 : OAI21_X1 port map( B1 => n14631, B2 => n14649, A => n18002, ZN => 
                           n14648);
   U15139 : INV_X1 port map( A => n14650, ZN => n17928);
   U15140 : OAI21_X1 port map( B1 => n14634, B2 => n14649, A => n18002, ZN => 
                           n14650);
   U15141 : INV_X1 port map( A => n14653, ZN => n17901);
   U15142 : OAI21_X1 port map( B1 => n14640, B2 => n14649, A => n18002, ZN => 
                           n14653);
   U15143 : INV_X1 port map( A => n14654, ZN => n17892);
   U15144 : OAI21_X1 port map( B1 => n14642, B2 => n14649, A => n18002, ZN => 
                           n14654);
   U15145 : INV_X1 port map( A => n14662, ZN => n17829);
   U15146 : OAI21_X1 port map( B1 => n14640, B2 => n14658, A => n18001, ZN => 
                           n14662);
   U15147 : INV_X1 port map( A => n14663, ZN => n17820);
   U15148 : OAI21_X1 port map( B1 => n14642, B2 => n14658, A => n18001, ZN => 
                           n14663);
   U15149 : INV_X1 port map( A => n14669, ZN => n17775);
   U15150 : OAI21_X1 port map( B1 => n14636, B2 => n14667, A => n18001, ZN => 
                           n14669);
   U15151 : INV_X1 port map( A => n14670, ZN => n17766);
   U15152 : OAI21_X1 port map( B1 => n14638, B2 => n14667, A => n18001, ZN => 
                           n14670);
   U15153 : INV_X1 port map( A => n14673, ZN => n17739);
   U15154 : OAI21_X1 port map( B1 => n14644, B2 => n14667, A => n18001, ZN => 
                           n14673);
   U15155 : INV_X1 port map( A => n14657, ZN => n17865);
   U15156 : OAI21_X1 port map( B1 => n14631, B2 => n14658, A => n18002, ZN => 
                           n14657);
   U15157 : INV_X1 port map( A => n14659, ZN => n17856);
   U15158 : OAI21_X1 port map( B1 => n14634, B2 => n14658, A => n18002, ZN => 
                           n14659);
   U15159 : INV_X1 port map( A => n14645, ZN => n17946);
   U15160 : OAI21_X1 port map( B1 => n14630, B2 => n14646, A => n18003, ZN => 
                           n14645);
   U15161 : INV_X1 port map( A => n14633, ZN => n18000);
   U15162 : OAI21_X1 port map( B1 => n14630, B2 => n14634, A => n18003, ZN => 
                           n14633);
   U15163 : INV_X1 port map( A => n14643, ZN => n17955);
   U15164 : OAI21_X1 port map( B1 => n14630, B2 => n14644, A => n18003, ZN => 
                           n14643);
   U15165 : INV_X1 port map( A => n14635, ZN => n17991);
   U15166 : OAI21_X1 port map( B1 => n14630, B2 => n14636, A => n18003, ZN => 
                           n14635);
   U15167 : INV_X1 port map( A => n14637, ZN => n17982);
   U15168 : OAI21_X1 port map( B1 => n14630, B2 => n14638, A => n18003, ZN => 
                           n14637);
   U15169 : INV_X1 port map( A => n14639, ZN => n17973);
   U15170 : OAI21_X1 port map( B1 => n14630, B2 => n14640, A => n18003, ZN => 
                           n14639);
   U15171 : INV_X1 port map( A => n14641, ZN => n17964);
   U15172 : OAI21_X1 port map( B1 => n14630, B2 => n14642, A => n18003, ZN => 
                           n14641);
   U15173 : AOI221_X1 port map( B1 => n17610, B2 => n12674, C1 => n17607, C2 =>
                           n12698, A => n15957, ZN => n15956);
   U15174 : OAI22_X1 port map( A1 => n16737, A2 => n17604, B1 => n17221, B2 => 
                           n17601, ZN => n15957);
   U15175 : AOI221_X1 port map( B1 => n17610, B2 => n12675, C1 => n17607, C2 =>
                           n12699, A => n15938, ZN => n15937);
   U15176 : OAI22_X1 port map( A1 => n16738, A2 => n17604, B1 => n17222, B2 => 
                           n17601, ZN => n15938);
   U15177 : AOI221_X1 port map( B1 => n17610, B2 => n12676, C1 => n17607, C2 =>
                           n12700, A => n15919, ZN => n15918);
   U15178 : OAI22_X1 port map( A1 => n16739, A2 => n17604, B1 => n17223, B2 => 
                           n17601, ZN => n15919);
   U15179 : AOI221_X1 port map( B1 => n17610, B2 => n12677, C1 => n17607, C2 =>
                           n12701, A => n15900, ZN => n15899);
   U15180 : OAI22_X1 port map( A1 => n16740, A2 => n17604, B1 => n17224, B2 => 
                           n17601, ZN => n15900);
   U15181 : AOI221_X1 port map( B1 => n17610, B2 => n12678, C1 => n17607, C2 =>
                           n12702, A => n15881, ZN => n15880);
   U15182 : OAI22_X1 port map( A1 => n16741, A2 => n17604, B1 => n17225, B2 => 
                           n17601, ZN => n15881);
   U15183 : AOI221_X1 port map( B1 => n17610, B2 => n12679, C1 => n17607, C2 =>
                           n12703, A => n15862, ZN => n15861);
   U15184 : OAI22_X1 port map( A1 => n16742, A2 => n17604, B1 => n17226, B2 => 
                           n17601, ZN => n15862);
   U15185 : AOI221_X1 port map( B1 => n17610, B2 => n12680, C1 => n17607, C2 =>
                           n12704, A => n15843, ZN => n15842);
   U15186 : OAI22_X1 port map( A1 => n16743, A2 => n17604, B1 => n17227, B2 => 
                           n17601, ZN => n15843);
   U15187 : AOI221_X1 port map( B1 => n17610, B2 => n12681, C1 => n17607, C2 =>
                           n12705, A => n15824, ZN => n15823);
   U15188 : OAI22_X1 port map( A1 => n16744, A2 => n17604, B1 => n17228, B2 => 
                           n17601, ZN => n15824);
   U15189 : AOI221_X1 port map( B1 => n17610, B2 => n12682, C1 => n17607, C2 =>
                           n12706, A => n15805, ZN => n15804);
   U15190 : OAI22_X1 port map( A1 => n16745, A2 => n17604, B1 => n17229, B2 => 
                           n17601, ZN => n15805);
   U15191 : AOI221_X1 port map( B1 => n17610, B2 => n12683, C1 => n17607, C2 =>
                           n12707, A => n15786, ZN => n15785);
   U15192 : OAI22_X1 port map( A1 => n16746, A2 => n17604, B1 => n17230, B2 => 
                           n17601, ZN => n15786);
   U15193 : AOI221_X1 port map( B1 => n17610, B2 => n12684, C1 => n17607, C2 =>
                           n12708, A => n15767, ZN => n15766);
   U15194 : OAI22_X1 port map( A1 => n16747, A2 => n17604, B1 => n17231, B2 => 
                           n17601, ZN => n15767);
   U15195 : AOI221_X1 port map( B1 => n17610, B2 => n12685, C1 => n17607, C2 =>
                           n12709, A => n15748, ZN => n15747);
   U15196 : OAI22_X1 port map( A1 => n16748, A2 => n17604, B1 => n17232, B2 => 
                           n17601, ZN => n15748);
   U15197 : AOI221_X1 port map( B1 => n17611, B2 => n12686, C1 => n17608, C2 =>
                           n12710, A => n15729, ZN => n15728);
   U15198 : OAI22_X1 port map( A1 => n16633, A2 => n17605, B1 => n17233, B2 => 
                           n17602, ZN => n15729);
   U15199 : AOI221_X1 port map( B1 => n17611, B2 => n12687, C1 => n17608, C2 =>
                           n12711, A => n15710, ZN => n15709);
   U15200 : OAI22_X1 port map( A1 => n16634, A2 => n17605, B1 => n17234, B2 => 
                           n17602, ZN => n15710);
   U15201 : AOI221_X1 port map( B1 => n17611, B2 => n12688, C1 => n17608, C2 =>
                           n12712, A => n15691, ZN => n15690);
   U15202 : OAI22_X1 port map( A1 => n16635, A2 => n17605, B1 => n17235, B2 => 
                           n17602, ZN => n15691);
   U15203 : AOI221_X1 port map( B1 => n17611, B2 => n12689, C1 => n17608, C2 =>
                           n12713, A => n15672, ZN => n15671);
   U15204 : OAI22_X1 port map( A1 => n16636, A2 => n17605, B1 => n17236, B2 => 
                           n17602, ZN => n15672);
   U15205 : AOI221_X1 port map( B1 => n17611, B2 => n12690, C1 => n17608, C2 =>
                           n12714, A => n15653, ZN => n15652);
   U15206 : OAI22_X1 port map( A1 => n16637, A2 => n17605, B1 => n17237, B2 => 
                           n17602, ZN => n15653);
   U15207 : AOI221_X1 port map( B1 => n17611, B2 => n12691, C1 => n17608, C2 =>
                           n12715, A => n15634, ZN => n15633);
   U15208 : OAI22_X1 port map( A1 => n16638, A2 => n17605, B1 => n17238, B2 => 
                           n17602, ZN => n15634);
   U15209 : AOI221_X1 port map( B1 => n17611, B2 => n12692, C1 => n17608, C2 =>
                           n12716, A => n15615, ZN => n15614);
   U15210 : OAI22_X1 port map( A1 => n16639, A2 => n17605, B1 => n17239, B2 => 
                           n17602, ZN => n15615);
   U15211 : AOI221_X1 port map( B1 => n17611, B2 => n12693, C1 => n17608, C2 =>
                           n12717, A => n15596, ZN => n15595);
   U15212 : OAI22_X1 port map( A1 => n16640, A2 => n17605, B1 => n17240, B2 => 
                           n17602, ZN => n15596);
   U15213 : AOI221_X1 port map( B1 => n17611, B2 => n12694, C1 => n17608, C2 =>
                           n12718, A => n15577, ZN => n15576);
   U15214 : OAI22_X1 port map( A1 => n16641, A2 => n17605, B1 => n17241, B2 => 
                           n17602, ZN => n15577);
   U15215 : AOI221_X1 port map( B1 => n17611, B2 => n12695, C1 => n17608, C2 =>
                           n12719, A => n15558, ZN => n15557);
   U15216 : OAI22_X1 port map( A1 => n16642, A2 => n17605, B1 => n17242, B2 => 
                           n17602, ZN => n15558);
   U15217 : AOI221_X1 port map( B1 => n17611, B2 => n12696, C1 => n17608, C2 =>
                           n12720, A => n15539, ZN => n15538);
   U15218 : OAI22_X1 port map( A1 => n16643, A2 => n17605, B1 => n17243, B2 => 
                           n17602, ZN => n15539);
   U15219 : AOI221_X1 port map( B1 => n17611, B2 => n12697, C1 => n17608, C2 =>
                           n12721, A => n15520, ZN => n15519);
   U15220 : OAI22_X1 port map( A1 => n16644, A2 => n17605, B1 => n17244, B2 => 
                           n17602, ZN => n15520);
   U15221 : AOI221_X1 port map( B1 => n17612, B2 => n12468, C1 => n17609, C2 =>
                           n12476, A => n15501, ZN => n15500);
   U15222 : OAI22_X1 port map( A1 => n16645, A2 => n17606, B1 => n16805, B2 => 
                           n17603, ZN => n15501);
   U15223 : AOI221_X1 port map( B1 => n17612, B2 => n12469, C1 => n17609, C2 =>
                           n12477, A => n15482, ZN => n15481);
   U15224 : OAI22_X1 port map( A1 => n16646, A2 => n17606, B1 => n16806, B2 => 
                           n17603, ZN => n15482);
   U15225 : AOI221_X1 port map( B1 => n17612, B2 => n12470, C1 => n17609, C2 =>
                           n12478, A => n15463, ZN => n15462);
   U15226 : OAI22_X1 port map( A1 => n16647, A2 => n17606, B1 => n16807, B2 => 
                           n17603, ZN => n15463);
   U15227 : AOI221_X1 port map( B1 => n17612, B2 => n12471, C1 => n17609, C2 =>
                           n12479, A => n15444, ZN => n15443);
   U15228 : OAI22_X1 port map( A1 => n16648, A2 => n17606, B1 => n16808, B2 => 
                           n17603, ZN => n15444);
   U15229 : AOI221_X1 port map( B1 => n17612, B2 => n12472, C1 => n17609, C2 =>
                           n12480, A => n15425, ZN => n15424);
   U15230 : OAI22_X1 port map( A1 => n16649, A2 => n17606, B1 => n16809, B2 => 
                           n17603, ZN => n15425);
   U15231 : AOI221_X1 port map( B1 => n17612, B2 => n12473, C1 => n17609, C2 =>
                           n12481, A => n15406, ZN => n15405);
   U15232 : OAI22_X1 port map( A1 => n16650, A2 => n17606, B1 => n16810, B2 => 
                           n17603, ZN => n15406);
   U15233 : AOI221_X1 port map( B1 => n17612, B2 => n12474, C1 => n17609, C2 =>
                           n12482, A => n15387, ZN => n15386);
   U15234 : OAI22_X1 port map( A1 => n16651, A2 => n17606, B1 => n16811, B2 => 
                           n17603, ZN => n15387);
   U15235 : AOI221_X1 port map( B1 => n17612, B2 => n12475, C1 => n17609, C2 =>
                           n12483, A => n15338, ZN => n15335);
   U15236 : OAI22_X1 port map( A1 => n16652, A2 => n17606, B1 => n16812, B2 => 
                           n17603, ZN => n15338);
   U15237 : AOI221_X1 port map( B1 => n17712, B2 => n12674, C1 => n17709, C2 =>
                           n12698, A => n15304, ZN => n15303);
   U15238 : OAI22_X1 port map( A1 => n16737, A2 => n17706, B1 => n17221, B2 => 
                           n17703, ZN => n15304);
   U15239 : AOI221_X1 port map( B1 => n17712, B2 => n12675, C1 => n17709, C2 =>
                           n12699, A => n15285, ZN => n15284);
   U15240 : OAI22_X1 port map( A1 => n16738, A2 => n17706, B1 => n17222, B2 => 
                           n17703, ZN => n15285);
   U15241 : AOI221_X1 port map( B1 => n17712, B2 => n12676, C1 => n17709, C2 =>
                           n12700, A => n15266, ZN => n15265);
   U15242 : OAI22_X1 port map( A1 => n16739, A2 => n17706, B1 => n17223, B2 => 
                           n17703, ZN => n15266);
   U15243 : AOI221_X1 port map( B1 => n17712, B2 => n12677, C1 => n17709, C2 =>
                           n12701, A => n15247, ZN => n15246);
   U15244 : OAI22_X1 port map( A1 => n16740, A2 => n17706, B1 => n17224, B2 => 
                           n17703, ZN => n15247);
   U15245 : AOI221_X1 port map( B1 => n17712, B2 => n12678, C1 => n17709, C2 =>
                           n12702, A => n15228, ZN => n15227);
   U15246 : OAI22_X1 port map( A1 => n16741, A2 => n17706, B1 => n17225, B2 => 
                           n17703, ZN => n15228);
   U15247 : AOI221_X1 port map( B1 => n17712, B2 => n12679, C1 => n17709, C2 =>
                           n12703, A => n15209, ZN => n15208);
   U15248 : OAI22_X1 port map( A1 => n16742, A2 => n17706, B1 => n17226, B2 => 
                           n17703, ZN => n15209);
   U15249 : AOI221_X1 port map( B1 => n17712, B2 => n12680, C1 => n17709, C2 =>
                           n12704, A => n15190, ZN => n15189);
   U15250 : OAI22_X1 port map( A1 => n16743, A2 => n17706, B1 => n17227, B2 => 
                           n17703, ZN => n15190);
   U15251 : AOI221_X1 port map( B1 => n17712, B2 => n12681, C1 => n17709, C2 =>
                           n12705, A => n15171, ZN => n15170);
   U15252 : OAI22_X1 port map( A1 => n16744, A2 => n17706, B1 => n17228, B2 => 
                           n17703, ZN => n15171);
   U15253 : AOI221_X1 port map( B1 => n17712, B2 => n12682, C1 => n17709, C2 =>
                           n12706, A => n15152, ZN => n15151);
   U15254 : OAI22_X1 port map( A1 => n16745, A2 => n17706, B1 => n17229, B2 => 
                           n17703, ZN => n15152);
   U15255 : AOI221_X1 port map( B1 => n17712, B2 => n12683, C1 => n17709, C2 =>
                           n12707, A => n15133, ZN => n15132);
   U15256 : OAI22_X1 port map( A1 => n16746, A2 => n17706, B1 => n17230, B2 => 
                           n17703, ZN => n15133);
   U15257 : AOI221_X1 port map( B1 => n17712, B2 => n12684, C1 => n17709, C2 =>
                           n12708, A => n15114, ZN => n15113);
   U15258 : OAI22_X1 port map( A1 => n16747, A2 => n17706, B1 => n17231, B2 => 
                           n17703, ZN => n15114);
   U15259 : AOI221_X1 port map( B1 => n17712, B2 => n12685, C1 => n17709, C2 =>
                           n12709, A => n15095, ZN => n15094);
   U15260 : OAI22_X1 port map( A1 => n16748, A2 => n17706, B1 => n17232, B2 => 
                           n17703, ZN => n15095);
   U15261 : AOI221_X1 port map( B1 => n17713, B2 => n12686, C1 => n17710, C2 =>
                           n12710, A => n15076, ZN => n15075);
   U15262 : OAI22_X1 port map( A1 => n16633, A2 => n17707, B1 => n17233, B2 => 
                           n17704, ZN => n15076);
   U15263 : AOI221_X1 port map( B1 => n17713, B2 => n12687, C1 => n17710, C2 =>
                           n12711, A => n15057, ZN => n15056);
   U15264 : OAI22_X1 port map( A1 => n16634, A2 => n17707, B1 => n17234, B2 => 
                           n17704, ZN => n15057);
   U15265 : AOI221_X1 port map( B1 => n17713, B2 => n12688, C1 => n17710, C2 =>
                           n12712, A => n15038, ZN => n15037);
   U15266 : OAI22_X1 port map( A1 => n16635, A2 => n17707, B1 => n17235, B2 => 
                           n17704, ZN => n15038);
   U15267 : AOI221_X1 port map( B1 => n17713, B2 => n12689, C1 => n17710, C2 =>
                           n12713, A => n15019, ZN => n15018);
   U15268 : OAI22_X1 port map( A1 => n16636, A2 => n17707, B1 => n17236, B2 => 
                           n17704, ZN => n15019);
   U15269 : AOI221_X1 port map( B1 => n17713, B2 => n12690, C1 => n17710, C2 =>
                           n12714, A => n15000, ZN => n14999);
   U15270 : OAI22_X1 port map( A1 => n16637, A2 => n17707, B1 => n17237, B2 => 
                           n17704, ZN => n15000);
   U15271 : AOI221_X1 port map( B1 => n17713, B2 => n12691, C1 => n17710, C2 =>
                           n12715, A => n14981, ZN => n14980);
   U15272 : OAI22_X1 port map( A1 => n16638, A2 => n17707, B1 => n17238, B2 => 
                           n17704, ZN => n14981);
   U15273 : AOI221_X1 port map( B1 => n17713, B2 => n12692, C1 => n17710, C2 =>
                           n12716, A => n14962, ZN => n14961);
   U15274 : OAI22_X1 port map( A1 => n16639, A2 => n17707, B1 => n17239, B2 => 
                           n17704, ZN => n14962);
   U15275 : AOI221_X1 port map( B1 => n17713, B2 => n12693, C1 => n17710, C2 =>
                           n12717, A => n14943, ZN => n14942);
   U15276 : OAI22_X1 port map( A1 => n16640, A2 => n17707, B1 => n17240, B2 => 
                           n17704, ZN => n14943);
   U15277 : AOI221_X1 port map( B1 => n17713, B2 => n12694, C1 => n17710, C2 =>
                           n12718, A => n14924, ZN => n14923);
   U15278 : OAI22_X1 port map( A1 => n16641, A2 => n17707, B1 => n17241, B2 => 
                           n17704, ZN => n14924);
   U15279 : AOI221_X1 port map( B1 => n17713, B2 => n12695, C1 => n17710, C2 =>
                           n12719, A => n14905, ZN => n14904);
   U15280 : OAI22_X1 port map( A1 => n16642, A2 => n17707, B1 => n17242, B2 => 
                           n17704, ZN => n14905);
   U15281 : AOI221_X1 port map( B1 => n17713, B2 => n12696, C1 => n17710, C2 =>
                           n12720, A => n14886, ZN => n14885);
   U15282 : OAI22_X1 port map( A1 => n16643, A2 => n17707, B1 => n17243, B2 => 
                           n17704, ZN => n14886);
   U15283 : AOI221_X1 port map( B1 => n17713, B2 => n12697, C1 => n17710, C2 =>
                           n12721, A => n14867, ZN => n14866);
   U15284 : OAI22_X1 port map( A1 => n16644, A2 => n17707, B1 => n17244, B2 => 
                           n17704, ZN => n14867);
   U15285 : AOI221_X1 port map( B1 => n17714, B2 => n12468, C1 => n17711, C2 =>
                           n12476, A => n14848, ZN => n14847);
   U15286 : OAI22_X1 port map( A1 => n16645, A2 => n17708, B1 => n16805, B2 => 
                           n17705, ZN => n14848);
   U15287 : AOI221_X1 port map( B1 => n17714, B2 => n12469, C1 => n17711, C2 =>
                           n12477, A => n14829, ZN => n14828);
   U15288 : OAI22_X1 port map( A1 => n16646, A2 => n17708, B1 => n16806, B2 => 
                           n17705, ZN => n14829);
   U15289 : AOI221_X1 port map( B1 => n17714, B2 => n12470, C1 => n17711, C2 =>
                           n12478, A => n14810, ZN => n14809);
   U15290 : OAI22_X1 port map( A1 => n16647, A2 => n17708, B1 => n16807, B2 => 
                           n17705, ZN => n14810);
   U15291 : AOI221_X1 port map( B1 => n17714, B2 => n12471, C1 => n17711, C2 =>
                           n12479, A => n14791, ZN => n14790);
   U15292 : OAI22_X1 port map( A1 => n16648, A2 => n17708, B1 => n16808, B2 => 
                           n17705, ZN => n14791);
   U15293 : AOI221_X1 port map( B1 => n17714, B2 => n12472, C1 => n17711, C2 =>
                           n12480, A => n14772, ZN => n14771);
   U15294 : OAI22_X1 port map( A1 => n16649, A2 => n17708, B1 => n16809, B2 => 
                           n17705, ZN => n14772);
   U15295 : AOI221_X1 port map( B1 => n17714, B2 => n12473, C1 => n17711, C2 =>
                           n12481, A => n14753, ZN => n14752);
   U15296 : OAI22_X1 port map( A1 => n16650, A2 => n17708, B1 => n16810, B2 => 
                           n17705, ZN => n14753);
   U15297 : AOI221_X1 port map( B1 => n17714, B2 => n12474, C1 => n17711, C2 =>
                           n12482, A => n14734, ZN => n14733);
   U15298 : OAI22_X1 port map( A1 => n16651, A2 => n17708, B1 => n16811, B2 => 
                           n17705, ZN => n14734);
   U15299 : AOI221_X1 port map( B1 => n17714, B2 => n12475, C1 => n17711, C2 =>
                           n12483, A => n14685, ZN => n14682);
   U15300 : OAI22_X1 port map( A1 => n16652, A2 => n17708, B1 => n16812, B2 => 
                           n17705, ZN => n14685);
   U15301 : OAI22_X1 port map( A1 => n17844, A2 => n18077, B1 => n14660, B2 => 
                           n17037, ZN => n3033);
   U15302 : OAI22_X1 port map( A1 => n17845, A2 => n18080, B1 => n14660, B2 => 
                           n17038, ZN => n3034);
   U15303 : OAI22_X1 port map( A1 => n17845, A2 => n18083, B1 => n14660, B2 => 
                           n17039, ZN => n3035);
   U15304 : OAI22_X1 port map( A1 => n17845, A2 => n18086, B1 => n14660, B2 => 
                           n17040, ZN => n3036);
   U15305 : OAI22_X1 port map( A1 => n17845, A2 => n18089, B1 => n14660, B2 => 
                           n17041, ZN => n3037);
   U15306 : OAI22_X1 port map( A1 => n17845, A2 => n18092, B1 => n14660, B2 => 
                           n17042, ZN => n3038);
   U15307 : OAI22_X1 port map( A1 => n17846, A2 => n18095, B1 => n14660, B2 => 
                           n17043, ZN => n3039);
   U15308 : OAI22_X1 port map( A1 => n17846, A2 => n18107, B1 => n14660, B2 => 
                           n17044, ZN => n3040);
   U15309 : OAI22_X1 port map( A1 => n17988, A2 => n18076, B1 => n9008, B2 => 
                           n14635, ZN => n3545);
   U15310 : OAI22_X1 port map( A1 => n17989, A2 => n18079, B1 => n8991, B2 => 
                           n14635, ZN => n3546);
   U15311 : OAI22_X1 port map( A1 => n17989, A2 => n18082, B1 => n8974, B2 => 
                           n14635, ZN => n3547);
   U15312 : OAI22_X1 port map( A1 => n17989, A2 => n18085, B1 => n8957, B2 => 
                           n14635, ZN => n3548);
   U15313 : OAI22_X1 port map( A1 => n17989, A2 => n18088, B1 => n8940, B2 => 
                           n14635, ZN => n3549);
   U15314 : OAI22_X1 port map( A1 => n17989, A2 => n18091, B1 => n8923, B2 => 
                           n14635, ZN => n3550);
   U15315 : OAI22_X1 port map( A1 => n17990, A2 => n18094, B1 => n8906, B2 => 
                           n14635, ZN => n3551);
   U15316 : OAI22_X1 port map( A1 => n17990, A2 => n18106, B1 => n8889, B2 => 
                           n14635, ZN => n3552);
   U15317 : OAI22_X1 port map( A1 => n17979, A2 => n18076, B1 => n9009, B2 => 
                           n14637, ZN => n3513);
   U15318 : OAI22_X1 port map( A1 => n17980, A2 => n18079, B1 => n8992, B2 => 
                           n14637, ZN => n3514);
   U15319 : OAI22_X1 port map( A1 => n17980, A2 => n18082, B1 => n8975, B2 => 
                           n14637, ZN => n3515);
   U15320 : OAI22_X1 port map( A1 => n17980, A2 => n18085, B1 => n8958, B2 => 
                           n14637, ZN => n3516);
   U15321 : OAI22_X1 port map( A1 => n17980, A2 => n18088, B1 => n8941, B2 => 
                           n14637, ZN => n3517);
   U15322 : OAI22_X1 port map( A1 => n17980, A2 => n18091, B1 => n8924, B2 => 
                           n14637, ZN => n3518);
   U15323 : OAI22_X1 port map( A1 => n17981, A2 => n18094, B1 => n8907, B2 => 
                           n14637, ZN => n3519);
   U15324 : OAI22_X1 port map( A1 => n17981, A2 => n18106, B1 => n8890, B2 => 
                           n14637, ZN => n3520);
   U15325 : OAI22_X1 port map( A1 => n17970, A2 => n18076, B1 => n6647, B2 => 
                           n14639, ZN => n3481);
   U15326 : OAI22_X1 port map( A1 => n17971, A2 => n18079, B1 => n6646, B2 => 
                           n14639, ZN => n3482);
   U15327 : OAI22_X1 port map( A1 => n17971, A2 => n18082, B1 => n6645, B2 => 
                           n14639, ZN => n3483);
   U15328 : OAI22_X1 port map( A1 => n17971, A2 => n18085, B1 => n6644, B2 => 
                           n14639, ZN => n3484);
   U15329 : OAI22_X1 port map( A1 => n17971, A2 => n18088, B1 => n6643, B2 => 
                           n14639, ZN => n3485);
   U15330 : OAI22_X1 port map( A1 => n17971, A2 => n18091, B1 => n6642, B2 => 
                           n14639, ZN => n3486);
   U15331 : OAI22_X1 port map( A1 => n17972, A2 => n18094, B1 => n6641, B2 => 
                           n14639, ZN => n3487);
   U15332 : OAI22_X1 port map( A1 => n17972, A2 => n18106, B1 => n6640, B2 => 
                           n14639, ZN => n3488);
   U15333 : OAI22_X1 port map( A1 => n17961, A2 => n18076, B1 => n6679, B2 => 
                           n14641, ZN => n3449);
   U15334 : OAI22_X1 port map( A1 => n17962, A2 => n18079, B1 => n6678, B2 => 
                           n14641, ZN => n3450);
   U15335 : OAI22_X1 port map( A1 => n17962, A2 => n18082, B1 => n6677, B2 => 
                           n14641, ZN => n3451);
   U15336 : OAI22_X1 port map( A1 => n17962, A2 => n18085, B1 => n6676, B2 => 
                           n14641, ZN => n3452);
   U15337 : OAI22_X1 port map( A1 => n17962, A2 => n18088, B1 => n6675, B2 => 
                           n14641, ZN => n3453);
   U15338 : OAI22_X1 port map( A1 => n17962, A2 => n18091, B1 => n6674, B2 => 
                           n14641, ZN => n3454);
   U15339 : OAI22_X1 port map( A1 => n17963, A2 => n18094, B1 => n6673, B2 => 
                           n14641, ZN => n3455);
   U15340 : OAI22_X1 port map( A1 => n17963, A2 => n18106, B1 => n6672, B2 => 
                           n14641, ZN => n3456);
   U15341 : OAI22_X1 port map( A1 => n17934, A2 => n18076, B1 => n9013, B2 => 
                           n14648, ZN => n3353);
   U15342 : OAI22_X1 port map( A1 => n17935, A2 => n18079, B1 => n8996, B2 => 
                           n14648, ZN => n3354);
   U15343 : OAI22_X1 port map( A1 => n17935, A2 => n18082, B1 => n8979, B2 => 
                           n14648, ZN => n3355);
   U15344 : OAI22_X1 port map( A1 => n17935, A2 => n18085, B1 => n8962, B2 => 
                           n14648, ZN => n3356);
   U15345 : OAI22_X1 port map( A1 => n17935, A2 => n18088, B1 => n8945, B2 => 
                           n14648, ZN => n3357);
   U15346 : OAI22_X1 port map( A1 => n17935, A2 => n18091, B1 => n8928, B2 => 
                           n14648, ZN => n3358);
   U15347 : OAI22_X1 port map( A1 => n17936, A2 => n18094, B1 => n8911, B2 => 
                           n14648, ZN => n3359);
   U15348 : OAI22_X1 port map( A1 => n17936, A2 => n18106, B1 => n8894, B2 => 
                           n14648, ZN => n3360);
   U15349 : OAI22_X1 port map( A1 => n17925, A2 => n18076, B1 => n9012, B2 => 
                           n14650, ZN => n3321);
   U15350 : OAI22_X1 port map( A1 => n17926, A2 => n18079, B1 => n8995, B2 => 
                           n14650, ZN => n3322);
   U15351 : OAI22_X1 port map( A1 => n17926, A2 => n18082, B1 => n8978, B2 => 
                           n14650, ZN => n3323);
   U15352 : OAI22_X1 port map( A1 => n17926, A2 => n18085, B1 => n8961, B2 => 
                           n14650, ZN => n3324);
   U15353 : OAI22_X1 port map( A1 => n17926, A2 => n18088, B1 => n8944, B2 => 
                           n14650, ZN => n3325);
   U15354 : OAI22_X1 port map( A1 => n17926, A2 => n18091, B1 => n8927, B2 => 
                           n14650, ZN => n3326);
   U15355 : OAI22_X1 port map( A1 => n17927, A2 => n18094, B1 => n8910, B2 => 
                           n14650, ZN => n3327);
   U15356 : OAI22_X1 port map( A1 => n17927, A2 => n18106, B1 => n8893, B2 => 
                           n14650, ZN => n3328);
   U15357 : OAI22_X1 port map( A1 => n17898, A2 => n18077, B1 => n9015, B2 => 
                           n14653, ZN => n3225);
   U15358 : OAI22_X1 port map( A1 => n17899, A2 => n18080, B1 => n8998, B2 => 
                           n14653, ZN => n3226);
   U15359 : OAI22_X1 port map( A1 => n17899, A2 => n18083, B1 => n8981, B2 => 
                           n14653, ZN => n3227);
   U15360 : OAI22_X1 port map( A1 => n17899, A2 => n18086, B1 => n8964, B2 => 
                           n14653, ZN => n3228);
   U15361 : OAI22_X1 port map( A1 => n17899, A2 => n18089, B1 => n8947, B2 => 
                           n14653, ZN => n3229);
   U15362 : OAI22_X1 port map( A1 => n17899, A2 => n18092, B1 => n8930, B2 => 
                           n14653, ZN => n3230);
   U15363 : OAI22_X1 port map( A1 => n17900, A2 => n18095, B1 => n8913, B2 => 
                           n14653, ZN => n3231);
   U15364 : OAI22_X1 port map( A1 => n17900, A2 => n18107, B1 => n8896, B2 => 
                           n14653, ZN => n3232);
   U15365 : OAI22_X1 port map( A1 => n17889, A2 => n18077, B1 => n9014, B2 => 
                           n14654, ZN => n3193);
   U15366 : OAI22_X1 port map( A1 => n17890, A2 => n18080, B1 => n8997, B2 => 
                           n14654, ZN => n3194);
   U15367 : OAI22_X1 port map( A1 => n17890, A2 => n18083, B1 => n8980, B2 => 
                           n14654, ZN => n3195);
   U15368 : OAI22_X1 port map( A1 => n17890, A2 => n18086, B1 => n8963, B2 => 
                           n14654, ZN => n3196);
   U15369 : OAI22_X1 port map( A1 => n17890, A2 => n18089, B1 => n8946, B2 => 
                           n14654, ZN => n3197);
   U15370 : OAI22_X1 port map( A1 => n17890, A2 => n18092, B1 => n8929, B2 => 
                           n14654, ZN => n3198);
   U15371 : OAI22_X1 port map( A1 => n17891, A2 => n18095, B1 => n8912, B2 => 
                           n14654, ZN => n3199);
   U15372 : OAI22_X1 port map( A1 => n17891, A2 => n18107, B1 => n8895, B2 => 
                           n14654, ZN => n3200);
   U15373 : OAI22_X1 port map( A1 => n17826, A2 => n18077, B1 => n9019, B2 => 
                           n14662, ZN => n2969);
   U15374 : OAI22_X1 port map( A1 => n17827, A2 => n18080, B1 => n9002, B2 => 
                           n14662, ZN => n2970);
   U15375 : OAI22_X1 port map( A1 => n17827, A2 => n18083, B1 => n8985, B2 => 
                           n14662, ZN => n2971);
   U15376 : OAI22_X1 port map( A1 => n17827, A2 => n18086, B1 => n8968, B2 => 
                           n14662, ZN => n2972);
   U15377 : OAI22_X1 port map( A1 => n17827, A2 => n18089, B1 => n8951, B2 => 
                           n14662, ZN => n2973);
   U15378 : OAI22_X1 port map( A1 => n17827, A2 => n18092, B1 => n8934, B2 => 
                           n14662, ZN => n2974);
   U15379 : OAI22_X1 port map( A1 => n17828, A2 => n18095, B1 => n8917, B2 => 
                           n14662, ZN => n2975);
   U15380 : OAI22_X1 port map( A1 => n17828, A2 => n18107, B1 => n8900, B2 => 
                           n14662, ZN => n2976);
   U15381 : OAI22_X1 port map( A1 => n17817, A2 => n18077, B1 => n9018, B2 => 
                           n14663, ZN => n2937);
   U15382 : OAI22_X1 port map( A1 => n17818, A2 => n18080, B1 => n9001, B2 => 
                           n14663, ZN => n2938);
   U15383 : OAI22_X1 port map( A1 => n17818, A2 => n18083, B1 => n8984, B2 => 
                           n14663, ZN => n2939);
   U15384 : OAI22_X1 port map( A1 => n17818, A2 => n18086, B1 => n8967, B2 => 
                           n14663, ZN => n2940);
   U15385 : OAI22_X1 port map( A1 => n17818, A2 => n18089, B1 => n8950, B2 => 
                           n14663, ZN => n2941);
   U15386 : OAI22_X1 port map( A1 => n17818, A2 => n18092, B1 => n8933, B2 => 
                           n14663, ZN => n2942);
   U15387 : OAI22_X1 port map( A1 => n17819, A2 => n18095, B1 => n8916, B2 => 
                           n14663, ZN => n2943);
   U15388 : OAI22_X1 port map( A1 => n17819, A2 => n18107, B1 => n8899, B2 => 
                           n14663, ZN => n2944);
   U15389 : OAI22_X1 port map( A1 => n17772, A2 => n18078, B1 => n9021, B2 => 
                           n14669, ZN => n2777);
   U15390 : OAI22_X1 port map( A1 => n17773, A2 => n18081, B1 => n9004, B2 => 
                           n14669, ZN => n2778);
   U15391 : OAI22_X1 port map( A1 => n17773, A2 => n18084, B1 => n8987, B2 => 
                           n14669, ZN => n2779);
   U15392 : OAI22_X1 port map( A1 => n17773, A2 => n18087, B1 => n8970, B2 => 
                           n14669, ZN => n2780);
   U15393 : OAI22_X1 port map( A1 => n17773, A2 => n18090, B1 => n8953, B2 => 
                           n14669, ZN => n2781);
   U15394 : OAI22_X1 port map( A1 => n17773, A2 => n18093, B1 => n8936, B2 => 
                           n14669, ZN => n2782);
   U15395 : OAI22_X1 port map( A1 => n17774, A2 => n18096, B1 => n8919, B2 => 
                           n14669, ZN => n2783);
   U15396 : OAI22_X1 port map( A1 => n17774, A2 => n18108, B1 => n8902, B2 => 
                           n14669, ZN => n2784);
   U15397 : OAI22_X1 port map( A1 => n17763, A2 => n18078, B1 => n9020, B2 => 
                           n14670, ZN => n2745);
   U15398 : OAI22_X1 port map( A1 => n17764, A2 => n18081, B1 => n9003, B2 => 
                           n14670, ZN => n2746);
   U15399 : OAI22_X1 port map( A1 => n17764, A2 => n18084, B1 => n8986, B2 => 
                           n14670, ZN => n2747);
   U15400 : OAI22_X1 port map( A1 => n17764, A2 => n18087, B1 => n8969, B2 => 
                           n14670, ZN => n2748);
   U15401 : OAI22_X1 port map( A1 => n17764, A2 => n18090, B1 => n8952, B2 => 
                           n14670, ZN => n2749);
   U15402 : OAI22_X1 port map( A1 => n17764, A2 => n18093, B1 => n8935, B2 => 
                           n14670, ZN => n2750);
   U15403 : OAI22_X1 port map( A1 => n17765, A2 => n18096, B1 => n8918, B2 => 
                           n14670, ZN => n2751);
   U15404 : OAI22_X1 port map( A1 => n17765, A2 => n18108, B1 => n8901, B2 => 
                           n14670, ZN => n2752);
   U15405 : OAI22_X1 port map( A1 => n17736, A2 => n18078, B1 => n9023, B2 => 
                           n14673, ZN => n2649);
   U15406 : OAI22_X1 port map( A1 => n17737, A2 => n18081, B1 => n9006, B2 => 
                           n14673, ZN => n2650);
   U15407 : OAI22_X1 port map( A1 => n17737, A2 => n18084, B1 => n8989, B2 => 
                           n14673, ZN => n2651);
   U15408 : OAI22_X1 port map( A1 => n17737, A2 => n18087, B1 => n8972, B2 => 
                           n14673, ZN => n2652);
   U15409 : OAI22_X1 port map( A1 => n17737, A2 => n18090, B1 => n8955, B2 => 
                           n14673, ZN => n2653);
   U15410 : OAI22_X1 port map( A1 => n17737, A2 => n18093, B1 => n8938, B2 => 
                           n14673, ZN => n2654);
   U15411 : OAI22_X1 port map( A1 => n17738, A2 => n18096, B1 => n8921, B2 => 
                           n14673, ZN => n2655);
   U15412 : OAI22_X1 port map( A1 => n17738, A2 => n18108, B1 => n8904, B2 => 
                           n14673, ZN => n2656);
   U15413 : OAI22_X1 port map( A1 => n17840, A2 => n18005, B1 => n17839, B2 => 
                           n17469, ZN => n3009);
   U15414 : OAI22_X1 port map( A1 => n17840, A2 => n18008, B1 => n17839, B2 => 
                           n17470, ZN => n3010);
   U15415 : OAI22_X1 port map( A1 => n17840, A2 => n18011, B1 => n17839, B2 => 
                           n17471, ZN => n3011);
   U15416 : OAI22_X1 port map( A1 => n17840, A2 => n18014, B1 => n17839, B2 => 
                           n17472, ZN => n3012);
   U15417 : OAI22_X1 port map( A1 => n17840, A2 => n18017, B1 => n17839, B2 => 
                           n17473, ZN => n3013);
   U15418 : OAI22_X1 port map( A1 => n17841, A2 => n18020, B1 => n17839, B2 => 
                           n17474, ZN => n3014);
   U15419 : OAI22_X1 port map( A1 => n17841, A2 => n18023, B1 => n17839, B2 => 
                           n17475, ZN => n3015);
   U15420 : OAI22_X1 port map( A1 => n17841, A2 => n18026, B1 => n17839, B2 => 
                           n17476, ZN => n3016);
   U15421 : OAI22_X1 port map( A1 => n17841, A2 => n18029, B1 => n17839, B2 => 
                           n17477, ZN => n3017);
   U15422 : OAI22_X1 port map( A1 => n17841, A2 => n18032, B1 => n17839, B2 => 
                           n17478, ZN => n3018);
   U15423 : OAI22_X1 port map( A1 => n17842, A2 => n18035, B1 => n17839, B2 => 
                           n17479, ZN => n3019);
   U15424 : OAI22_X1 port map( A1 => n17842, A2 => n18038, B1 => n17839, B2 => 
                           n17480, ZN => n3020);
   U15425 : OAI22_X1 port map( A1 => n17842, A2 => n18041, B1 => n14660, B2 => 
                           n17481, ZN => n3021);
   U15426 : OAI22_X1 port map( A1 => n17842, A2 => n18044, B1 => n14660, B2 => 
                           n17482, ZN => n3022);
   U15427 : OAI22_X1 port map( A1 => n17842, A2 => n18047, B1 => n14660, B2 => 
                           n17483, ZN => n3023);
   U15428 : OAI22_X1 port map( A1 => n17843, A2 => n18050, B1 => n17839, B2 => 
                           n17484, ZN => n3024);
   U15429 : OAI22_X1 port map( A1 => n17843, A2 => n18053, B1 => n17839, B2 => 
                           n17485, ZN => n3025);
   U15430 : OAI22_X1 port map( A1 => n17843, A2 => n18056, B1 => n17839, B2 => 
                           n17486, ZN => n3026);
   U15431 : OAI22_X1 port map( A1 => n17843, A2 => n18059, B1 => n17839, B2 => 
                           n17487, ZN => n3027);
   U15432 : OAI22_X1 port map( A1 => n17843, A2 => n18062, B1 => n17839, B2 => 
                           n17488, ZN => n3028);
   U15433 : OAI22_X1 port map( A1 => n17844, A2 => n18065, B1 => n17839, B2 => 
                           n17489, ZN => n3029);
   U15434 : OAI22_X1 port map( A1 => n17844, A2 => n18068, B1 => n17839, B2 => 
                           n17490, ZN => n3030);
   U15435 : OAI22_X1 port map( A1 => n17844, A2 => n18071, B1 => n17839, B2 => 
                           n17491, ZN => n3031);
   U15436 : OAI22_X1 port map( A1 => n17844, A2 => n18074, B1 => n17839, B2 => 
                           n17492, ZN => n3032);
   U15437 : OAI22_X1 port map( A1 => n9430, A2 => n14674, B1 => n17722, B2 => 
                           n18006, ZN => n2593);
   U15438 : OAI22_X1 port map( A1 => n9413, A2 => n17721, B1 => n17722, B2 => 
                           n18009, ZN => n2594);
   U15439 : OAI22_X1 port map( A1 => n9396, A2 => n17721, B1 => n17722, B2 => 
                           n18012, ZN => n2595);
   U15440 : OAI22_X1 port map( A1 => n9379, A2 => n17721, B1 => n17722, B2 => 
                           n18015, ZN => n2596);
   U15441 : OAI22_X1 port map( A1 => n9362, A2 => n17721, B1 => n17723, B2 => 
                           n18018, ZN => n2597);
   U15442 : OAI22_X1 port map( A1 => n9345, A2 => n17721, B1 => n17723, B2 => 
                           n18021, ZN => n2598);
   U15443 : OAI22_X1 port map( A1 => n9328, A2 => n17721, B1 => n17723, B2 => 
                           n18024, ZN => n2599);
   U15444 : OAI22_X1 port map( A1 => n9311, A2 => n17721, B1 => n17723, B2 => 
                           n18027, ZN => n2600);
   U15445 : OAI22_X1 port map( A1 => n9294, A2 => n17721, B1 => n17724, B2 => 
                           n18030, ZN => n2601);
   U15446 : OAI22_X1 port map( A1 => n9277, A2 => n17721, B1 => n17724, B2 => 
                           n18033, ZN => n2602);
   U15447 : OAI22_X1 port map( A1 => n9260, A2 => n17721, B1 => n17724, B2 => 
                           n18036, ZN => n2603);
   U15448 : OAI22_X1 port map( A1 => n9243, A2 => n17721, B1 => n17724, B2 => 
                           n18039, ZN => n2604);
   U15449 : OAI22_X1 port map( A1 => n9226, A2 => n14674, B1 => n17725, B2 => 
                           n18042, ZN => n2605);
   U15450 : OAI22_X1 port map( A1 => n9209, A2 => n17721, B1 => n17725, B2 => 
                           n18045, ZN => n2606);
   U15451 : OAI22_X1 port map( A1 => n9192, A2 => n14674, B1 => n17725, B2 => 
                           n18048, ZN => n2607);
   U15452 : OAI22_X1 port map( A1 => n9175, A2 => n17721, B1 => n17725, B2 => 
                           n18051, ZN => n2608);
   U15453 : OAI22_X1 port map( A1 => n9158, A2 => n14674, B1 => n17726, B2 => 
                           n18054, ZN => n2609);
   U15454 : OAI22_X1 port map( A1 => n9141, A2 => n17721, B1 => n17726, B2 => 
                           n18057, ZN => n2610);
   U15455 : OAI22_X1 port map( A1 => n9124, A2 => n14674, B1 => n17726, B2 => 
                           n18060, ZN => n2611);
   U15456 : OAI22_X1 port map( A1 => n9107, A2 => n17721, B1 => n17726, B2 => 
                           n18063, ZN => n2612);
   U15457 : OAI22_X1 port map( A1 => n9090, A2 => n14674, B1 => n17727, B2 => 
                           n18066, ZN => n2613);
   U15458 : OAI22_X1 port map( A1 => n9073, A2 => n17721, B1 => n17727, B2 => 
                           n18069, ZN => n2614);
   U15459 : OAI22_X1 port map( A1 => n9056, A2 => n14674, B1 => n17727, B2 => 
                           n18072, ZN => n2615);
   U15460 : OAI22_X1 port map( A1 => n9039, A2 => n17721, B1 => n17727, B2 => 
                           n18075, ZN => n2616);
   U15461 : OAI22_X1 port map( A1 => n9022, A2 => n14674, B1 => n17728, B2 => 
                           n18078, ZN => n2617);
   U15462 : OAI22_X1 port map( A1 => n9005, A2 => n17721, B1 => n17728, B2 => 
                           n18081, ZN => n2618);
   U15463 : OAI22_X1 port map( A1 => n8988, A2 => n14674, B1 => n17728, B2 => 
                           n18084, ZN => n2619);
   U15464 : OAI22_X1 port map( A1 => n8971, A2 => n17721, B1 => n17728, B2 => 
                           n18087, ZN => n2620);
   U15465 : OAI22_X1 port map( A1 => n8954, A2 => n14674, B1 => n17729, B2 => 
                           n18090, ZN => n2621);
   U15466 : OAI22_X1 port map( A1 => n8937, A2 => n17721, B1 => n17729, B2 => 
                           n18093, ZN => n2622);
   U15467 : OAI22_X1 port map( A1 => n8920, A2 => n14674, B1 => n17729, B2 => 
                           n18096, ZN => n2623);
   U15468 : OAI22_X1 port map( A1 => n8903, A2 => n17721, B1 => n17729, B2 => 
                           n18108, ZN => n2624);
   U15469 : OAI22_X1 port map( A1 => n17984, A2 => n18004, B1 => n9416, B2 => 
                           n17983, ZN => n3521);
   U15470 : OAI22_X1 port map( A1 => n17984, A2 => n18007, B1 => n9399, B2 => 
                           n17983, ZN => n3522);
   U15471 : OAI22_X1 port map( A1 => n17984, A2 => n18010, B1 => n9382, B2 => 
                           n17983, ZN => n3523);
   U15472 : OAI22_X1 port map( A1 => n17984, A2 => n18013, B1 => n9365, B2 => 
                           n17983, ZN => n3524);
   U15473 : OAI22_X1 port map( A1 => n17984, A2 => n18016, B1 => n9348, B2 => 
                           n17983, ZN => n3525);
   U15474 : OAI22_X1 port map( A1 => n17985, A2 => n18019, B1 => n9331, B2 => 
                           n17983, ZN => n3526);
   U15475 : OAI22_X1 port map( A1 => n17985, A2 => n18022, B1 => n9314, B2 => 
                           n17983, ZN => n3527);
   U15476 : OAI22_X1 port map( A1 => n17985, A2 => n18025, B1 => n9297, B2 => 
                           n17983, ZN => n3528);
   U15477 : OAI22_X1 port map( A1 => n17985, A2 => n18028, B1 => n9280, B2 => 
                           n17983, ZN => n3529);
   U15478 : OAI22_X1 port map( A1 => n17985, A2 => n18031, B1 => n9263, B2 => 
                           n17983, ZN => n3530);
   U15479 : OAI22_X1 port map( A1 => n17986, A2 => n18034, B1 => n9246, B2 => 
                           n17983, ZN => n3531);
   U15480 : OAI22_X1 port map( A1 => n17986, A2 => n18037, B1 => n9229, B2 => 
                           n17983, ZN => n3532);
   U15481 : OAI22_X1 port map( A1 => n17986, A2 => n18040, B1 => n9212, B2 => 
                           n14635, ZN => n3533);
   U15482 : OAI22_X1 port map( A1 => n17986, A2 => n18043, B1 => n9195, B2 => 
                           n14635, ZN => n3534);
   U15483 : OAI22_X1 port map( A1 => n17986, A2 => n18046, B1 => n9178, B2 => 
                           n14635, ZN => n3535);
   U15484 : OAI22_X1 port map( A1 => n17987, A2 => n18049, B1 => n9161, B2 => 
                           n17983, ZN => n3536);
   U15485 : OAI22_X1 port map( A1 => n17987, A2 => n18052, B1 => n9144, B2 => 
                           n17983, ZN => n3537);
   U15486 : OAI22_X1 port map( A1 => n17987, A2 => n18055, B1 => n9127, B2 => 
                           n17983, ZN => n3538);
   U15487 : OAI22_X1 port map( A1 => n17987, A2 => n18058, B1 => n9110, B2 => 
                           n17983, ZN => n3539);
   U15488 : OAI22_X1 port map( A1 => n17987, A2 => n18061, B1 => n9093, B2 => 
                           n17983, ZN => n3540);
   U15489 : OAI22_X1 port map( A1 => n17988, A2 => n18064, B1 => n9076, B2 => 
                           n17983, ZN => n3541);
   U15490 : OAI22_X1 port map( A1 => n17988, A2 => n18067, B1 => n9059, B2 => 
                           n17983, ZN => n3542);
   U15491 : OAI22_X1 port map( A1 => n17988, A2 => n18070, B1 => n9042, B2 => 
                           n17983, ZN => n3543);
   U15492 : OAI22_X1 port map( A1 => n17988, A2 => n18073, B1 => n9025, B2 => 
                           n17983, ZN => n3544);
   U15493 : OAI22_X1 port map( A1 => n17975, A2 => n18004, B1 => n9417, B2 => 
                           n17974, ZN => n3489);
   U15494 : OAI22_X1 port map( A1 => n17975, A2 => n18007, B1 => n9400, B2 => 
                           n17974, ZN => n3490);
   U15495 : OAI22_X1 port map( A1 => n17975, A2 => n18010, B1 => n9383, B2 => 
                           n17974, ZN => n3491);
   U15496 : OAI22_X1 port map( A1 => n17975, A2 => n18013, B1 => n9366, B2 => 
                           n17974, ZN => n3492);
   U15497 : OAI22_X1 port map( A1 => n17975, A2 => n18016, B1 => n9349, B2 => 
                           n17974, ZN => n3493);
   U15498 : OAI22_X1 port map( A1 => n17976, A2 => n18019, B1 => n9332, B2 => 
                           n17974, ZN => n3494);
   U15499 : OAI22_X1 port map( A1 => n17976, A2 => n18022, B1 => n9315, B2 => 
                           n17974, ZN => n3495);
   U15500 : OAI22_X1 port map( A1 => n17976, A2 => n18025, B1 => n9298, B2 => 
                           n17974, ZN => n3496);
   U15501 : OAI22_X1 port map( A1 => n17976, A2 => n18028, B1 => n9281, B2 => 
                           n17974, ZN => n3497);
   U15502 : OAI22_X1 port map( A1 => n17976, A2 => n18031, B1 => n9264, B2 => 
                           n17974, ZN => n3498);
   U15503 : OAI22_X1 port map( A1 => n17977, A2 => n18034, B1 => n9247, B2 => 
                           n17974, ZN => n3499);
   U15504 : OAI22_X1 port map( A1 => n17977, A2 => n18037, B1 => n9230, B2 => 
                           n17974, ZN => n3500);
   U15505 : OAI22_X1 port map( A1 => n17977, A2 => n18040, B1 => n9213, B2 => 
                           n14637, ZN => n3501);
   U15506 : OAI22_X1 port map( A1 => n17977, A2 => n18043, B1 => n9196, B2 => 
                           n14637, ZN => n3502);
   U15507 : OAI22_X1 port map( A1 => n17977, A2 => n18046, B1 => n9179, B2 => 
                           n14637, ZN => n3503);
   U15508 : OAI22_X1 port map( A1 => n17978, A2 => n18049, B1 => n9162, B2 => 
                           n17974, ZN => n3504);
   U15509 : OAI22_X1 port map( A1 => n17978, A2 => n18052, B1 => n9145, B2 => 
                           n17974, ZN => n3505);
   U15510 : OAI22_X1 port map( A1 => n17978, A2 => n18055, B1 => n9128, B2 => 
                           n17974, ZN => n3506);
   U15511 : OAI22_X1 port map( A1 => n17978, A2 => n18058, B1 => n9111, B2 => 
                           n17974, ZN => n3507);
   U15512 : OAI22_X1 port map( A1 => n17978, A2 => n18061, B1 => n9094, B2 => 
                           n17974, ZN => n3508);
   U15513 : OAI22_X1 port map( A1 => n17979, A2 => n18064, B1 => n9077, B2 => 
                           n17974, ZN => n3509);
   U15514 : OAI22_X1 port map( A1 => n17979, A2 => n18067, B1 => n9060, B2 => 
                           n17974, ZN => n3510);
   U15515 : OAI22_X1 port map( A1 => n17979, A2 => n18070, B1 => n9043, B2 => 
                           n17974, ZN => n3511);
   U15516 : OAI22_X1 port map( A1 => n17979, A2 => n18073, B1 => n9026, B2 => 
                           n17974, ZN => n3512);
   U15517 : OAI22_X1 port map( A1 => n17966, A2 => n18004, B1 => n6671, B2 => 
                           n17965, ZN => n3457);
   U15518 : OAI22_X1 port map( A1 => n17966, A2 => n18007, B1 => n6670, B2 => 
                           n17965, ZN => n3458);
   U15519 : OAI22_X1 port map( A1 => n17966, A2 => n18010, B1 => n6669, B2 => 
                           n17965, ZN => n3459);
   U15520 : OAI22_X1 port map( A1 => n17966, A2 => n18013, B1 => n6668, B2 => 
                           n17965, ZN => n3460);
   U15521 : OAI22_X1 port map( A1 => n17966, A2 => n18016, B1 => n6667, B2 => 
                           n17965, ZN => n3461);
   U15522 : OAI22_X1 port map( A1 => n17967, A2 => n18019, B1 => n6666, B2 => 
                           n17965, ZN => n3462);
   U15523 : OAI22_X1 port map( A1 => n17967, A2 => n18022, B1 => n6665, B2 => 
                           n17965, ZN => n3463);
   U15524 : OAI22_X1 port map( A1 => n17967, A2 => n18025, B1 => n6664, B2 => 
                           n17965, ZN => n3464);
   U15525 : OAI22_X1 port map( A1 => n17967, A2 => n18028, B1 => n6663, B2 => 
                           n17965, ZN => n3465);
   U15526 : OAI22_X1 port map( A1 => n17967, A2 => n18031, B1 => n6662, B2 => 
                           n17965, ZN => n3466);
   U15527 : OAI22_X1 port map( A1 => n17968, A2 => n18034, B1 => n6661, B2 => 
                           n17965, ZN => n3467);
   U15528 : OAI22_X1 port map( A1 => n17968, A2 => n18037, B1 => n6660, B2 => 
                           n17965, ZN => n3468);
   U15529 : OAI22_X1 port map( A1 => n17968, A2 => n18040, B1 => n6659, B2 => 
                           n14639, ZN => n3469);
   U15530 : OAI22_X1 port map( A1 => n17968, A2 => n18043, B1 => n6658, B2 => 
                           n14639, ZN => n3470);
   U15531 : OAI22_X1 port map( A1 => n17968, A2 => n18046, B1 => n6657, B2 => 
                           n14639, ZN => n3471);
   U15532 : OAI22_X1 port map( A1 => n17969, A2 => n18049, B1 => n6656, B2 => 
                           n17965, ZN => n3472);
   U15533 : OAI22_X1 port map( A1 => n17969, A2 => n18052, B1 => n6655, B2 => 
                           n17965, ZN => n3473);
   U15534 : OAI22_X1 port map( A1 => n17969, A2 => n18055, B1 => n6654, B2 => 
                           n17965, ZN => n3474);
   U15535 : OAI22_X1 port map( A1 => n17969, A2 => n18058, B1 => n6653, B2 => 
                           n17965, ZN => n3475);
   U15536 : OAI22_X1 port map( A1 => n17969, A2 => n18061, B1 => n6652, B2 => 
                           n17965, ZN => n3476);
   U15537 : OAI22_X1 port map( A1 => n17970, A2 => n18064, B1 => n6651, B2 => 
                           n17965, ZN => n3477);
   U15538 : OAI22_X1 port map( A1 => n17970, A2 => n18067, B1 => n6650, B2 => 
                           n17965, ZN => n3478);
   U15539 : OAI22_X1 port map( A1 => n17970, A2 => n18070, B1 => n6649, B2 => 
                           n17965, ZN => n3479);
   U15540 : OAI22_X1 port map( A1 => n17970, A2 => n18073, B1 => n6648, B2 => 
                           n17965, ZN => n3480);
   U15541 : OAI22_X1 port map( A1 => n17957, A2 => n18004, B1 => n6703, B2 => 
                           n17956, ZN => n3425);
   U15542 : OAI22_X1 port map( A1 => n17957, A2 => n18007, B1 => n6702, B2 => 
                           n17956, ZN => n3426);
   U15543 : OAI22_X1 port map( A1 => n17957, A2 => n18010, B1 => n6701, B2 => 
                           n17956, ZN => n3427);
   U15544 : OAI22_X1 port map( A1 => n17957, A2 => n18013, B1 => n6700, B2 => 
                           n17956, ZN => n3428);
   U15545 : OAI22_X1 port map( A1 => n17957, A2 => n18016, B1 => n6699, B2 => 
                           n17956, ZN => n3429);
   U15546 : OAI22_X1 port map( A1 => n17958, A2 => n18019, B1 => n6698, B2 => 
                           n17956, ZN => n3430);
   U15547 : OAI22_X1 port map( A1 => n17958, A2 => n18022, B1 => n6697, B2 => 
                           n17956, ZN => n3431);
   U15548 : OAI22_X1 port map( A1 => n17958, A2 => n18025, B1 => n6696, B2 => 
                           n17956, ZN => n3432);
   U15549 : OAI22_X1 port map( A1 => n17958, A2 => n18028, B1 => n6695, B2 => 
                           n17956, ZN => n3433);
   U15550 : OAI22_X1 port map( A1 => n17958, A2 => n18031, B1 => n6694, B2 => 
                           n17956, ZN => n3434);
   U15551 : OAI22_X1 port map( A1 => n17959, A2 => n18034, B1 => n6693, B2 => 
                           n17956, ZN => n3435);
   U15552 : OAI22_X1 port map( A1 => n17959, A2 => n18037, B1 => n6692, B2 => 
                           n17956, ZN => n3436);
   U15553 : OAI22_X1 port map( A1 => n17959, A2 => n18040, B1 => n6691, B2 => 
                           n14641, ZN => n3437);
   U15554 : OAI22_X1 port map( A1 => n17959, A2 => n18043, B1 => n6690, B2 => 
                           n14641, ZN => n3438);
   U15555 : OAI22_X1 port map( A1 => n17959, A2 => n18046, B1 => n6689, B2 => 
                           n14641, ZN => n3439);
   U15556 : OAI22_X1 port map( A1 => n17960, A2 => n18049, B1 => n6688, B2 => 
                           n17956, ZN => n3440);
   U15557 : OAI22_X1 port map( A1 => n17960, A2 => n18052, B1 => n6687, B2 => 
                           n17956, ZN => n3441);
   U15558 : OAI22_X1 port map( A1 => n17960, A2 => n18055, B1 => n6686, B2 => 
                           n17956, ZN => n3442);
   U15559 : OAI22_X1 port map( A1 => n17960, A2 => n18058, B1 => n6685, B2 => 
                           n17956, ZN => n3443);
   U15560 : OAI22_X1 port map( A1 => n17960, A2 => n18061, B1 => n6684, B2 => 
                           n17956, ZN => n3444);
   U15561 : OAI22_X1 port map( A1 => n17961, A2 => n18064, B1 => n6683, B2 => 
                           n17956, ZN => n3445);
   U15562 : OAI22_X1 port map( A1 => n17961, A2 => n18067, B1 => n6682, B2 => 
                           n17956, ZN => n3446);
   U15563 : OAI22_X1 port map( A1 => n17961, A2 => n18070, B1 => n6681, B2 => 
                           n17956, ZN => n3447);
   U15564 : OAI22_X1 port map( A1 => n17961, A2 => n18073, B1 => n6680, B2 => 
                           n17956, ZN => n3448);
   U15565 : OAI22_X1 port map( A1 => n17930, A2 => n18004, B1 => n9421, B2 => 
                           n17929, ZN => n3329);
   U15566 : OAI22_X1 port map( A1 => n17930, A2 => n18007, B1 => n9404, B2 => 
                           n17929, ZN => n3330);
   U15567 : OAI22_X1 port map( A1 => n17930, A2 => n18010, B1 => n9387, B2 => 
                           n17929, ZN => n3331);
   U15568 : OAI22_X1 port map( A1 => n17930, A2 => n18013, B1 => n9370, B2 => 
                           n17929, ZN => n3332);
   U15569 : OAI22_X1 port map( A1 => n17930, A2 => n18016, B1 => n9353, B2 => 
                           n17929, ZN => n3333);
   U15570 : OAI22_X1 port map( A1 => n17931, A2 => n18019, B1 => n9336, B2 => 
                           n17929, ZN => n3334);
   U15571 : OAI22_X1 port map( A1 => n17931, A2 => n18022, B1 => n9319, B2 => 
                           n17929, ZN => n3335);
   U15572 : OAI22_X1 port map( A1 => n17931, A2 => n18025, B1 => n9302, B2 => 
                           n17929, ZN => n3336);
   U15573 : OAI22_X1 port map( A1 => n17931, A2 => n18028, B1 => n9285, B2 => 
                           n17929, ZN => n3337);
   U15574 : OAI22_X1 port map( A1 => n17931, A2 => n18031, B1 => n9268, B2 => 
                           n17929, ZN => n3338);
   U15575 : OAI22_X1 port map( A1 => n17932, A2 => n18034, B1 => n9251, B2 => 
                           n17929, ZN => n3339);
   U15576 : OAI22_X1 port map( A1 => n17932, A2 => n18037, B1 => n9234, B2 => 
                           n17929, ZN => n3340);
   U15577 : OAI22_X1 port map( A1 => n17932, A2 => n18040, B1 => n9217, B2 => 
                           n14648, ZN => n3341);
   U15578 : OAI22_X1 port map( A1 => n17932, A2 => n18043, B1 => n9200, B2 => 
                           n14648, ZN => n3342);
   U15579 : OAI22_X1 port map( A1 => n17932, A2 => n18046, B1 => n9183, B2 => 
                           n14648, ZN => n3343);
   U15580 : OAI22_X1 port map( A1 => n17933, A2 => n18049, B1 => n9166, B2 => 
                           n17929, ZN => n3344);
   U15581 : OAI22_X1 port map( A1 => n17933, A2 => n18052, B1 => n9149, B2 => 
                           n17929, ZN => n3345);
   U15582 : OAI22_X1 port map( A1 => n17933, A2 => n18055, B1 => n9132, B2 => 
                           n17929, ZN => n3346);
   U15583 : OAI22_X1 port map( A1 => n17933, A2 => n18058, B1 => n9115, B2 => 
                           n17929, ZN => n3347);
   U15584 : OAI22_X1 port map( A1 => n17933, A2 => n18061, B1 => n9098, B2 => 
                           n17929, ZN => n3348);
   U15585 : OAI22_X1 port map( A1 => n17934, A2 => n18064, B1 => n9081, B2 => 
                           n17929, ZN => n3349);
   U15586 : OAI22_X1 port map( A1 => n17934, A2 => n18067, B1 => n9064, B2 => 
                           n17929, ZN => n3350);
   U15587 : OAI22_X1 port map( A1 => n17934, A2 => n18070, B1 => n9047, B2 => 
                           n17929, ZN => n3351);
   U15588 : OAI22_X1 port map( A1 => n17934, A2 => n18073, B1 => n9030, B2 => 
                           n17929, ZN => n3352);
   U15589 : OAI22_X1 port map( A1 => n17921, A2 => n18004, B1 => n9420, B2 => 
                           n17920, ZN => n3297);
   U15590 : OAI22_X1 port map( A1 => n17921, A2 => n18007, B1 => n9403, B2 => 
                           n17920, ZN => n3298);
   U15591 : OAI22_X1 port map( A1 => n17921, A2 => n18010, B1 => n9386, B2 => 
                           n17920, ZN => n3299);
   U15592 : OAI22_X1 port map( A1 => n17921, A2 => n18013, B1 => n9369, B2 => 
                           n17920, ZN => n3300);
   U15593 : OAI22_X1 port map( A1 => n17921, A2 => n18016, B1 => n9352, B2 => 
                           n17920, ZN => n3301);
   U15594 : OAI22_X1 port map( A1 => n17922, A2 => n18019, B1 => n9335, B2 => 
                           n17920, ZN => n3302);
   U15595 : OAI22_X1 port map( A1 => n17922, A2 => n18022, B1 => n9318, B2 => 
                           n17920, ZN => n3303);
   U15596 : OAI22_X1 port map( A1 => n17922, A2 => n18025, B1 => n9301, B2 => 
                           n17920, ZN => n3304);
   U15597 : OAI22_X1 port map( A1 => n17922, A2 => n18028, B1 => n9284, B2 => 
                           n17920, ZN => n3305);
   U15598 : OAI22_X1 port map( A1 => n17922, A2 => n18031, B1 => n9267, B2 => 
                           n17920, ZN => n3306);
   U15599 : OAI22_X1 port map( A1 => n17923, A2 => n18034, B1 => n9250, B2 => 
                           n17920, ZN => n3307);
   U15600 : OAI22_X1 port map( A1 => n17923, A2 => n18037, B1 => n9233, B2 => 
                           n17920, ZN => n3308);
   U15601 : OAI22_X1 port map( A1 => n17923, A2 => n18040, B1 => n9216, B2 => 
                           n14650, ZN => n3309);
   U15602 : OAI22_X1 port map( A1 => n17923, A2 => n18043, B1 => n9199, B2 => 
                           n14650, ZN => n3310);
   U15603 : OAI22_X1 port map( A1 => n17923, A2 => n18046, B1 => n9182, B2 => 
                           n14650, ZN => n3311);
   U15604 : OAI22_X1 port map( A1 => n17924, A2 => n18049, B1 => n9165, B2 => 
                           n17920, ZN => n3312);
   U15605 : OAI22_X1 port map( A1 => n17924, A2 => n18052, B1 => n9148, B2 => 
                           n17920, ZN => n3313);
   U15606 : OAI22_X1 port map( A1 => n17924, A2 => n18055, B1 => n9131, B2 => 
                           n17920, ZN => n3314);
   U15607 : OAI22_X1 port map( A1 => n17924, A2 => n18058, B1 => n9114, B2 => 
                           n17920, ZN => n3315);
   U15608 : OAI22_X1 port map( A1 => n17924, A2 => n18061, B1 => n9097, B2 => 
                           n17920, ZN => n3316);
   U15609 : OAI22_X1 port map( A1 => n17925, A2 => n18064, B1 => n9080, B2 => 
                           n17920, ZN => n3317);
   U15610 : OAI22_X1 port map( A1 => n17925, A2 => n18067, B1 => n9063, B2 => 
                           n17920, ZN => n3318);
   U15611 : OAI22_X1 port map( A1 => n17925, A2 => n18070, B1 => n9046, B2 => 
                           n17920, ZN => n3319);
   U15612 : OAI22_X1 port map( A1 => n17925, A2 => n18073, B1 => n9029, B2 => 
                           n17920, ZN => n3320);
   U15613 : OAI22_X1 port map( A1 => n17894, A2 => n18005, B1 => n9423, B2 => 
                           n17893, ZN => n3201);
   U15614 : OAI22_X1 port map( A1 => n17894, A2 => n18008, B1 => n9406, B2 => 
                           n17893, ZN => n3202);
   U15615 : OAI22_X1 port map( A1 => n17894, A2 => n18011, B1 => n9389, B2 => 
                           n17893, ZN => n3203);
   U15616 : OAI22_X1 port map( A1 => n17894, A2 => n18014, B1 => n9372, B2 => 
                           n17893, ZN => n3204);
   U15617 : OAI22_X1 port map( A1 => n17894, A2 => n18017, B1 => n9355, B2 => 
                           n17893, ZN => n3205);
   U15618 : OAI22_X1 port map( A1 => n17895, A2 => n18020, B1 => n9338, B2 => 
                           n17893, ZN => n3206);
   U15619 : OAI22_X1 port map( A1 => n17895, A2 => n18023, B1 => n9321, B2 => 
                           n17893, ZN => n3207);
   U15620 : OAI22_X1 port map( A1 => n17895, A2 => n18026, B1 => n9304, B2 => 
                           n17893, ZN => n3208);
   U15621 : OAI22_X1 port map( A1 => n17895, A2 => n18029, B1 => n9287, B2 => 
                           n17893, ZN => n3209);
   U15622 : OAI22_X1 port map( A1 => n17895, A2 => n18032, B1 => n9270, B2 => 
                           n17893, ZN => n3210);
   U15623 : OAI22_X1 port map( A1 => n17896, A2 => n18035, B1 => n9253, B2 => 
                           n17893, ZN => n3211);
   U15624 : OAI22_X1 port map( A1 => n17896, A2 => n18038, B1 => n9236, B2 => 
                           n17893, ZN => n3212);
   U15625 : OAI22_X1 port map( A1 => n17896, A2 => n18041, B1 => n9219, B2 => 
                           n14653, ZN => n3213);
   U15626 : OAI22_X1 port map( A1 => n17896, A2 => n18044, B1 => n9202, B2 => 
                           n14653, ZN => n3214);
   U15627 : OAI22_X1 port map( A1 => n17896, A2 => n18047, B1 => n9185, B2 => 
                           n14653, ZN => n3215);
   U15628 : OAI22_X1 port map( A1 => n17897, A2 => n18050, B1 => n9168, B2 => 
                           n17893, ZN => n3216);
   U15629 : OAI22_X1 port map( A1 => n17897, A2 => n18053, B1 => n9151, B2 => 
                           n17893, ZN => n3217);
   U15630 : OAI22_X1 port map( A1 => n17897, A2 => n18056, B1 => n9134, B2 => 
                           n17893, ZN => n3218);
   U15631 : OAI22_X1 port map( A1 => n17897, A2 => n18059, B1 => n9117, B2 => 
                           n17893, ZN => n3219);
   U15632 : OAI22_X1 port map( A1 => n17897, A2 => n18062, B1 => n9100, B2 => 
                           n17893, ZN => n3220);
   U15633 : OAI22_X1 port map( A1 => n17898, A2 => n18065, B1 => n9083, B2 => 
                           n17893, ZN => n3221);
   U15634 : OAI22_X1 port map( A1 => n17898, A2 => n18068, B1 => n9066, B2 => 
                           n17893, ZN => n3222);
   U15635 : OAI22_X1 port map( A1 => n17898, A2 => n18071, B1 => n9049, B2 => 
                           n17893, ZN => n3223);
   U15636 : OAI22_X1 port map( A1 => n17898, A2 => n18074, B1 => n9032, B2 => 
                           n17893, ZN => n3224);
   U15637 : OAI22_X1 port map( A1 => n17885, A2 => n18005, B1 => n9422, B2 => 
                           n17884, ZN => n3169);
   U15638 : OAI22_X1 port map( A1 => n17885, A2 => n18008, B1 => n9405, B2 => 
                           n17884, ZN => n3170);
   U15639 : OAI22_X1 port map( A1 => n17885, A2 => n18011, B1 => n9388, B2 => 
                           n17884, ZN => n3171);
   U15640 : OAI22_X1 port map( A1 => n17885, A2 => n18014, B1 => n9371, B2 => 
                           n17884, ZN => n3172);
   U15641 : OAI22_X1 port map( A1 => n17885, A2 => n18017, B1 => n9354, B2 => 
                           n17884, ZN => n3173);
   U15642 : OAI22_X1 port map( A1 => n17886, A2 => n18020, B1 => n9337, B2 => 
                           n17884, ZN => n3174);
   U15643 : OAI22_X1 port map( A1 => n17886, A2 => n18023, B1 => n9320, B2 => 
                           n17884, ZN => n3175);
   U15644 : OAI22_X1 port map( A1 => n17886, A2 => n18026, B1 => n9303, B2 => 
                           n17884, ZN => n3176);
   U15645 : OAI22_X1 port map( A1 => n17886, A2 => n18029, B1 => n9286, B2 => 
                           n17884, ZN => n3177);
   U15646 : OAI22_X1 port map( A1 => n17886, A2 => n18032, B1 => n9269, B2 => 
                           n17884, ZN => n3178);
   U15647 : OAI22_X1 port map( A1 => n17887, A2 => n18035, B1 => n9252, B2 => 
                           n17884, ZN => n3179);
   U15648 : OAI22_X1 port map( A1 => n17887, A2 => n18038, B1 => n9235, B2 => 
                           n17884, ZN => n3180);
   U15649 : OAI22_X1 port map( A1 => n17887, A2 => n18041, B1 => n9218, B2 => 
                           n14654, ZN => n3181);
   U15650 : OAI22_X1 port map( A1 => n17887, A2 => n18044, B1 => n9201, B2 => 
                           n14654, ZN => n3182);
   U15651 : OAI22_X1 port map( A1 => n17887, A2 => n18047, B1 => n9184, B2 => 
                           n14654, ZN => n3183);
   U15652 : OAI22_X1 port map( A1 => n17888, A2 => n18050, B1 => n9167, B2 => 
                           n17884, ZN => n3184);
   U15653 : OAI22_X1 port map( A1 => n17888, A2 => n18053, B1 => n9150, B2 => 
                           n17884, ZN => n3185);
   U15654 : OAI22_X1 port map( A1 => n17888, A2 => n18056, B1 => n9133, B2 => 
                           n17884, ZN => n3186);
   U15655 : OAI22_X1 port map( A1 => n17888, A2 => n18059, B1 => n9116, B2 => 
                           n17884, ZN => n3187);
   U15656 : OAI22_X1 port map( A1 => n17888, A2 => n18062, B1 => n9099, B2 => 
                           n17884, ZN => n3188);
   U15657 : OAI22_X1 port map( A1 => n17889, A2 => n18065, B1 => n9082, B2 => 
                           n17884, ZN => n3189);
   U15658 : OAI22_X1 port map( A1 => n17889, A2 => n18068, B1 => n9065, B2 => 
                           n17884, ZN => n3190);
   U15659 : OAI22_X1 port map( A1 => n17889, A2 => n18071, B1 => n9048, B2 => 
                           n17884, ZN => n3191);
   U15660 : OAI22_X1 port map( A1 => n17889, A2 => n18074, B1 => n9031, B2 => 
                           n17884, ZN => n3192);
   U15661 : OAI22_X1 port map( A1 => n17822, A2 => n18005, B1 => n9427, B2 => 
                           n17821, ZN => n2945);
   U15662 : OAI22_X1 port map( A1 => n17822, A2 => n18008, B1 => n9410, B2 => 
                           n17821, ZN => n2946);
   U15663 : OAI22_X1 port map( A1 => n17822, A2 => n18011, B1 => n9393, B2 => 
                           n17821, ZN => n2947);
   U15664 : OAI22_X1 port map( A1 => n17822, A2 => n18014, B1 => n9376, B2 => 
                           n17821, ZN => n2948);
   U15665 : OAI22_X1 port map( A1 => n17822, A2 => n18017, B1 => n9359, B2 => 
                           n17821, ZN => n2949);
   U15666 : OAI22_X1 port map( A1 => n17823, A2 => n18020, B1 => n9342, B2 => 
                           n17821, ZN => n2950);
   U15667 : OAI22_X1 port map( A1 => n17823, A2 => n18023, B1 => n9325, B2 => 
                           n17821, ZN => n2951);
   U15668 : OAI22_X1 port map( A1 => n17823, A2 => n18026, B1 => n9308, B2 => 
                           n17821, ZN => n2952);
   U15669 : OAI22_X1 port map( A1 => n17823, A2 => n18029, B1 => n9291, B2 => 
                           n17821, ZN => n2953);
   U15670 : OAI22_X1 port map( A1 => n17823, A2 => n18032, B1 => n9274, B2 => 
                           n17821, ZN => n2954);
   U15671 : OAI22_X1 port map( A1 => n17824, A2 => n18035, B1 => n9257, B2 => 
                           n17821, ZN => n2955);
   U15672 : OAI22_X1 port map( A1 => n17824, A2 => n18038, B1 => n9240, B2 => 
                           n17821, ZN => n2956);
   U15673 : OAI22_X1 port map( A1 => n17824, A2 => n18041, B1 => n9223, B2 => 
                           n14662, ZN => n2957);
   U15674 : OAI22_X1 port map( A1 => n17824, A2 => n18044, B1 => n9206, B2 => 
                           n14662, ZN => n2958);
   U15675 : OAI22_X1 port map( A1 => n17824, A2 => n18047, B1 => n9189, B2 => 
                           n14662, ZN => n2959);
   U15676 : OAI22_X1 port map( A1 => n17825, A2 => n18050, B1 => n9172, B2 => 
                           n17821, ZN => n2960);
   U15677 : OAI22_X1 port map( A1 => n17825, A2 => n18053, B1 => n9155, B2 => 
                           n17821, ZN => n2961);
   U15678 : OAI22_X1 port map( A1 => n17825, A2 => n18056, B1 => n9138, B2 => 
                           n17821, ZN => n2962);
   U15679 : OAI22_X1 port map( A1 => n17825, A2 => n18059, B1 => n9121, B2 => 
                           n17821, ZN => n2963);
   U15680 : OAI22_X1 port map( A1 => n17825, A2 => n18062, B1 => n9104, B2 => 
                           n17821, ZN => n2964);
   U15681 : OAI22_X1 port map( A1 => n17826, A2 => n18065, B1 => n9087, B2 => 
                           n17821, ZN => n2965);
   U15682 : OAI22_X1 port map( A1 => n17826, A2 => n18068, B1 => n9070, B2 => 
                           n17821, ZN => n2966);
   U15683 : OAI22_X1 port map( A1 => n17826, A2 => n18071, B1 => n9053, B2 => 
                           n17821, ZN => n2967);
   U15684 : OAI22_X1 port map( A1 => n17826, A2 => n18074, B1 => n9036, B2 => 
                           n17821, ZN => n2968);
   U15685 : OAI22_X1 port map( A1 => n17813, A2 => n18005, B1 => n9426, B2 => 
                           n17812, ZN => n2913);
   U15686 : OAI22_X1 port map( A1 => n17813, A2 => n18008, B1 => n9409, B2 => 
                           n17812, ZN => n2914);
   U15687 : OAI22_X1 port map( A1 => n17813, A2 => n18011, B1 => n9392, B2 => 
                           n17812, ZN => n2915);
   U15688 : OAI22_X1 port map( A1 => n17813, A2 => n18014, B1 => n9375, B2 => 
                           n17812, ZN => n2916);
   U15689 : OAI22_X1 port map( A1 => n17813, A2 => n18017, B1 => n9358, B2 => 
                           n17812, ZN => n2917);
   U15690 : OAI22_X1 port map( A1 => n17814, A2 => n18020, B1 => n9341, B2 => 
                           n17812, ZN => n2918);
   U15691 : OAI22_X1 port map( A1 => n17814, A2 => n18023, B1 => n9324, B2 => 
                           n17812, ZN => n2919);
   U15692 : OAI22_X1 port map( A1 => n17814, A2 => n18026, B1 => n9307, B2 => 
                           n17812, ZN => n2920);
   U15693 : OAI22_X1 port map( A1 => n17814, A2 => n18029, B1 => n9290, B2 => 
                           n17812, ZN => n2921);
   U15694 : OAI22_X1 port map( A1 => n17814, A2 => n18032, B1 => n9273, B2 => 
                           n17812, ZN => n2922);
   U15695 : OAI22_X1 port map( A1 => n17815, A2 => n18035, B1 => n9256, B2 => 
                           n17812, ZN => n2923);
   U15696 : OAI22_X1 port map( A1 => n17815, A2 => n18038, B1 => n9239, B2 => 
                           n17812, ZN => n2924);
   U15697 : OAI22_X1 port map( A1 => n17815, A2 => n18041, B1 => n9222, B2 => 
                           n14663, ZN => n2925);
   U15698 : OAI22_X1 port map( A1 => n17815, A2 => n18044, B1 => n9205, B2 => 
                           n14663, ZN => n2926);
   U15699 : OAI22_X1 port map( A1 => n17815, A2 => n18047, B1 => n9188, B2 => 
                           n14663, ZN => n2927);
   U15700 : OAI22_X1 port map( A1 => n17816, A2 => n18050, B1 => n9171, B2 => 
                           n17812, ZN => n2928);
   U15701 : OAI22_X1 port map( A1 => n17816, A2 => n18053, B1 => n9154, B2 => 
                           n17812, ZN => n2929);
   U15702 : OAI22_X1 port map( A1 => n17816, A2 => n18056, B1 => n9137, B2 => 
                           n17812, ZN => n2930);
   U15703 : OAI22_X1 port map( A1 => n17816, A2 => n18059, B1 => n9120, B2 => 
                           n17812, ZN => n2931);
   U15704 : OAI22_X1 port map( A1 => n17816, A2 => n18062, B1 => n9103, B2 => 
                           n17812, ZN => n2932);
   U15705 : OAI22_X1 port map( A1 => n17817, A2 => n18065, B1 => n9086, B2 => 
                           n17812, ZN => n2933);
   U15706 : OAI22_X1 port map( A1 => n17817, A2 => n18068, B1 => n9069, B2 => 
                           n17812, ZN => n2934);
   U15707 : OAI22_X1 port map( A1 => n17817, A2 => n18071, B1 => n9052, B2 => 
                           n17812, ZN => n2935);
   U15708 : OAI22_X1 port map( A1 => n17817, A2 => n18074, B1 => n9035, B2 => 
                           n17812, ZN => n2936);
   U15709 : OAI22_X1 port map( A1 => n17768, A2 => n18006, B1 => n9429, B2 => 
                           n17767, ZN => n2753);
   U15710 : OAI22_X1 port map( A1 => n17768, A2 => n18009, B1 => n9412, B2 => 
                           n17767, ZN => n2754);
   U15711 : OAI22_X1 port map( A1 => n17768, A2 => n18012, B1 => n9395, B2 => 
                           n17767, ZN => n2755);
   U15712 : OAI22_X1 port map( A1 => n17768, A2 => n18015, B1 => n9378, B2 => 
                           n17767, ZN => n2756);
   U15713 : OAI22_X1 port map( A1 => n17768, A2 => n18018, B1 => n9361, B2 => 
                           n17767, ZN => n2757);
   U15714 : OAI22_X1 port map( A1 => n17769, A2 => n18021, B1 => n9344, B2 => 
                           n17767, ZN => n2758);
   U15715 : OAI22_X1 port map( A1 => n17769, A2 => n18024, B1 => n9327, B2 => 
                           n17767, ZN => n2759);
   U15716 : OAI22_X1 port map( A1 => n17769, A2 => n18027, B1 => n9310, B2 => 
                           n17767, ZN => n2760);
   U15717 : OAI22_X1 port map( A1 => n17769, A2 => n18030, B1 => n9293, B2 => 
                           n17767, ZN => n2761);
   U15718 : OAI22_X1 port map( A1 => n17769, A2 => n18033, B1 => n9276, B2 => 
                           n17767, ZN => n2762);
   U15719 : OAI22_X1 port map( A1 => n17770, A2 => n18036, B1 => n9259, B2 => 
                           n17767, ZN => n2763);
   U15720 : OAI22_X1 port map( A1 => n17770, A2 => n18039, B1 => n9242, B2 => 
                           n17767, ZN => n2764);
   U15721 : OAI22_X1 port map( A1 => n17770, A2 => n18042, B1 => n9225, B2 => 
                           n14669, ZN => n2765);
   U15722 : OAI22_X1 port map( A1 => n17770, A2 => n18045, B1 => n9208, B2 => 
                           n14669, ZN => n2766);
   U15723 : OAI22_X1 port map( A1 => n17770, A2 => n18048, B1 => n9191, B2 => 
                           n14669, ZN => n2767);
   U15724 : OAI22_X1 port map( A1 => n17771, A2 => n18051, B1 => n9174, B2 => 
                           n17767, ZN => n2768);
   U15725 : OAI22_X1 port map( A1 => n17771, A2 => n18054, B1 => n9157, B2 => 
                           n17767, ZN => n2769);
   U15726 : OAI22_X1 port map( A1 => n17771, A2 => n18057, B1 => n9140, B2 => 
                           n17767, ZN => n2770);
   U15727 : OAI22_X1 port map( A1 => n17771, A2 => n18060, B1 => n9123, B2 => 
                           n17767, ZN => n2771);
   U15728 : OAI22_X1 port map( A1 => n17771, A2 => n18063, B1 => n9106, B2 => 
                           n17767, ZN => n2772);
   U15729 : OAI22_X1 port map( A1 => n17772, A2 => n18066, B1 => n9089, B2 => 
                           n17767, ZN => n2773);
   U15730 : OAI22_X1 port map( A1 => n17772, A2 => n18069, B1 => n9072, B2 => 
                           n17767, ZN => n2774);
   U15731 : OAI22_X1 port map( A1 => n17772, A2 => n18072, B1 => n9055, B2 => 
                           n17767, ZN => n2775);
   U15732 : OAI22_X1 port map( A1 => n17772, A2 => n18075, B1 => n9038, B2 => 
                           n17767, ZN => n2776);
   U15733 : OAI22_X1 port map( A1 => n17759, A2 => n18006, B1 => n9428, B2 => 
                           n17758, ZN => n2721);
   U15734 : OAI22_X1 port map( A1 => n17759, A2 => n18009, B1 => n9411, B2 => 
                           n17758, ZN => n2722);
   U15735 : OAI22_X1 port map( A1 => n17759, A2 => n18012, B1 => n9394, B2 => 
                           n17758, ZN => n2723);
   U15736 : OAI22_X1 port map( A1 => n17759, A2 => n18015, B1 => n9377, B2 => 
                           n17758, ZN => n2724);
   U15737 : OAI22_X1 port map( A1 => n17759, A2 => n18018, B1 => n9360, B2 => 
                           n17758, ZN => n2725);
   U15738 : OAI22_X1 port map( A1 => n17760, A2 => n18021, B1 => n9343, B2 => 
                           n17758, ZN => n2726);
   U15739 : OAI22_X1 port map( A1 => n17760, A2 => n18024, B1 => n9326, B2 => 
                           n17758, ZN => n2727);
   U15740 : OAI22_X1 port map( A1 => n17760, A2 => n18027, B1 => n9309, B2 => 
                           n17758, ZN => n2728);
   U15741 : OAI22_X1 port map( A1 => n17760, A2 => n18030, B1 => n9292, B2 => 
                           n17758, ZN => n2729);
   U15742 : OAI22_X1 port map( A1 => n17760, A2 => n18033, B1 => n9275, B2 => 
                           n17758, ZN => n2730);
   U15743 : OAI22_X1 port map( A1 => n17761, A2 => n18036, B1 => n9258, B2 => 
                           n17758, ZN => n2731);
   U15744 : OAI22_X1 port map( A1 => n17761, A2 => n18039, B1 => n9241, B2 => 
                           n17758, ZN => n2732);
   U15745 : OAI22_X1 port map( A1 => n17761, A2 => n18042, B1 => n9224, B2 => 
                           n14670, ZN => n2733);
   U15746 : OAI22_X1 port map( A1 => n17761, A2 => n18045, B1 => n9207, B2 => 
                           n14670, ZN => n2734);
   U15747 : OAI22_X1 port map( A1 => n17761, A2 => n18048, B1 => n9190, B2 => 
                           n14670, ZN => n2735);
   U15748 : OAI22_X1 port map( A1 => n17762, A2 => n18051, B1 => n9173, B2 => 
                           n17758, ZN => n2736);
   U15749 : OAI22_X1 port map( A1 => n17762, A2 => n18054, B1 => n9156, B2 => 
                           n17758, ZN => n2737);
   U15750 : OAI22_X1 port map( A1 => n17762, A2 => n18057, B1 => n9139, B2 => 
                           n17758, ZN => n2738);
   U15751 : OAI22_X1 port map( A1 => n17762, A2 => n18060, B1 => n9122, B2 => 
                           n17758, ZN => n2739);
   U15752 : OAI22_X1 port map( A1 => n17762, A2 => n18063, B1 => n9105, B2 => 
                           n17758, ZN => n2740);
   U15753 : OAI22_X1 port map( A1 => n17763, A2 => n18066, B1 => n9088, B2 => 
                           n17758, ZN => n2741);
   U15754 : OAI22_X1 port map( A1 => n17763, A2 => n18069, B1 => n9071, B2 => 
                           n17758, ZN => n2742);
   U15755 : OAI22_X1 port map( A1 => n17763, A2 => n18072, B1 => n9054, B2 => 
                           n17758, ZN => n2743);
   U15756 : OAI22_X1 port map( A1 => n17763, A2 => n18075, B1 => n9037, B2 => 
                           n17758, ZN => n2744);
   U15757 : OAI22_X1 port map( A1 => n17732, A2 => n18006, B1 => n9431, B2 => 
                           n17731, ZN => n2625);
   U15758 : OAI22_X1 port map( A1 => n17732, A2 => n18009, B1 => n9414, B2 => 
                           n17731, ZN => n2626);
   U15759 : OAI22_X1 port map( A1 => n17732, A2 => n18012, B1 => n9397, B2 => 
                           n17731, ZN => n2627);
   U15760 : OAI22_X1 port map( A1 => n17732, A2 => n18015, B1 => n9380, B2 => 
                           n17731, ZN => n2628);
   U15761 : OAI22_X1 port map( A1 => n17732, A2 => n18018, B1 => n9363, B2 => 
                           n17731, ZN => n2629);
   U15762 : OAI22_X1 port map( A1 => n17733, A2 => n18021, B1 => n9346, B2 => 
                           n17731, ZN => n2630);
   U15763 : OAI22_X1 port map( A1 => n17733, A2 => n18024, B1 => n9329, B2 => 
                           n17731, ZN => n2631);
   U15764 : OAI22_X1 port map( A1 => n17733, A2 => n18027, B1 => n9312, B2 => 
                           n17731, ZN => n2632);
   U15765 : OAI22_X1 port map( A1 => n17733, A2 => n18030, B1 => n9295, B2 => 
                           n17731, ZN => n2633);
   U15766 : OAI22_X1 port map( A1 => n17733, A2 => n18033, B1 => n9278, B2 => 
                           n17731, ZN => n2634);
   U15767 : OAI22_X1 port map( A1 => n17734, A2 => n18036, B1 => n9261, B2 => 
                           n17731, ZN => n2635);
   U15768 : OAI22_X1 port map( A1 => n17734, A2 => n18039, B1 => n9244, B2 => 
                           n17731, ZN => n2636);
   U15769 : OAI22_X1 port map( A1 => n17734, A2 => n18042, B1 => n9227, B2 => 
                           n14673, ZN => n2637);
   U15770 : OAI22_X1 port map( A1 => n17734, A2 => n18045, B1 => n9210, B2 => 
                           n14673, ZN => n2638);
   U15771 : OAI22_X1 port map( A1 => n17734, A2 => n18048, B1 => n9193, B2 => 
                           n14673, ZN => n2639);
   U15772 : OAI22_X1 port map( A1 => n17735, A2 => n18051, B1 => n9176, B2 => 
                           n17731, ZN => n2640);
   U15773 : OAI22_X1 port map( A1 => n17735, A2 => n18054, B1 => n9159, B2 => 
                           n17731, ZN => n2641);
   U15774 : OAI22_X1 port map( A1 => n17735, A2 => n18057, B1 => n9142, B2 => 
                           n17731, ZN => n2642);
   U15775 : OAI22_X1 port map( A1 => n17735, A2 => n18060, B1 => n9125, B2 => 
                           n17731, ZN => n2643);
   U15776 : OAI22_X1 port map( A1 => n17735, A2 => n18063, B1 => n9108, B2 => 
                           n17731, ZN => n2644);
   U15777 : OAI22_X1 port map( A1 => n17736, A2 => n18066, B1 => n9091, B2 => 
                           n17731, ZN => n2645);
   U15778 : OAI22_X1 port map( A1 => n17736, A2 => n18069, B1 => n9074, B2 => 
                           n17731, ZN => n2646);
   U15779 : OAI22_X1 port map( A1 => n17736, A2 => n18072, B1 => n9057, B2 => 
                           n17731, ZN => n2647);
   U15780 : OAI22_X1 port map( A1 => n17736, A2 => n18075, B1 => n9040, B2 => 
                           n17731, ZN => n2648);
   U15781 : OAI21_X1 port map( B1 => n9415, B2 => n17615, A => n15950, ZN => 
                           n2529);
   U15782 : OAI21_X1 port map( B1 => n15951, B2 => n15952, A => n17618, ZN => 
                           n15950);
   U15783 : NAND4_X1 port map( A1 => n15969, A2 => n15970, A3 => n15971, A4 => 
                           n15972, ZN => n15951);
   U15784 : NAND4_X1 port map( A1 => n15953, A2 => n15954, A3 => n15955, A4 => 
                           n15956, ZN => n15952);
   U15785 : OAI21_X1 port map( B1 => n9398, B2 => n17615, A => n15931, ZN => 
                           n2530);
   U15786 : OAI21_X1 port map( B1 => n15932, B2 => n15933, A => n17618, ZN => 
                           n15931);
   U15787 : NAND4_X1 port map( A1 => n15942, A2 => n15943, A3 => n15944, A4 => 
                           n15945, ZN => n15932);
   U15788 : NAND4_X1 port map( A1 => n15934, A2 => n15935, A3 => n15936, A4 => 
                           n15937, ZN => n15933);
   U15789 : OAI21_X1 port map( B1 => n9381, B2 => n17615, A => n15912, ZN => 
                           n2531);
   U15790 : OAI21_X1 port map( B1 => n15913, B2 => n15914, A => n17617, ZN => 
                           n15912);
   U15791 : NAND4_X1 port map( A1 => n15923, A2 => n15924, A3 => n15925, A4 => 
                           n15926, ZN => n15913);
   U15792 : NAND4_X1 port map( A1 => n15915, A2 => n15916, A3 => n15917, A4 => 
                           n15918, ZN => n15914);
   U15793 : OAI21_X1 port map( B1 => n9364, B2 => n17615, A => n15893, ZN => 
                           n2532);
   U15794 : OAI21_X1 port map( B1 => n15894, B2 => n15895, A => n17617, ZN => 
                           n15893);
   U15795 : NAND4_X1 port map( A1 => n15904, A2 => n15905, A3 => n15906, A4 => 
                           n15907, ZN => n15894);
   U15796 : NAND4_X1 port map( A1 => n15896, A2 => n15897, A3 => n15898, A4 => 
                           n15899, ZN => n15895);
   U15797 : OAI21_X1 port map( B1 => n9347, B2 => n17615, A => n15874, ZN => 
                           n2533);
   U15798 : OAI21_X1 port map( B1 => n15875, B2 => n15876, A => n17617, ZN => 
                           n15874);
   U15799 : NAND4_X1 port map( A1 => n15885, A2 => n15886, A3 => n15887, A4 => 
                           n15888, ZN => n15875);
   U15800 : NAND4_X1 port map( A1 => n15877, A2 => n15878, A3 => n15879, A4 => 
                           n15880, ZN => n15876);
   U15801 : OAI21_X1 port map( B1 => n9330, B2 => n17615, A => n15855, ZN => 
                           n2534);
   U15802 : OAI21_X1 port map( B1 => n15856, B2 => n15857, A => n17616, ZN => 
                           n15855);
   U15803 : NAND4_X1 port map( A1 => n15866, A2 => n15867, A3 => n15868, A4 => 
                           n15869, ZN => n15856);
   U15804 : NAND4_X1 port map( A1 => n15858, A2 => n15859, A3 => n15860, A4 => 
                           n15861, ZN => n15857);
   U15805 : OAI21_X1 port map( B1 => n9313, B2 => n17615, A => n15836, ZN => 
                           n2535);
   U15806 : OAI21_X1 port map( B1 => n15837, B2 => n15838, A => n17617, ZN => 
                           n15836);
   U15807 : NAND4_X1 port map( A1 => n15847, A2 => n15848, A3 => n15849, A4 => 
                           n15850, ZN => n15837);
   U15808 : NAND4_X1 port map( A1 => n15839, A2 => n15840, A3 => n15841, A4 => 
                           n15842, ZN => n15838);
   U15809 : OAI21_X1 port map( B1 => n9279, B2 => n17615, A => n15798, ZN => 
                           n2537);
   U15810 : OAI21_X1 port map( B1 => n15799, B2 => n15800, A => n17616, ZN => 
                           n15798);
   U15811 : NAND4_X1 port map( A1 => n15809, A2 => n15810, A3 => n15811, A4 => 
                           n15812, ZN => n15799);
   U15812 : NAND4_X1 port map( A1 => n15801, A2 => n15802, A3 => n15803, A4 => 
                           n15804, ZN => n15800);
   U15813 : OAI21_X1 port map( B1 => n8887, B2 => n17717, A => n15297, ZN => 
                           n2561);
   U15814 : OAI21_X1 port map( B1 => n15298, B2 => n15299, A => n17720, ZN => 
                           n15297);
   U15815 : NAND4_X1 port map( A1 => n15316, A2 => n15317, A3 => n15318, A4 => 
                           n15319, ZN => n15298);
   U15816 : NAND4_X1 port map( A1 => n15300, A2 => n15301, A3 => n15302, A4 => 
                           n15303, ZN => n15299);
   U15817 : OAI21_X1 port map( B1 => n8886, B2 => n17717, A => n15278, ZN => 
                           n2562);
   U15818 : OAI21_X1 port map( B1 => n15279, B2 => n15280, A => n17720, ZN => 
                           n15278);
   U15819 : NAND4_X1 port map( A1 => n15289, A2 => n15290, A3 => n15291, A4 => 
                           n15292, ZN => n15279);
   U15820 : NAND4_X1 port map( A1 => n15281, A2 => n15282, A3 => n15283, A4 => 
                           n15284, ZN => n15280);
   U15821 : OAI21_X1 port map( B1 => n8885, B2 => n17717, A => n15259, ZN => 
                           n2563);
   U15822 : OAI21_X1 port map( B1 => n15260, B2 => n15261, A => n17719, ZN => 
                           n15259);
   U15823 : NAND4_X1 port map( A1 => n15270, A2 => n15271, A3 => n15272, A4 => 
                           n15273, ZN => n15260);
   U15824 : NAND4_X1 port map( A1 => n15262, A2 => n15263, A3 => n15264, A4 => 
                           n15265, ZN => n15261);
   U15825 : OAI21_X1 port map( B1 => n8884, B2 => n17717, A => n15240, ZN => 
                           n2564);
   U15826 : OAI21_X1 port map( B1 => n15241, B2 => n15242, A => n17719, ZN => 
                           n15240);
   U15827 : NAND4_X1 port map( A1 => n15251, A2 => n15252, A3 => n15253, A4 => 
                           n15254, ZN => n15241);
   U15828 : NAND4_X1 port map( A1 => n15243, A2 => n15244, A3 => n15245, A4 => 
                           n15246, ZN => n15242);
   U15829 : OAI21_X1 port map( B1 => n8883, B2 => n17717, A => n15221, ZN => 
                           n2565);
   U15830 : OAI21_X1 port map( B1 => n15222, B2 => n15223, A => n17719, ZN => 
                           n15221);
   U15831 : NAND4_X1 port map( A1 => n15232, A2 => n15233, A3 => n15234, A4 => 
                           n15235, ZN => n15222);
   U15832 : NAND4_X1 port map( A1 => n15224, A2 => n15225, A3 => n15226, A4 => 
                           n15227, ZN => n15223);
   U15833 : OAI21_X1 port map( B1 => n8882, B2 => n17717, A => n15202, ZN => 
                           n2566);
   U15834 : OAI21_X1 port map( B1 => n15203, B2 => n15204, A => n17718, ZN => 
                           n15202);
   U15835 : NAND4_X1 port map( A1 => n15213, A2 => n15214, A3 => n15215, A4 => 
                           n15216, ZN => n15203);
   U15836 : NAND4_X1 port map( A1 => n15205, A2 => n15206, A3 => n15207, A4 => 
                           n15208, ZN => n15204);
   U15837 : OAI21_X1 port map( B1 => n8881, B2 => n17717, A => n15183, ZN => 
                           n2567);
   U15838 : OAI21_X1 port map( B1 => n15184, B2 => n15185, A => n17719, ZN => 
                           n15183);
   U15839 : NAND4_X1 port map( A1 => n15194, A2 => n15195, A3 => n15196, A4 => 
                           n15197, ZN => n15184);
   U15840 : NAND4_X1 port map( A1 => n15186, A2 => n15187, A3 => n15188, A4 => 
                           n15189, ZN => n15185);
   U15841 : OAI21_X1 port map( B1 => n8879, B2 => n17717, A => n15145, ZN => 
                           n2569);
   U15842 : OAI21_X1 port map( B1 => n15146, B2 => n15147, A => n17718, ZN => 
                           n15145);
   U15843 : NAND4_X1 port map( A1 => n15156, A2 => n15157, A3 => n15158, A4 => 
                           n15159, ZN => n15146);
   U15844 : NAND4_X1 port map( A1 => n15148, A2 => n15149, A3 => n15150, A4 => 
                           n15151, ZN => n15147);
   U15845 : OAI21_X1 port map( B1 => n9296, B2 => n17614, A => n15817, ZN => 
                           n2536);
   U15846 : OAI21_X1 port map( B1 => n15818, B2 => n15819, A => n17616, ZN => 
                           n15817);
   U15847 : NAND4_X1 port map( A1 => n15828, A2 => n15829, A3 => n15830, A4 => 
                           n15831, ZN => n15818);
   U15848 : NAND4_X1 port map( A1 => n15820, A2 => n15821, A3 => n15822, A4 => 
                           n15823, ZN => n15819);
   U15849 : OAI21_X1 port map( B1 => n9262, B2 => n17614, A => n15779, ZN => 
                           n2538);
   U15850 : OAI21_X1 port map( B1 => n15780, B2 => n15781, A => n17616, ZN => 
                           n15779);
   U15851 : NAND4_X1 port map( A1 => n15790, A2 => n15791, A3 => n15792, A4 => 
                           n15793, ZN => n15780);
   U15852 : NAND4_X1 port map( A1 => n15782, A2 => n15783, A3 => n15784, A4 => 
                           n15785, ZN => n15781);
   U15853 : OAI21_X1 port map( B1 => n9245, B2 => n17614, A => n15760, ZN => 
                           n2539);
   U15854 : OAI21_X1 port map( B1 => n15761, B2 => n15762, A => n17615, ZN => 
                           n15760);
   U15855 : NAND4_X1 port map( A1 => n15771, A2 => n15772, A3 => n15773, A4 => 
                           n15774, ZN => n15761);
   U15856 : NAND4_X1 port map( A1 => n15763, A2 => n15764, A3 => n15765, A4 => 
                           n15766, ZN => n15762);
   U15857 : OAI21_X1 port map( B1 => n9228, B2 => n17614, A => n15741, ZN => 
                           n2540);
   U15858 : OAI21_X1 port map( B1 => n15742, B2 => n15743, A => n17615, ZN => 
                           n15741);
   U15859 : NAND4_X1 port map( A1 => n15752, A2 => n15753, A3 => n15754, A4 => 
                           n15755, ZN => n15742);
   U15860 : NAND4_X1 port map( A1 => n15744, A2 => n15745, A3 => n15746, A4 => 
                           n15747, ZN => n15743);
   U15861 : OAI21_X1 port map( B1 => n9211, B2 => n17614, A => n15722, ZN => 
                           n2541);
   U15862 : OAI21_X1 port map( B1 => n15723, B2 => n15724, A => n17616, ZN => 
                           n15722);
   U15863 : NAND4_X1 port map( A1 => n15733, A2 => n15734, A3 => n15735, A4 => 
                           n15736, ZN => n15723);
   U15864 : NAND4_X1 port map( A1 => n15725, A2 => n15726, A3 => n15727, A4 => 
                           n15728, ZN => n15724);
   U15865 : OAI21_X1 port map( B1 => n9194, B2 => n17614, A => n15703, ZN => 
                           n2542);
   U15866 : OAI21_X1 port map( B1 => n15704, B2 => n15705, A => n17615, ZN => 
                           n15703);
   U15867 : NAND4_X1 port map( A1 => n15714, A2 => n15715, A3 => n15716, A4 => 
                           n15717, ZN => n15704);
   U15868 : NAND4_X1 port map( A1 => n15706, A2 => n15707, A3 => n15708, A4 => 
                           n15709, ZN => n15705);
   U15869 : OAI21_X1 port map( B1 => n9177, B2 => n17614, A => n15684, ZN => 
                           n2543);
   U15870 : OAI21_X1 port map( B1 => n15685, B2 => n15686, A => n17615, ZN => 
                           n15684);
   U15871 : NAND4_X1 port map( A1 => n15695, A2 => n15696, A3 => n15697, A4 => 
                           n15698, ZN => n15685);
   U15872 : NAND4_X1 port map( A1 => n15687, A2 => n15688, A3 => n15689, A4 => 
                           n15690, ZN => n15686);
   U15873 : OAI21_X1 port map( B1 => n9160, B2 => n17614, A => n15665, ZN => 
                           n2544);
   U15874 : OAI21_X1 port map( B1 => n15666, B2 => n15667, A => n17616, ZN => 
                           n15665);
   U15875 : NAND4_X1 port map( A1 => n15676, A2 => n15677, A3 => n15678, A4 => 
                           n15679, ZN => n15666);
   U15876 : NAND4_X1 port map( A1 => n15668, A2 => n15669, A3 => n15670, A4 => 
                           n15671, ZN => n15667);
   U15877 : OAI21_X1 port map( B1 => n9143, B2 => n17614, A => n15646, ZN => 
                           n2545);
   U15878 : OAI21_X1 port map( B1 => n15647, B2 => n15648, A => n17616, ZN => 
                           n15646);
   U15879 : NAND4_X1 port map( A1 => n15657, A2 => n15658, A3 => n15659, A4 => 
                           n15660, ZN => n15647);
   U15880 : NAND4_X1 port map( A1 => n15649, A2 => n15650, A3 => n15651, A4 => 
                           n15652, ZN => n15648);
   U15881 : OAI21_X1 port map( B1 => n9126, B2 => n17614, A => n15627, ZN => 
                           n2546);
   U15882 : OAI21_X1 port map( B1 => n15628, B2 => n15629, A => n17616, ZN => 
                           n15627);
   U15883 : NAND4_X1 port map( A1 => n15638, A2 => n15639, A3 => n15640, A4 => 
                           n15641, ZN => n15628);
   U15884 : NAND4_X1 port map( A1 => n15630, A2 => n15631, A3 => n15632, A4 => 
                           n15633, ZN => n15629);
   U15885 : OAI21_X1 port map( B1 => n9109, B2 => n17614, A => n15608, ZN => 
                           n2547);
   U15886 : OAI21_X1 port map( B1 => n15609, B2 => n15610, A => n17616, ZN => 
                           n15608);
   U15887 : NAND4_X1 port map( A1 => n15619, A2 => n15620, A3 => n15621, A4 => 
                           n15622, ZN => n15609);
   U15888 : NAND4_X1 port map( A1 => n15611, A2 => n15612, A3 => n15613, A4 => 
                           n15614, ZN => n15610);
   U15889 : OAI21_X1 port map( B1 => n9092, B2 => n17613, A => n15589, ZN => 
                           n2548);
   U15890 : OAI21_X1 port map( B1 => n15590, B2 => n15591, A => n17616, ZN => 
                           n15589);
   U15891 : NAND4_X1 port map( A1 => n15600, A2 => n15601, A3 => n15602, A4 => 
                           n15603, ZN => n15590);
   U15892 : NAND4_X1 port map( A1 => n15592, A2 => n15593, A3 => n15594, A4 => 
                           n15595, ZN => n15591);
   U15893 : OAI21_X1 port map( B1 => n9075, B2 => n17613, A => n15570, ZN => 
                           n2549);
   U15894 : OAI21_X1 port map( B1 => n15571, B2 => n15572, A => n17616, ZN => 
                           n15570);
   U15895 : NAND4_X1 port map( A1 => n15581, A2 => n15582, A3 => n15583, A4 => 
                           n15584, ZN => n15571);
   U15896 : NAND4_X1 port map( A1 => n15573, A2 => n15574, A3 => n15575, A4 => 
                           n15576, ZN => n15572);
   U15897 : OAI21_X1 port map( B1 => n9058, B2 => n17613, A => n15551, ZN => 
                           n2550);
   U15898 : OAI21_X1 port map( B1 => n15552, B2 => n15553, A => n17617, ZN => 
                           n15551);
   U15899 : NAND4_X1 port map( A1 => n15562, A2 => n15563, A3 => n15564, A4 => 
                           n15565, ZN => n15552);
   U15900 : NAND4_X1 port map( A1 => n15554, A2 => n15555, A3 => n15556, A4 => 
                           n15557, ZN => n15553);
   U15901 : OAI21_X1 port map( B1 => n9041, B2 => n17613, A => n15532, ZN => 
                           n2551);
   U15902 : OAI21_X1 port map( B1 => n15533, B2 => n15534, A => n17616, ZN => 
                           n15532);
   U15903 : NAND4_X1 port map( A1 => n15543, A2 => n15544, A3 => n15545, A4 => 
                           n15546, ZN => n15533);
   U15904 : NAND4_X1 port map( A1 => n15535, A2 => n15536, A3 => n15537, A4 => 
                           n15538, ZN => n15534);
   U15905 : OAI21_X1 port map( B1 => n9024, B2 => n17613, A => n15513, ZN => 
                           n2552);
   U15906 : OAI21_X1 port map( B1 => n15514, B2 => n15515, A => n17617, ZN => 
                           n15513);
   U15907 : NAND4_X1 port map( A1 => n15524, A2 => n15525, A3 => n15526, A4 => 
                           n15527, ZN => n15514);
   U15908 : NAND4_X1 port map( A1 => n15516, A2 => n15517, A3 => n15518, A4 => 
                           n15519, ZN => n15515);
   U15909 : OAI21_X1 port map( B1 => n9007, B2 => n17613, A => n15494, ZN => 
                           n2553);
   U15910 : OAI21_X1 port map( B1 => n15495, B2 => n15496, A => n17617, ZN => 
                           n15494);
   U15911 : NAND4_X1 port map( A1 => n15505, A2 => n15506, A3 => n15507, A4 => 
                           n15508, ZN => n15495);
   U15912 : NAND4_X1 port map( A1 => n15497, A2 => n15498, A3 => n15499, A4 => 
                           n15500, ZN => n15496);
   U15913 : OAI21_X1 port map( B1 => n8990, B2 => n17613, A => n15475, ZN => 
                           n2554);
   U15914 : OAI21_X1 port map( B1 => n15476, B2 => n15477, A => n17617, ZN => 
                           n15475);
   U15915 : NAND4_X1 port map( A1 => n15486, A2 => n15487, A3 => n15488, A4 => 
                           n15489, ZN => n15476);
   U15916 : NAND4_X1 port map( A1 => n15478, A2 => n15479, A3 => n15480, A4 => 
                           n15481, ZN => n15477);
   U15917 : OAI21_X1 port map( B1 => n8973, B2 => n17613, A => n15456, ZN => 
                           n2555);
   U15918 : OAI21_X1 port map( B1 => n15457, B2 => n15458, A => n17617, ZN => 
                           n15456);
   U15919 : NAND4_X1 port map( A1 => n15467, A2 => n15468, A3 => n15469, A4 => 
                           n15470, ZN => n15457);
   U15920 : NAND4_X1 port map( A1 => n15459, A2 => n15460, A3 => n15461, A4 => 
                           n15462, ZN => n15458);
   U15921 : OAI21_X1 port map( B1 => n8956, B2 => n17613, A => n15437, ZN => 
                           n2556);
   U15922 : OAI21_X1 port map( B1 => n15438, B2 => n15439, A => n17617, ZN => 
                           n15437);
   U15923 : NAND4_X1 port map( A1 => n15448, A2 => n15449, A3 => n15450, A4 => 
                           n15451, ZN => n15438);
   U15924 : NAND4_X1 port map( A1 => n15440, A2 => n15441, A3 => n15442, A4 => 
                           n15443, ZN => n15439);
   U15925 : OAI21_X1 port map( B1 => n8939, B2 => n17613, A => n15418, ZN => 
                           n2557);
   U15926 : OAI21_X1 port map( B1 => n15419, B2 => n15420, A => n17617, ZN => 
                           n15418);
   U15927 : NAND4_X1 port map( A1 => n15429, A2 => n15430, A3 => n15431, A4 => 
                           n15432, ZN => n15419);
   U15928 : NAND4_X1 port map( A1 => n15421, A2 => n15422, A3 => n15423, A4 => 
                           n15424, ZN => n15420);
   U15929 : OAI21_X1 port map( B1 => n8922, B2 => n17613, A => n15399, ZN => 
                           n2558);
   U15930 : OAI21_X1 port map( B1 => n15400, B2 => n15401, A => n17617, ZN => 
                           n15399);
   U15931 : NAND4_X1 port map( A1 => n15410, A2 => n15411, A3 => n15412, A4 => 
                           n15413, ZN => n15400);
   U15932 : NAND4_X1 port map( A1 => n15402, A2 => n15403, A3 => n15404, A4 => 
                           n15405, ZN => n15401);
   U15933 : OAI21_X1 port map( B1 => n8905, B2 => n17613, A => n15380, ZN => 
                           n2559);
   U15934 : OAI21_X1 port map( B1 => n15381, B2 => n15382, A => n17618, ZN => 
                           n15380);
   U15935 : NAND4_X1 port map( A1 => n15391, A2 => n15392, A3 => n15393, A4 => 
                           n15394, ZN => n15381);
   U15936 : NAND4_X1 port map( A1 => n15383, A2 => n15384, A3 => n15385, A4 => 
                           n15386, ZN => n15382);
   U15937 : OAI21_X1 port map( B1 => n8888, B2 => n17614, A => n15329, ZN => 
                           n2560);
   U15938 : OAI21_X1 port map( B1 => n15330, B2 => n15331, A => n17618, ZN => 
                           n15329);
   U15939 : NAND4_X1 port map( A1 => n15356, A2 => n15357, A3 => n15358, A4 => 
                           n15359, ZN => n15330);
   U15940 : NAND4_X1 port map( A1 => n15332, A2 => n15333, A3 => n15334, A4 => 
                           n15335, ZN => n15331);
   U15941 : OAI21_X1 port map( B1 => n8880, B2 => n17716, A => n15164, ZN => 
                           n2568);
   U15942 : OAI21_X1 port map( B1 => n15165, B2 => n15166, A => n17718, ZN => 
                           n15164);
   U15943 : NAND4_X1 port map( A1 => n15175, A2 => n15176, A3 => n15177, A4 => 
                           n15178, ZN => n15165);
   U15944 : NAND4_X1 port map( A1 => n15167, A2 => n15168, A3 => n15169, A4 => 
                           n15170, ZN => n15166);
   U15945 : OAI21_X1 port map( B1 => n8878, B2 => n17716, A => n15126, ZN => 
                           n2570);
   U15946 : OAI21_X1 port map( B1 => n15127, B2 => n15128, A => n17718, ZN => 
                           n15126);
   U15947 : NAND4_X1 port map( A1 => n15137, A2 => n15138, A3 => n15139, A4 => 
                           n15140, ZN => n15127);
   U15948 : NAND4_X1 port map( A1 => n15129, A2 => n15130, A3 => n15131, A4 => 
                           n15132, ZN => n15128);
   U15949 : OAI21_X1 port map( B1 => n8877, B2 => n17716, A => n15107, ZN => 
                           n2571);
   U15950 : OAI21_X1 port map( B1 => n15108, B2 => n15109, A => n17717, ZN => 
                           n15107);
   U15951 : NAND4_X1 port map( A1 => n15118, A2 => n15119, A3 => n15120, A4 => 
                           n15121, ZN => n15108);
   U15952 : NAND4_X1 port map( A1 => n15110, A2 => n15111, A3 => n15112, A4 => 
                           n15113, ZN => n15109);
   U15953 : OAI21_X1 port map( B1 => n8876, B2 => n17716, A => n15088, ZN => 
                           n2572);
   U15954 : OAI21_X1 port map( B1 => n15089, B2 => n15090, A => n17717, ZN => 
                           n15088);
   U15955 : NAND4_X1 port map( A1 => n15099, A2 => n15100, A3 => n15101, A4 => 
                           n15102, ZN => n15089);
   U15956 : NAND4_X1 port map( A1 => n15091, A2 => n15092, A3 => n15093, A4 => 
                           n15094, ZN => n15090);
   U15957 : OAI21_X1 port map( B1 => n8875, B2 => n17716, A => n15069, ZN => 
                           n2573);
   U15958 : OAI21_X1 port map( B1 => n15070, B2 => n15071, A => n17718, ZN => 
                           n15069);
   U15959 : NAND4_X1 port map( A1 => n15080, A2 => n15081, A3 => n15082, A4 => 
                           n15083, ZN => n15070);
   U15960 : NAND4_X1 port map( A1 => n15072, A2 => n15073, A3 => n15074, A4 => 
                           n15075, ZN => n15071);
   U15961 : OAI21_X1 port map( B1 => n8874, B2 => n17716, A => n15050, ZN => 
                           n2574);
   U15962 : OAI21_X1 port map( B1 => n15051, B2 => n15052, A => n17717, ZN => 
                           n15050);
   U15963 : NAND4_X1 port map( A1 => n15061, A2 => n15062, A3 => n15063, A4 => 
                           n15064, ZN => n15051);
   U15964 : NAND4_X1 port map( A1 => n15053, A2 => n15054, A3 => n15055, A4 => 
                           n15056, ZN => n15052);
   U15965 : OAI21_X1 port map( B1 => n8873, B2 => n17716, A => n15031, ZN => 
                           n2575);
   U15966 : OAI21_X1 port map( B1 => n15032, B2 => n15033, A => n17717, ZN => 
                           n15031);
   U15967 : NAND4_X1 port map( A1 => n15042, A2 => n15043, A3 => n15044, A4 => 
                           n15045, ZN => n15032);
   U15968 : NAND4_X1 port map( A1 => n15034, A2 => n15035, A3 => n15036, A4 => 
                           n15037, ZN => n15033);
   U15969 : OAI21_X1 port map( B1 => n8872, B2 => n17716, A => n15012, ZN => 
                           n2576);
   U15970 : OAI21_X1 port map( B1 => n15013, B2 => n15014, A => n17718, ZN => 
                           n15012);
   U15971 : NAND4_X1 port map( A1 => n15023, A2 => n15024, A3 => n15025, A4 => 
                           n15026, ZN => n15013);
   U15972 : NAND4_X1 port map( A1 => n15015, A2 => n15016, A3 => n15017, A4 => 
                           n15018, ZN => n15014);
   U15973 : OAI21_X1 port map( B1 => n8871, B2 => n17716, A => n14993, ZN => 
                           n2577);
   U15974 : OAI21_X1 port map( B1 => n14994, B2 => n14995, A => n17718, ZN => 
                           n14993);
   U15975 : NAND4_X1 port map( A1 => n15004, A2 => n15005, A3 => n15006, A4 => 
                           n15007, ZN => n14994);
   U15976 : NAND4_X1 port map( A1 => n14996, A2 => n14997, A3 => n14998, A4 => 
                           n14999, ZN => n14995);
   U15977 : OAI21_X1 port map( B1 => n8870, B2 => n17716, A => n14974, ZN => 
                           n2578);
   U15978 : OAI21_X1 port map( B1 => n14975, B2 => n14976, A => n17718, ZN => 
                           n14974);
   U15979 : NAND4_X1 port map( A1 => n14985, A2 => n14986, A3 => n14987, A4 => 
                           n14988, ZN => n14975);
   U15980 : NAND4_X1 port map( A1 => n14977, A2 => n14978, A3 => n14979, A4 => 
                           n14980, ZN => n14976);
   U15981 : OAI21_X1 port map( B1 => n8869, B2 => n17716, A => n14955, ZN => 
                           n2579);
   U15982 : OAI21_X1 port map( B1 => n14956, B2 => n14957, A => n17718, ZN => 
                           n14955);
   U15983 : NAND4_X1 port map( A1 => n14966, A2 => n14967, A3 => n14968, A4 => 
                           n14969, ZN => n14956);
   U15984 : NAND4_X1 port map( A1 => n14958, A2 => n14959, A3 => n14960, A4 => 
                           n14961, ZN => n14957);
   U15985 : OAI21_X1 port map( B1 => n8868, B2 => n17715, A => n14936, ZN => 
                           n2580);
   U15986 : OAI21_X1 port map( B1 => n14937, B2 => n14938, A => n17718, ZN => 
                           n14936);
   U15987 : NAND4_X1 port map( A1 => n14947, A2 => n14948, A3 => n14949, A4 => 
                           n14950, ZN => n14937);
   U15988 : NAND4_X1 port map( A1 => n14939, A2 => n14940, A3 => n14941, A4 => 
                           n14942, ZN => n14938);
   U15989 : OAI21_X1 port map( B1 => n8867, B2 => n17715, A => n14917, ZN => 
                           n2581);
   U15990 : OAI21_X1 port map( B1 => n14918, B2 => n14919, A => n17718, ZN => 
                           n14917);
   U15991 : NAND4_X1 port map( A1 => n14928, A2 => n14929, A3 => n14930, A4 => 
                           n14931, ZN => n14918);
   U15992 : NAND4_X1 port map( A1 => n14920, A2 => n14921, A3 => n14922, A4 => 
                           n14923, ZN => n14919);
   U15993 : OAI21_X1 port map( B1 => n8866, B2 => n17715, A => n14898, ZN => 
                           n2582);
   U15994 : OAI21_X1 port map( B1 => n14899, B2 => n14900, A => n17719, ZN => 
                           n14898);
   U15995 : NAND4_X1 port map( A1 => n14909, A2 => n14910, A3 => n14911, A4 => 
                           n14912, ZN => n14899);
   U15996 : NAND4_X1 port map( A1 => n14901, A2 => n14902, A3 => n14903, A4 => 
                           n14904, ZN => n14900);
   U15997 : OAI21_X1 port map( B1 => n8865, B2 => n17715, A => n14879, ZN => 
                           n2583);
   U15998 : OAI21_X1 port map( B1 => n14880, B2 => n14881, A => n17718, ZN => 
                           n14879);
   U15999 : NAND4_X1 port map( A1 => n14890, A2 => n14891, A3 => n14892, A4 => 
                           n14893, ZN => n14880);
   U16000 : NAND4_X1 port map( A1 => n14882, A2 => n14883, A3 => n14884, A4 => 
                           n14885, ZN => n14881);
   U16001 : OAI21_X1 port map( B1 => n8864, B2 => n17715, A => n14860, ZN => 
                           n2584);
   U16002 : OAI21_X1 port map( B1 => n14861, B2 => n14862, A => n17719, ZN => 
                           n14860);
   U16003 : NAND4_X1 port map( A1 => n14871, A2 => n14872, A3 => n14873, A4 => 
                           n14874, ZN => n14861);
   U16004 : NAND4_X1 port map( A1 => n14863, A2 => n14864, A3 => n14865, A4 => 
                           n14866, ZN => n14862);
   U16005 : OAI21_X1 port map( B1 => n8863, B2 => n17715, A => n14841, ZN => 
                           n2585);
   U16006 : OAI21_X1 port map( B1 => n14842, B2 => n14843, A => n17719, ZN => 
                           n14841);
   U16007 : NAND4_X1 port map( A1 => n14852, A2 => n14853, A3 => n14854, A4 => 
                           n14855, ZN => n14842);
   U16008 : NAND4_X1 port map( A1 => n14844, A2 => n14845, A3 => n14846, A4 => 
                           n14847, ZN => n14843);
   U16009 : OAI21_X1 port map( B1 => n8862, B2 => n17715, A => n14822, ZN => 
                           n2586);
   U16010 : OAI21_X1 port map( B1 => n14823, B2 => n14824, A => n17719, ZN => 
                           n14822);
   U16011 : NAND4_X1 port map( A1 => n14833, A2 => n14834, A3 => n14835, A4 => 
                           n14836, ZN => n14823);
   U16012 : NAND4_X1 port map( A1 => n14825, A2 => n14826, A3 => n14827, A4 => 
                           n14828, ZN => n14824);
   U16013 : OAI21_X1 port map( B1 => n8861, B2 => n17715, A => n14803, ZN => 
                           n2587);
   U16014 : OAI21_X1 port map( B1 => n14804, B2 => n14805, A => n17719, ZN => 
                           n14803);
   U16015 : NAND4_X1 port map( A1 => n14814, A2 => n14815, A3 => n14816, A4 => 
                           n14817, ZN => n14804);
   U16016 : NAND4_X1 port map( A1 => n14806, A2 => n14807, A3 => n14808, A4 => 
                           n14809, ZN => n14805);
   U16017 : OAI21_X1 port map( B1 => n8860, B2 => n17715, A => n14784, ZN => 
                           n2588);
   U16018 : OAI21_X1 port map( B1 => n14785, B2 => n14786, A => n17719, ZN => 
                           n14784);
   U16019 : NAND4_X1 port map( A1 => n14795, A2 => n14796, A3 => n14797, A4 => 
                           n14798, ZN => n14785);
   U16020 : NAND4_X1 port map( A1 => n14787, A2 => n14788, A3 => n14789, A4 => 
                           n14790, ZN => n14786);
   U16021 : OAI21_X1 port map( B1 => n8859, B2 => n17715, A => n14765, ZN => 
                           n2589);
   U16022 : OAI21_X1 port map( B1 => n14766, B2 => n14767, A => n17719, ZN => 
                           n14765);
   U16023 : NAND4_X1 port map( A1 => n14776, A2 => n14777, A3 => n14778, A4 => 
                           n14779, ZN => n14766);
   U16024 : NAND4_X1 port map( A1 => n14768, A2 => n14769, A3 => n14770, A4 => 
                           n14771, ZN => n14767);
   U16025 : OAI21_X1 port map( B1 => n8858, B2 => n17715, A => n14746, ZN => 
                           n2590);
   U16026 : OAI21_X1 port map( B1 => n14747, B2 => n14748, A => n17719, ZN => 
                           n14746);
   U16027 : NAND4_X1 port map( A1 => n14757, A2 => n14758, A3 => n14759, A4 => 
                           n14760, ZN => n14747);
   U16028 : NAND4_X1 port map( A1 => n14749, A2 => n14750, A3 => n14751, A4 => 
                           n14752, ZN => n14748);
   U16029 : OAI21_X1 port map( B1 => n8857, B2 => n17715, A => n14727, ZN => 
                           n2591);
   U16030 : OAI21_X1 port map( B1 => n14728, B2 => n14729, A => n17720, ZN => 
                           n14727);
   U16031 : NAND4_X1 port map( A1 => n14738, A2 => n14739, A3 => n14740, A4 => 
                           n14741, ZN => n14728);
   U16032 : NAND4_X1 port map( A1 => n14730, A2 => n14731, A3 => n14732, A4 => 
                           n14733, ZN => n14729);
   U16033 : OAI21_X1 port map( B1 => n8856, B2 => n17716, A => n14676, ZN => 
                           n2592);
   U16034 : OAI21_X1 port map( B1 => n14677, B2 => n14678, A => n17720, ZN => 
                           n14676);
   U16035 : NAND4_X1 port map( A1 => n14703, A2 => n14704, A3 => n14705, A4 => 
                           n14706, ZN => n14677);
   U16036 : NAND4_X1 port map( A1 => n14679, A2 => n14680, A3 => n14681, A4 => 
                           n14682, ZN => n14678);
   U16037 : OAI22_X1 port map( A1 => n17831, A2 => n18005, B1 => n17830, B2 => 
                           n17493, ZN => n2977);
   U16038 : OAI22_X1 port map( A1 => n17831, A2 => n18008, B1 => n17830, B2 => 
                           n17494, ZN => n2978);
   U16039 : OAI22_X1 port map( A1 => n17831, A2 => n18011, B1 => n17830, B2 => 
                           n17495, ZN => n2979);
   U16040 : OAI22_X1 port map( A1 => n17831, A2 => n18014, B1 => n17830, B2 => 
                           n17496, ZN => n2980);
   U16041 : OAI22_X1 port map( A1 => n17831, A2 => n18017, B1 => n17830, B2 => 
                           n17497, ZN => n2981);
   U16042 : OAI22_X1 port map( A1 => n17832, A2 => n18020, B1 => n17830, B2 => 
                           n17498, ZN => n2982);
   U16043 : OAI22_X1 port map( A1 => n17832, A2 => n18023, B1 => n17830, B2 => 
                           n17499, ZN => n2983);
   U16044 : OAI22_X1 port map( A1 => n17832, A2 => n18026, B1 => n17830, B2 => 
                           n17500, ZN => n2984);
   U16045 : OAI22_X1 port map( A1 => n17832, A2 => n18029, B1 => n17830, B2 => 
                           n17501, ZN => n2985);
   U16046 : OAI22_X1 port map( A1 => n17832, A2 => n18032, B1 => n17830, B2 => 
                           n17502, ZN => n2986);
   U16047 : OAI22_X1 port map( A1 => n17833, A2 => n18035, B1 => n17830, B2 => 
                           n17503, ZN => n2987);
   U16048 : OAI22_X1 port map( A1 => n17833, A2 => n18038, B1 => n17830, B2 => 
                           n17504, ZN => n2988);
   U16049 : OAI22_X1 port map( A1 => n17833, A2 => n18041, B1 => n14661, B2 => 
                           n17505, ZN => n2989);
   U16050 : OAI22_X1 port map( A1 => n17833, A2 => n18044, B1 => n14661, B2 => 
                           n17506, ZN => n2990);
   U16051 : OAI22_X1 port map( A1 => n17833, A2 => n18047, B1 => n14661, B2 => 
                           n17507, ZN => n2991);
   U16052 : OAI22_X1 port map( A1 => n17834, A2 => n18050, B1 => n17830, B2 => 
                           n17508, ZN => n2992);
   U16053 : OAI22_X1 port map( A1 => n17834, A2 => n18053, B1 => n17830, B2 => 
                           n17509, ZN => n2993);
   U16054 : OAI22_X1 port map( A1 => n17834, A2 => n18056, B1 => n17830, B2 => 
                           n17510, ZN => n2994);
   U16055 : OAI22_X1 port map( A1 => n17834, A2 => n18059, B1 => n17830, B2 => 
                           n17511, ZN => n2995);
   U16056 : OAI22_X1 port map( A1 => n17834, A2 => n18062, B1 => n17830, B2 => 
                           n17512, ZN => n2996);
   U16057 : OAI22_X1 port map( A1 => n17835, A2 => n18065, B1 => n17830, B2 => 
                           n17513, ZN => n2997);
   U16058 : OAI22_X1 port map( A1 => n17835, A2 => n18068, B1 => n17830, B2 => 
                           n17514, ZN => n2998);
   U16059 : OAI22_X1 port map( A1 => n17835, A2 => n18071, B1 => n17830, B2 => 
                           n17515, ZN => n2999);
   U16060 : OAI22_X1 port map( A1 => n17835, A2 => n18074, B1 => n17830, B2 => 
                           n17516, ZN => n3000);
   U16061 : OAI22_X1 port map( A1 => n17835, A2 => n18077, B1 => n14661, B2 => 
                           n17045, ZN => n3001);
   U16062 : OAI22_X1 port map( A1 => n17836, A2 => n18080, B1 => n14661, B2 => 
                           n17046, ZN => n3002);
   U16063 : OAI22_X1 port map( A1 => n17836, A2 => n18083, B1 => n14661, B2 => 
                           n17047, ZN => n3003);
   U16064 : OAI22_X1 port map( A1 => n17836, A2 => n18086, B1 => n14661, B2 => 
                           n17048, ZN => n3004);
   U16065 : OAI22_X1 port map( A1 => n17836, A2 => n18089, B1 => n14661, B2 => 
                           n17049, ZN => n3005);
   U16066 : OAI22_X1 port map( A1 => n17836, A2 => n18092, B1 => n14661, B2 => 
                           n17050, ZN => n3006);
   U16067 : OAI22_X1 port map( A1 => n17837, A2 => n18095, B1 => n14661, B2 => 
                           n17051, ZN => n3007);
   U16068 : OAI22_X1 port map( A1 => n17837, A2 => n18107, B1 => n14661, B2 => 
                           n17052, ZN => n3008);
   U16069 : NOR3_X1 port map( A1 => ADDR_RD2(3), A2 => ADDR_RD2(4), A3 => 
                           n13572, ZN => n15974);
   U16070 : NOR3_X1 port map( A1 => ADDR_RD1(3), A2 => ADDR_RD1(4), A3 => 
                           n13568, ZN => n15321);
   U16071 : NOR2_X1 port map( A1 => n13571, A2 => ADDR_RD2(2), ZN => n15961);
   U16072 : NOR2_X1 port map( A1 => n13567, A2 => ADDR_RD1(2), ZN => n15308);
   U16073 : NOR2_X1 port map( A1 => n13570, A2 => ADDR_RD2(1), ZN => n15964);
   U16074 : NOR2_X1 port map( A1 => n13566, A2 => ADDR_RD1(1), ZN => n15311);
   U16075 : NOR3_X1 port map( A1 => ADDR_RD2(3), A2 => ADDR_RD2(4), A3 => 
                           ADDR_RD2(0), ZN => n15975);
   U16076 : NOR3_X1 port map( A1 => ADDR_RD1(3), A2 => ADDR_RD1(4), A3 => 
                           ADDR_RD1(0), ZN => n15322);
   U16077 : NOR3_X1 port map( A1 => n13572, A2 => ADDR_RD2(4), A3 => n13569, ZN
                           => n15979);
   U16078 : NOR3_X1 port map( A1 => n13568, A2 => ADDR_RD1(4), A3 => n13565, ZN
                           => n15326);
   U16079 : NOR3_X1 port map( A1 => ADDR_RD2(0), A2 => ADDR_RD2(4), A3 => 
                           n13569, ZN => n15978);
   U16080 : NOR3_X1 port map( A1 => ADDR_RD1(0), A2 => ADDR_RD1(4), A3 => 
                           n13565, ZN => n15325);
   U16081 : AND3_X1 port map( A1 => EN, A2 => n18111, A3 => RD2, ZN => n15328);
   U16082 : AND3_X1 port map( A1 => EN, A2 => n18111, A3 => RD1, ZN => n14675);
   U16083 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => n18111, ZN => n14629);
   U16084 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => n18111, ZN => n14628);
   U16085 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => n18111, ZN => n14627);
   U16086 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => n18111, ZN => n14626);
   U16087 : NAND2_X1 port map( A1 => DATA_IN(4), A2 => n18111, ZN => n14625);
   U16088 : NAND2_X1 port map( A1 => DATA_IN(5), A2 => n18111, ZN => n14624);
   U16089 : NAND2_X1 port map( A1 => DATA_IN(6), A2 => n18111, ZN => n14623);
   U16090 : NAND2_X1 port map( A1 => DATA_IN(7), A2 => n18111, ZN => n14622);
   U16091 : AND3_X1 port map( A1 => n13572, A2 => n13569, A3 => ADDR_RD2(4), ZN
                           => n15958);
   U16092 : AND3_X1 port map( A1 => n13568, A2 => n13565, A3 => ADDR_RD1(4), ZN
                           => n15305);
   U16093 : AND3_X1 port map( A1 => ADDR_RD2(0), A2 => n13569, A3 => 
                           ADDR_RD2(4), ZN => n15960);
   U16094 : AND3_X1 port map( A1 => ADDR_RD2(3), A2 => n13572, A3 => 
                           ADDR_RD2(4), ZN => n15966);
   U16095 : AND3_X1 port map( A1 => ADDR_RD1(0), A2 => n13565, A3 => 
                           ADDR_RD1(4), ZN => n15307);
   U16096 : AND3_X1 port map( A1 => ADDR_RD1(3), A2 => n13568, A3 => 
                           ADDR_RD1(4), ZN => n15313);
   U16097 : AND3_X1 port map( A1 => ADDR_RD2(3), A2 => ADDR_RD2(0), A3 => 
                           ADDR_RD2(4), ZN => n15967);
   U16098 : AND3_X1 port map( A1 => ADDR_RD1(3), A2 => ADDR_RD1(0), A3 => 
                           ADDR_RD1(4), ZN => n15314);
   U16099 : NAND2_X1 port map( A1 => DATA_IN(8), A2 => n18110, ZN => n14621);
   U16100 : NAND2_X1 port map( A1 => DATA_IN(9), A2 => n18110, ZN => n14620);
   U16101 : NAND2_X1 port map( A1 => DATA_IN(10), A2 => n18110, ZN => n14619);
   U16102 : NAND2_X1 port map( A1 => DATA_IN(11), A2 => n18110, ZN => n14618);
   U16103 : NAND2_X1 port map( A1 => DATA_IN(12), A2 => n18110, ZN => n14617);
   U16104 : NAND2_X1 port map( A1 => DATA_IN(13), A2 => n18110, ZN => n14616);
   U16105 : NAND2_X1 port map( A1 => DATA_IN(14), A2 => n18110, ZN => n14615);
   U16106 : NAND2_X1 port map( A1 => DATA_IN(15), A2 => n18110, ZN => n14614);
   U16107 : NAND2_X1 port map( A1 => DATA_IN(16), A2 => n18110, ZN => n14613);
   U16108 : NAND2_X1 port map( A1 => DATA_IN(17), A2 => n18110, ZN => n14612);
   U16109 : NAND2_X1 port map( A1 => DATA_IN(18), A2 => n18110, ZN => n14611);
   U16110 : NAND2_X1 port map( A1 => DATA_IN(19), A2 => n18110, ZN => n14610);
   U16111 : NAND2_X1 port map( A1 => DATA_IN(20), A2 => n18109, ZN => n14609);
   U16112 : NAND2_X1 port map( A1 => DATA_IN(21), A2 => n18109, ZN => n14608);
   U16113 : NAND2_X1 port map( A1 => DATA_IN(22), A2 => n18109, ZN => n14607);
   U16114 : NAND2_X1 port map( A1 => DATA_IN(23), A2 => n18109, ZN => n14606);
   U16115 : NAND2_X1 port map( A1 => DATA_IN(24), A2 => n18109, ZN => n14605);
   U16116 : NAND2_X1 port map( A1 => DATA_IN(25), A2 => n18109, ZN => n14604);
   U16117 : NAND2_X1 port map( A1 => DATA_IN(26), A2 => n18109, ZN => n14603);
   U16118 : NAND2_X1 port map( A1 => DATA_IN(27), A2 => n18109, ZN => n14602);
   U16119 : NAND2_X1 port map( A1 => DATA_IN(28), A2 => n18109, ZN => n14601);
   U16120 : NAND2_X1 port map( A1 => DATA_IN(29), A2 => n18109, ZN => n14600);
   U16121 : NAND2_X1 port map( A1 => DATA_IN(30), A2 => n18109, ZN => n14599);
   U16122 : NAND2_X1 port map( A1 => DATA_IN(31), A2 => n18109, ZN => n14597);
   U16123 : NAND2_X1 port map( A1 => RST, A2 => EN, ZN => n14632);
   U16124 : INV_X1 port map( A => ADDR_RD2(3), ZN => n13569);
   U16125 : INV_X1 port map( A => ADDR_RD1(3), ZN => n13565);
   U16126 : INV_X1 port map( A => ADDR_RD2(0), ZN => n13572);
   U16127 : INV_X1 port map( A => ADDR_RD1(0), ZN => n13568);
   U16128 : AND2_X1 port map( A1 => WR, A2 => EN, ZN => n14647);
   U16129 : INV_X1 port map( A => RST, ZN => n13559);
   U16130 : INV_X1 port map( A => ADDR_WR(2), ZN => n13562);
   U16131 : INV_X1 port map( A => ADDR_WR(0), ZN => n13564);
   U16132 : INV_X1 port map( A => ADDR_WR(1), ZN => n13563);
   U16133 : INV_X1 port map( A => ADDR_RD2(1), ZN => n13571);
   U16134 : INV_X1 port map( A => ADDR_RD1(1), ZN => n13567);
   U16135 : INV_X1 port map( A => ADDR_RD2(2), ZN => n13570);
   U16136 : INV_X1 port map( A => ADDR_RD1(2), ZN => n13566);
   U16137 : INV_X1 port map( A => ADDR_WR(4), ZN => n13560);
   U16138 : INV_X1 port map( A => ADDR_WR(3), ZN => n13561);
   U16139 : CLKBUF_X1 port map( A => n15328, Z => n17618);
   U16140 : CLKBUF_X1 port map( A => n14675, Z => n17720);

end SYN_beh;
