
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95;

architecture SYN_ARCH2 of ND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94;

architecture SYN_ARCH2 of ND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH2 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH2 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH2 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH2 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH2 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH2 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH2 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH2 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH2 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH2 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH2 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH2 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH2 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH2 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH2 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH2 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH2 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH2 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH2 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH2 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH2 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH2 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH2 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH2 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH2 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH2 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH2 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH2 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH2 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH2 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH2 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH2 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH2 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH2 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH2 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH2 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH2 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH2 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH2 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH2 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH2 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH2 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH2 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH2 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH2 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH2 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH2 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH2 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH2 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH2 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH2 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH2 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH2 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH2 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH2 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH2 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH2 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH2 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH2 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH2 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH2 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH2 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH2 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH2 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH2 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH2 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH2 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH2 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH2 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH2 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH2 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH2 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH2 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH2 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH2 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH2 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH2 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH2 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH2 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH2 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH2 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH2 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH2 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH2 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH2 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH2 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH2 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH2 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH2 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH2 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH2 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH2 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH2 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity MUX21_GENERIC_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_7;

architecture SYN_STRUCT of MUX21_GENERIC_NBIT4_7 is

   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal S_INV, NAND_OUT_A_3_port, NAND_OUT_A_2_port, NAND_OUT_A_1_port, 
      NAND_OUT_A_0_port, NAND_OUT_B_3_port, NAND_OUT_B_2_port, 
      NAND_OUT_B_1_port, NAND_OUT_B_0_port : std_logic;

begin
   
   INV : IV_7 port map( A => SEL, Y => S_INV);
   A_NAND_i_0 : ND2_84 port map( A => SEL, B => B(0), Y => NAND_OUT_A_0_port);
   B_NAND_i_0 : ND2_83 port map( A => S_INV, B => A(0), Y => NAND_OUT_B_0_port)
                           ;
   NAND_OUT_i_0 : ND2_82 port map( A => NAND_OUT_A_0_port, B => 
                           NAND_OUT_B_0_port, Y => Y(0));
   A_NAND_i_1 : ND2_81 port map( A => SEL, B => B(1), Y => NAND_OUT_A_1_port);
   B_NAND_i_1 : ND2_80 port map( A => S_INV, B => A(1), Y => NAND_OUT_B_1_port)
                           ;
   NAND_OUT_i_1 : ND2_79 port map( A => NAND_OUT_A_1_port, B => 
                           NAND_OUT_B_1_port, Y => Y(1));
   A_NAND_i_2 : ND2_78 port map( A => SEL, B => B(2), Y => NAND_OUT_A_2_port);
   B_NAND_i_2 : ND2_77 port map( A => S_INV, B => A(2), Y => NAND_OUT_B_2_port)
                           ;
   NAND_OUT_i_2 : ND2_76 port map( A => NAND_OUT_A_2_port, B => 
                           NAND_OUT_B_2_port, Y => Y(2));
   A_NAND_i_3 : ND2_75 port map( A => SEL, B => B(3), Y => NAND_OUT_A_3_port);
   B_NAND_i_3 : ND2_74 port map( A => S_INV, B => A(3), Y => NAND_OUT_B_3_port)
                           ;
   NAND_OUT_i_3 : ND2_73 port map( A => NAND_OUT_A_3_port, B => 
                           NAND_OUT_B_3_port, Y => Y(3));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity MUX21_GENERIC_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_6;

architecture SYN_STRUCT of MUX21_GENERIC_NBIT4_6 is

   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal S_INV, NAND_OUT_A_3_port, NAND_OUT_A_2_port, NAND_OUT_A_1_port, 
      NAND_OUT_A_0_port, NAND_OUT_B_3_port, NAND_OUT_B_2_port, 
      NAND_OUT_B_1_port, NAND_OUT_B_0_port : std_logic;

begin
   
   INV : IV_6 port map( A => SEL, Y => S_INV);
   A_NAND_i_0 : ND2_72 port map( A => SEL, B => B(0), Y => NAND_OUT_A_0_port);
   B_NAND_i_0 : ND2_71 port map( A => S_INV, B => A(0), Y => NAND_OUT_B_0_port)
                           ;
   NAND_OUT_i_0 : ND2_70 port map( A => NAND_OUT_A_0_port, B => 
                           NAND_OUT_B_0_port, Y => Y(0));
   A_NAND_i_1 : ND2_69 port map( A => SEL, B => B(1), Y => NAND_OUT_A_1_port);
   B_NAND_i_1 : ND2_68 port map( A => S_INV, B => A(1), Y => NAND_OUT_B_1_port)
                           ;
   NAND_OUT_i_1 : ND2_67 port map( A => NAND_OUT_A_1_port, B => 
                           NAND_OUT_B_1_port, Y => Y(1));
   A_NAND_i_2 : ND2_66 port map( A => SEL, B => B(2), Y => NAND_OUT_A_2_port);
   B_NAND_i_2 : ND2_65 port map( A => S_INV, B => A(2), Y => NAND_OUT_B_2_port)
                           ;
   NAND_OUT_i_2 : ND2_64 port map( A => NAND_OUT_A_2_port, B => 
                           NAND_OUT_B_2_port, Y => Y(2));
   A_NAND_i_3 : ND2_63 port map( A => SEL, B => B(3), Y => NAND_OUT_A_3_port);
   B_NAND_i_3 : ND2_62 port map( A => S_INV, B => A(3), Y => NAND_OUT_B_3_port)
                           ;
   NAND_OUT_i_3 : ND2_61 port map( A => NAND_OUT_A_3_port, B => 
                           NAND_OUT_B_3_port, Y => Y(3));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity MUX21_GENERIC_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_5;

architecture SYN_STRUCT of MUX21_GENERIC_NBIT4_5 is

   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal S_INV, NAND_OUT_A_3_port, NAND_OUT_A_2_port, NAND_OUT_A_1_port, 
      NAND_OUT_A_0_port, NAND_OUT_B_3_port, NAND_OUT_B_2_port, 
      NAND_OUT_B_1_port, NAND_OUT_B_0_port : std_logic;

begin
   
   INV : IV_5 port map( A => SEL, Y => S_INV);
   A_NAND_i_0 : ND2_60 port map( A => SEL, B => B(0), Y => NAND_OUT_A_0_port);
   B_NAND_i_0 : ND2_59 port map( A => S_INV, B => A(0), Y => NAND_OUT_B_0_port)
                           ;
   NAND_OUT_i_0 : ND2_58 port map( A => NAND_OUT_A_0_port, B => 
                           NAND_OUT_B_0_port, Y => Y(0));
   A_NAND_i_1 : ND2_57 port map( A => SEL, B => B(1), Y => NAND_OUT_A_1_port);
   B_NAND_i_1 : ND2_56 port map( A => S_INV, B => A(1), Y => NAND_OUT_B_1_port)
                           ;
   NAND_OUT_i_1 : ND2_55 port map( A => NAND_OUT_A_1_port, B => 
                           NAND_OUT_B_1_port, Y => Y(1));
   A_NAND_i_2 : ND2_54 port map( A => SEL, B => B(2), Y => NAND_OUT_A_2_port);
   B_NAND_i_2 : ND2_53 port map( A => S_INV, B => A(2), Y => NAND_OUT_B_2_port)
                           ;
   NAND_OUT_i_2 : ND2_52 port map( A => NAND_OUT_A_2_port, B => 
                           NAND_OUT_B_2_port, Y => Y(2));
   A_NAND_i_3 : ND2_51 port map( A => SEL, B => B(3), Y => NAND_OUT_A_3_port);
   B_NAND_i_3 : ND2_50 port map( A => S_INV, B => A(3), Y => NAND_OUT_B_3_port)
                           ;
   NAND_OUT_i_3 : ND2_49 port map( A => NAND_OUT_A_3_port, B => 
                           NAND_OUT_B_3_port, Y => Y(3));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity MUX21_GENERIC_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_4;

architecture SYN_STRUCT of MUX21_GENERIC_NBIT4_4 is

   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal S_INV, NAND_OUT_A_3_port, NAND_OUT_A_2_port, NAND_OUT_A_1_port, 
      NAND_OUT_A_0_port, NAND_OUT_B_3_port, NAND_OUT_B_2_port, 
      NAND_OUT_B_1_port, NAND_OUT_B_0_port : std_logic;

begin
   
   INV : IV_4 port map( A => SEL, Y => S_INV);
   A_NAND_i_0 : ND2_48 port map( A => SEL, B => B(0), Y => NAND_OUT_A_0_port);
   B_NAND_i_0 : ND2_47 port map( A => S_INV, B => A(0), Y => NAND_OUT_B_0_port)
                           ;
   NAND_OUT_i_0 : ND2_46 port map( A => NAND_OUT_A_0_port, B => 
                           NAND_OUT_B_0_port, Y => Y(0));
   A_NAND_i_1 : ND2_45 port map( A => SEL, B => B(1), Y => NAND_OUT_A_1_port);
   B_NAND_i_1 : ND2_44 port map( A => S_INV, B => A(1), Y => NAND_OUT_B_1_port)
                           ;
   NAND_OUT_i_1 : ND2_43 port map( A => NAND_OUT_A_1_port, B => 
                           NAND_OUT_B_1_port, Y => Y(1));
   A_NAND_i_2 : ND2_42 port map( A => SEL, B => B(2), Y => NAND_OUT_A_2_port);
   B_NAND_i_2 : ND2_41 port map( A => S_INV, B => A(2), Y => NAND_OUT_B_2_port)
                           ;
   NAND_OUT_i_2 : ND2_40 port map( A => NAND_OUT_A_2_port, B => 
                           NAND_OUT_B_2_port, Y => Y(2));
   A_NAND_i_3 : ND2_39 port map( A => SEL, B => B(3), Y => NAND_OUT_A_3_port);
   B_NAND_i_3 : ND2_38 port map( A => S_INV, B => A(3), Y => NAND_OUT_B_3_port)
                           ;
   NAND_OUT_i_3 : ND2_37 port map( A => NAND_OUT_A_3_port, B => 
                           NAND_OUT_B_3_port, Y => Y(3));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity MUX21_GENERIC_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_3;

architecture SYN_STRUCT of MUX21_GENERIC_NBIT4_3 is

   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal S_INV, NAND_OUT_A_3_port, NAND_OUT_A_2_port, NAND_OUT_A_1_port, 
      NAND_OUT_A_0_port, NAND_OUT_B_3_port, NAND_OUT_B_2_port, 
      NAND_OUT_B_1_port, NAND_OUT_B_0_port : std_logic;

begin
   
   INV : IV_3 port map( A => SEL, Y => S_INV);
   A_NAND_i_0 : ND2_36 port map( A => SEL, B => B(0), Y => NAND_OUT_A_0_port);
   B_NAND_i_0 : ND2_35 port map( A => S_INV, B => A(0), Y => NAND_OUT_B_0_port)
                           ;
   NAND_OUT_i_0 : ND2_34 port map( A => NAND_OUT_A_0_port, B => 
                           NAND_OUT_B_0_port, Y => Y(0));
   A_NAND_i_1 : ND2_33 port map( A => SEL, B => B(1), Y => NAND_OUT_A_1_port);
   B_NAND_i_1 : ND2_32 port map( A => S_INV, B => A(1), Y => NAND_OUT_B_1_port)
                           ;
   NAND_OUT_i_1 : ND2_31 port map( A => NAND_OUT_A_1_port, B => 
                           NAND_OUT_B_1_port, Y => Y(1));
   A_NAND_i_2 : ND2_30 port map( A => SEL, B => B(2), Y => NAND_OUT_A_2_port);
   B_NAND_i_2 : ND2_29 port map( A => S_INV, B => A(2), Y => NAND_OUT_B_2_port)
                           ;
   NAND_OUT_i_2 : ND2_28 port map( A => NAND_OUT_A_2_port, B => 
                           NAND_OUT_B_2_port, Y => Y(2));
   A_NAND_i_3 : ND2_27 port map( A => SEL, B => B(3), Y => NAND_OUT_A_3_port);
   B_NAND_i_3 : ND2_26 port map( A => S_INV, B => A(3), Y => NAND_OUT_B_3_port)
                           ;
   NAND_OUT_i_3 : ND2_25 port map( A => NAND_OUT_A_3_port, B => 
                           NAND_OUT_B_3_port, Y => Y(3));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity MUX21_GENERIC_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_2;

architecture SYN_STRUCT of MUX21_GENERIC_NBIT4_2 is

   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal S_INV, NAND_OUT_A_3_port, NAND_OUT_A_2_port, NAND_OUT_A_1_port, 
      NAND_OUT_A_0_port, NAND_OUT_B_3_port, NAND_OUT_B_2_port, 
      NAND_OUT_B_1_port, NAND_OUT_B_0_port : std_logic;

begin
   
   INV : IV_2 port map( A => SEL, Y => S_INV);
   A_NAND_i_0 : ND2_24 port map( A => SEL, B => B(0), Y => NAND_OUT_A_0_port);
   B_NAND_i_0 : ND2_23 port map( A => S_INV, B => A(0), Y => NAND_OUT_B_0_port)
                           ;
   NAND_OUT_i_0 : ND2_22 port map( A => NAND_OUT_A_0_port, B => 
                           NAND_OUT_B_0_port, Y => Y(0));
   A_NAND_i_1 : ND2_21 port map( A => SEL, B => B(1), Y => NAND_OUT_A_1_port);
   B_NAND_i_1 : ND2_20 port map( A => S_INV, B => A(1), Y => NAND_OUT_B_1_port)
                           ;
   NAND_OUT_i_1 : ND2_19 port map( A => NAND_OUT_A_1_port, B => 
                           NAND_OUT_B_1_port, Y => Y(1));
   A_NAND_i_2 : ND2_18 port map( A => SEL, B => B(2), Y => NAND_OUT_A_2_port);
   B_NAND_i_2 : ND2_17 port map( A => S_INV, B => A(2), Y => NAND_OUT_B_2_port)
                           ;
   NAND_OUT_i_2 : ND2_16 port map( A => NAND_OUT_A_2_port, B => 
                           NAND_OUT_B_2_port, Y => Y(2));
   A_NAND_i_3 : ND2_15 port map( A => SEL, B => B(3), Y => NAND_OUT_A_3_port);
   B_NAND_i_3 : ND2_14 port map( A => S_INV, B => A(3), Y => NAND_OUT_B_3_port)
                           ;
   NAND_OUT_i_3 : ND2_13 port map( A => NAND_OUT_A_3_port, B => 
                           NAND_OUT_B_3_port, Y => Y(3));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity MUX21_GENERIC_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_1;

architecture SYN_STRUCT of MUX21_GENERIC_NBIT4_1 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal S_INV, NAND_OUT_A_3_port, NAND_OUT_A_2_port, NAND_OUT_A_1_port, 
      NAND_OUT_A_0_port, NAND_OUT_B_3_port, NAND_OUT_B_2_port, 
      NAND_OUT_B_1_port, NAND_OUT_B_0_port : std_logic;

begin
   
   INV : IV_1 port map( A => SEL, Y => S_INV);
   A_NAND_i_0 : ND2_12 port map( A => SEL, B => B(0), Y => NAND_OUT_A_0_port);
   B_NAND_i_0 : ND2_11 port map( A => S_INV, B => A(0), Y => NAND_OUT_B_0_port)
                           ;
   NAND_OUT_i_0 : ND2_10 port map( A => NAND_OUT_A_0_port, B => 
                           NAND_OUT_B_0_port, Y => Y(0));
   A_NAND_i_1 : ND2_9 port map( A => SEL, B => B(1), Y => NAND_OUT_A_1_port);
   B_NAND_i_1 : ND2_8 port map( A => S_INV, B => A(1), Y => NAND_OUT_B_1_port);
   NAND_OUT_i_1 : ND2_7 port map( A => NAND_OUT_A_1_port, B => 
                           NAND_OUT_B_1_port, Y => Y(1));
   A_NAND_i_2 : ND2_6 port map( A => SEL, B => B(2), Y => NAND_OUT_A_2_port);
   B_NAND_i_2 : ND2_5 port map( A => S_INV, B => A(2), Y => NAND_OUT_B_2_port);
   NAND_OUT_i_2 : ND2_4 port map( A => NAND_OUT_A_2_port, B => 
                           NAND_OUT_B_2_port, Y => Y(2));
   A_NAND_i_3 : ND2_3 port map( A => SEL, B => B(3), Y => NAND_OUT_A_3_port);
   B_NAND_i_3 : ND2_2 port map( A => S_INV, B => A(3), Y => NAND_OUT_B_3_port);
   NAND_OUT_i_3 : ND2_1 port map( A => NAND_OUT_A_3_port, B => 
                           NAND_OUT_B_3_port, Y => Y(3));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_15;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_15 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_14;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_14 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_13;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_13 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_12;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_12 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_11;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_11 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_10;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_10 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_9;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_9 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_8;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_8 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_7;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_7 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_6;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_6 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_5;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_5 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_4;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_4 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_3;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_3 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_2;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_2 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_1;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_1 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CARRY_SELECT_BLOCK_GENERIC_NBIT4_7 is

   port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
         out std_logic_vector (3 downto 0));

end CARRY_SELECT_BLOCK_GENERIC_NBIT4_7;

architecture SYN_STRUCTURAL of CARRY_SELECT_BLOCK_GENERIC_NBIT4_7 is

   component MUX21_GENERIC_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GENERIC_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1000, n_1001 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GENERIC_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1000);
   RCA1 : RCA_GENERIC_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1001);
   MUX : MUX21_GENERIC_NBIT4_7 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => C_IN, Y(3) => S(3), Y(2) 
                           => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CARRY_SELECT_BLOCK_GENERIC_NBIT4_6 is

   port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
         out std_logic_vector (3 downto 0));

end CARRY_SELECT_BLOCK_GENERIC_NBIT4_6;

architecture SYN_STRUCTURAL of CARRY_SELECT_BLOCK_GENERIC_NBIT4_6 is

   component MUX21_GENERIC_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GENERIC_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1002, n_1003 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GENERIC_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1002);
   RCA1 : RCA_GENERIC_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1003);
   MUX : MUX21_GENERIC_NBIT4_6 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => C_IN, Y(3) => S(3), Y(2) 
                           => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CARRY_SELECT_BLOCK_GENERIC_NBIT4_5 is

   port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
         out std_logic_vector (3 downto 0));

end CARRY_SELECT_BLOCK_GENERIC_NBIT4_5;

architecture SYN_STRUCTURAL of CARRY_SELECT_BLOCK_GENERIC_NBIT4_5 is

   component MUX21_GENERIC_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GENERIC_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1004, n_1005 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GENERIC_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1004);
   RCA1 : RCA_GENERIC_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1005);
   MUX : MUX21_GENERIC_NBIT4_5 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => C_IN, Y(3) => S(3), Y(2) 
                           => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CARRY_SELECT_BLOCK_GENERIC_NBIT4_4 is

   port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
         out std_logic_vector (3 downto 0));

end CARRY_SELECT_BLOCK_GENERIC_NBIT4_4;

architecture SYN_STRUCTURAL of CARRY_SELECT_BLOCK_GENERIC_NBIT4_4 is

   component MUX21_GENERIC_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GENERIC_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1006, n_1007 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GENERIC_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1006);
   RCA1 : RCA_GENERIC_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1007);
   MUX : MUX21_GENERIC_NBIT4_4 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => C_IN, Y(3) => S(3), Y(2) 
                           => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CARRY_SELECT_BLOCK_GENERIC_NBIT4_3 is

   port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
         out std_logic_vector (3 downto 0));

end CARRY_SELECT_BLOCK_GENERIC_NBIT4_3;

architecture SYN_STRUCTURAL of CARRY_SELECT_BLOCK_GENERIC_NBIT4_3 is

   component MUX21_GENERIC_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GENERIC_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1008, n_1009 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GENERIC_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1008);
   RCA1 : RCA_GENERIC_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1009);
   MUX : MUX21_GENERIC_NBIT4_3 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => C_IN, Y(3) => S(3), Y(2) 
                           => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CARRY_SELECT_BLOCK_GENERIC_NBIT4_2 is

   port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
         out std_logic_vector (3 downto 0));

end CARRY_SELECT_BLOCK_GENERIC_NBIT4_2;

architecture SYN_STRUCTURAL of CARRY_SELECT_BLOCK_GENERIC_NBIT4_2 is

   component MUX21_GENERIC_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GENERIC_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1010, n_1011 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GENERIC_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1010);
   RCA1 : RCA_GENERIC_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1011);
   MUX : MUX21_GENERIC_NBIT4_2 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => C_IN, Y(3) => S(3), Y(2) 
                           => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CARRY_SELECT_BLOCK_GENERIC_NBIT4_1 is

   port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
         out std_logic_vector (3 downto 0));

end CARRY_SELECT_BLOCK_GENERIC_NBIT4_1;

architecture SYN_STRUCTURAL of CARRY_SELECT_BLOCK_GENERIC_NBIT4_1 is

   component MUX21_GENERIC_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GENERIC_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1012, n_1013 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GENERIC_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1012);
   RCA1 : RCA_GENERIC_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1013);
   MUX : MUX21_GENERIC_NBIT4_1 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => C_IN, Y(3) => S(3), Y(2) 
                           => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_27 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_27;

architecture SYN_beh of PG_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_26 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_26;

architecture SYN_beh of PG_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_25 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_25;

architecture SYN_beh of PG_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_24 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_24;

architecture SYN_beh of PG_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_23 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_23;

architecture SYN_beh of PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_22 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_22;

architecture SYN_beh of PG_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_21 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_21;

architecture SYN_beh of PG_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_20 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_20;

architecture SYN_beh of PG_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_19 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_19;

architecture SYN_beh of PG_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_18 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_18;

architecture SYN_beh of PG_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_17 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_17;

architecture SYN_beh of PG_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_16 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_16;

architecture SYN_beh of PG_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_15 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_15;

architecture SYN_beh of PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_14 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_14;

architecture SYN_beh of PG_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_13 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_13;

architecture SYN_beh of PG_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_12 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_12;

architecture SYN_beh of PG_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_11 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_11;

architecture SYN_beh of PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_10 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_10;

architecture SYN_beh of PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_9 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_9;

architecture SYN_beh of PG_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_8 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_8;

architecture SYN_beh of PG_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_7 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_7;

architecture SYN_beh of PG_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_6 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_6;

architecture SYN_beh of PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_5 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_5;

architecture SYN_beh of PG_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_4 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_4;

architecture SYN_beh of PG_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_3 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_3;

architecture SYN_beh of PG_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_2 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_2;

architecture SYN_beh of PG_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_1 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_1;

architecture SYN_beh of PG_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_9 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_9;

architecture SYN_beh of G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_8 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_8;

architecture SYN_beh of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_7 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_7;

architecture SYN_beh of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_6 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_6;

architecture SYN_beh of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_5 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_5;

architecture SYN_beh of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_4 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_4;

architecture SYN_beh of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_3 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_3;

architecture SYN_beh of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_2 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_2;

architecture SYN_beh of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_1 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_1;

architecture SYN_beh of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_31 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_31;

architecture SYN_beh of pgb_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_30 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_30;

architecture SYN_beh of pgb_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_29 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_29;

architecture SYN_beh of pgb_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_28 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_28;

architecture SYN_beh of pgb_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_27 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_27;

architecture SYN_beh of pgb_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_26 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_26;

architecture SYN_beh of pgb_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_25 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_25;

architecture SYN_beh of pgb_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_24 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_24;

architecture SYN_beh of pgb_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_23 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_23;

architecture SYN_beh of pgb_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_22 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_22;

architecture SYN_beh of pgb_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_21 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_21;

architecture SYN_beh of pgb_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_20 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_20;

architecture SYN_beh of pgb_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_19 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_19;

architecture SYN_beh of pgb_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_18 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_18;

architecture SYN_beh of pgb_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_17 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_17;

architecture SYN_beh of pgb_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_16 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_16;

architecture SYN_beh of pgb_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_15 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_15;

architecture SYN_beh of pgb_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_14 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_14;

architecture SYN_beh of pgb_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_13 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_13;

architecture SYN_beh of pgb_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_12 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_12;

architecture SYN_beh of pgb_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_11 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_11;

architecture SYN_beh of pgb_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_10 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_10;

architecture SYN_beh of pgb_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_9 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_9;

architecture SYN_beh of pgb_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_8 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_8;

architecture SYN_beh of pgb_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_7 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_7;

architecture SYN_beh of pgb_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_6 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_6;

architecture SYN_beh of pgb_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_5 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_5;

architecture SYN_beh of pgb_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_4 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_4;

architecture SYN_beh of pgb_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_3 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_3;

architecture SYN_beh of pgb_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_2 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_2;

architecture SYN_beh of pgb_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_1 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_1;

architecture SYN_beh of pgb_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity ND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0;

architecture SYN_ARCH2 of ND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity MUX21_GENERIC_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_0;

architecture SYN_STRUCT of MUX21_GENERIC_NBIT4_0 is

   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal S_INV, NAND_OUT_A_3_port, NAND_OUT_A_2_port, NAND_OUT_A_1_port, 
      NAND_OUT_A_0_port, NAND_OUT_B_3_port, NAND_OUT_B_2_port, 
      NAND_OUT_B_1_port, NAND_OUT_B_0_port : std_logic;

begin
   
   INV : IV_0 port map( A => SEL, Y => S_INV);
   A_NAND_i_0 : ND2_0 port map( A => SEL, B => B(0), Y => NAND_OUT_A_0_port);
   B_NAND_i_0 : ND2_95 port map( A => S_INV, B => A(0), Y => NAND_OUT_B_0_port)
                           ;
   NAND_OUT_i_0 : ND2_94 port map( A => NAND_OUT_A_0_port, B => 
                           NAND_OUT_B_0_port, Y => Y(0));
   A_NAND_i_1 : ND2_93 port map( A => SEL, B => B(1), Y => NAND_OUT_A_1_port);
   B_NAND_i_1 : ND2_92 port map( A => S_INV, B => A(1), Y => NAND_OUT_B_1_port)
                           ;
   NAND_OUT_i_1 : ND2_91 port map( A => NAND_OUT_A_1_port, B => 
                           NAND_OUT_B_1_port, Y => Y(1));
   A_NAND_i_2 : ND2_90 port map( A => SEL, B => B(2), Y => NAND_OUT_A_2_port);
   B_NAND_i_2 : ND2_89 port map( A => S_INV, B => A(2), Y => NAND_OUT_B_2_port)
                           ;
   NAND_OUT_i_2 : ND2_88 port map( A => NAND_OUT_A_2_port, B => 
                           NAND_OUT_B_2_port, Y => Y(2));
   A_NAND_i_3 : ND2_87 port map( A => SEL, B => B(3), Y => NAND_OUT_A_3_port);
   B_NAND_i_3 : ND2_86 port map( A => S_INV, B => A(3), Y => NAND_OUT_B_3_port)
                           ;
   NAND_OUT_i_3 : ND2_85 port map( A => NAND_OUT_A_3_port, B => 
                           NAND_OUT_B_3_port, Y => Y(3));

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity RCA_GENERIC_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GENERIC_NBIT4_0;

architecture SYN_BEHAVIORAL of RCA_GENERIC_NBIT4_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_55_2_carry_1_port, add_1_root_add_55_2_carry_2_port, 
      add_1_root_add_55_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_55_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_55_2_carry_1_port, S => S(0));
   add_1_root_add_55_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_55_2_carry_1_port, CO => 
                           add_1_root_add_55_2_carry_2_port, S => S(1));
   add_1_root_add_55_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_55_2_carry_2_port, CO => 
                           add_1_root_add_55_2_carry_3_port, S => S(2));
   add_1_root_add_55_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_55_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CARRY_SELECT_BLOCK_GENERIC_NBIT4_0 is

   port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
         out std_logic_vector (3 downto 0));

end CARRY_SELECT_BLOCK_GENERIC_NBIT4_0;

architecture SYN_STRUCTURAL of CARRY_SELECT_BLOCK_GENERIC_NBIT4_0 is

   component MUX21_GENERIC_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GENERIC_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GENERIC_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1014, n_1015 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GENERIC_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1014);
   RCA1 : RCA_GENERIC_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1015);
   MUX : MUX21_GENERIC_NBIT4_0 port map( A(3) => S0_3_port, A(2) => S0_2_port, 
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => C_IN, Y(3) => S(3), Y(2) 
                           => S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity PG_0 is

   port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);

end PG_0;

architecture SYN_beh of PG_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);
   U3 : AND2_X1 port map( A1 => Pdkj, A2 => Pik, ZN => Pij);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity G_0 is

   port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);

end G_0;

architecture SYN_beh of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Gij);
   U2 : AOI21_X1 port map( B1 => Pik, B2 => Gdkj, A => Gik, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity pgb_0 is

   port( ai, bi : in std_logic;  p, g : out std_logic);

end pgb_0;

architecture SYN_beh of pgb_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => bi, B => ai, Z => p);
   U2 : AND2_X1 port map( A1 => bi, A2 => ai, ZN => g);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity SUM_GENERATOR_GENERIC_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_GENERIC_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_STRUCTURAL of SUM_GENERATOR_GENERIC_NBIT_PER_BLOCK4_NBLOCKS8 
   is

   component CARRY_SELECT_BLOCK_GENERIC_NBIT4_1
      port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S :
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SELECT_BLOCK_GENERIC_NBIT4_2
      port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S :
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SELECT_BLOCK_GENERIC_NBIT4_3
      port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S :
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SELECT_BLOCK_GENERIC_NBIT4_4
      port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S :
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SELECT_BLOCK_GENERIC_NBIT4_5
      port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S :
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SELECT_BLOCK_GENERIC_NBIT4_6
      port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S :
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SELECT_BLOCK_GENERIC_NBIT4_7
      port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S :
            out std_logic_vector (3 downto 0));
   end component;
   
   component CARRY_SELECT_BLOCK_GENERIC_NBIT4_0
      port( C_IN : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S :
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CARRYSELBLOCK_i_1 : CARRY_SELECT_BLOCK_GENERIC_NBIT4_0 port map( C_IN => 
                           Ci(0), A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));
   CARRYSELBLOCK_i_2 : CARRY_SELECT_BLOCK_GENERIC_NBIT4_7 port map( C_IN => 
                           Ci(1), A(3) => A(7), A(2) => A(6), A(1) => A(5), 
                           A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1) => 
                           B(5), B(0) => B(4), S(3) => S(7), S(2) => S(6), S(1)
                           => S(5), S(0) => S(4));
   CARRYSELBLOCK_i_3 : CARRY_SELECT_BLOCK_GENERIC_NBIT4_6 port map( C_IN => 
                           Ci(2), A(3) => A(11), A(2) => A(10), A(1) => A(9), 
                           A(0) => A(8), B(3) => B(11), B(2) => B(10), B(1) => 
                           B(9), B(0) => B(8), S(3) => S(11), S(2) => S(10), 
                           S(1) => S(9), S(0) => S(8));
   CARRYSELBLOCK_i_4 : CARRY_SELECT_BLOCK_GENERIC_NBIT4_5 port map( C_IN => 
                           Ci(3), A(3) => A(15), A(2) => A(14), A(1) => A(13), 
                           A(0) => A(12), B(3) => B(15), B(2) => B(14), B(1) =>
                           B(13), B(0) => B(12), S(3) => S(15), S(2) => S(14), 
                           S(1) => S(13), S(0) => S(12));
   CARRYSELBLOCK_i_5 : CARRY_SELECT_BLOCK_GENERIC_NBIT4_4 port map( C_IN => 
                           Ci(4), A(3) => A(19), A(2) => A(18), A(1) => A(17), 
                           A(0) => A(16), B(3) => B(19), B(2) => B(18), B(1) =>
                           B(17), B(0) => B(16), S(3) => S(19), S(2) => S(18), 
                           S(1) => S(17), S(0) => S(16));
   CARRYSELBLOCK_i_6 : CARRY_SELECT_BLOCK_GENERIC_NBIT4_3 port map( C_IN => 
                           Ci(5), A(3) => A(23), A(2) => A(22), A(1) => A(21), 
                           A(0) => A(20), B(3) => B(23), B(2) => B(22), B(1) =>
                           B(21), B(0) => B(20), S(3) => S(23), S(2) => S(22), 
                           S(1) => S(21), S(0) => S(20));
   CARRYSELBLOCK_i_7 : CARRY_SELECT_BLOCK_GENERIC_NBIT4_2 port map( C_IN => 
                           Ci(6), A(3) => A(27), A(2) => A(26), A(1) => A(25), 
                           A(0) => A(24), B(3) => B(27), B(2) => B(26), B(1) =>
                           B(25), B(0) => B(24), S(3) => S(27), S(2) => S(26), 
                           S(1) => S(25), S(0) => S(24));
   CARRYSELBLOCK_i_8 : CARRY_SELECT_BLOCK_GENERIC_NBIT4_1 port map( C_IN => 
                           Ci(7), A(3) => A(31), A(2) => A(30), A(1) => A(29), 
                           A(0) => A(28), B(3) => B(31), B(2) => B(30), B(1) =>
                           B(29), B(0) => B(28), S(3) => S(31), S(2) => S(30), 
                           S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity CLA_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CLA_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_structural_generic of CLA_NBIT32_NBIT_PER_BLOCK4 is

   component G_1
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_1
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_2
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_3
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_4
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_5
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component G_2
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_6
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_7
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_8
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_9
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component G_3
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_10
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_11
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_12
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_13
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component G_4
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_14
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_15
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_16
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_17
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component G_5
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_18
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_19
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_20
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_21
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component G_6
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_22
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_23
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_24
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component G_7
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_25
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_26
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component PG_27
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component G_8
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component G_9
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component PG_0
      port( Pik, Pdkj, Gik, Gdkj : in std_logic;  Pij, Gij : out std_logic);
   end component;
   
   component pgb_1
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_2
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_3
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_4
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_5
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_6
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_7
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_8
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_9
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_10
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_11
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_12
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_13
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_14
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_15
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_16
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_17
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_18
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_19
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_20
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_21
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_22
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_23
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_24
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_25
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_26
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_27
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_28
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_29
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_30
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component pgb_31
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   component G_0
      port( Pik, Gik, Gdkj : in std_logic;  Gij : out std_logic);
   end component;
   
   component pgb_0
      port( ai, bi : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port, g_pgb00_G00, p_pgb00_G00, gi_matrix_0_0_port, 
      gi_matrix_0_1_port, gi_matrix_0_2_port, gi_matrix_0_3_port, 
      gi_matrix_0_4_port, gi_matrix_0_5_port, gi_matrix_0_6_port, 
      gi_matrix_0_7_port, gi_matrix_0_8_port, gi_matrix_0_9_port, 
      gi_matrix_0_10_port, gi_matrix_0_11_port, gi_matrix_0_12_port, 
      gi_matrix_0_13_port, gi_matrix_0_14_port, gi_matrix_0_15_port, 
      gi_matrix_0_16_port, gi_matrix_0_17_port, gi_matrix_0_18_port, 
      gi_matrix_0_19_port, gi_matrix_0_20_port, gi_matrix_0_21_port, 
      gi_matrix_0_22_port, gi_matrix_0_23_port, gi_matrix_0_24_port, 
      gi_matrix_0_25_port, gi_matrix_0_26_port, gi_matrix_0_27_port, 
      gi_matrix_0_28_port, gi_matrix_0_29_port, gi_matrix_0_30_port, 
      gi_matrix_0_31_port, gi_matrix_1_1_port, gi_matrix_1_3_port, 
      gi_matrix_1_5_port, gi_matrix_1_7_port, gi_matrix_1_9_port, 
      gi_matrix_1_11_port, gi_matrix_1_13_port, gi_matrix_1_15_port, 
      gi_matrix_1_17_port, gi_matrix_1_19_port, gi_matrix_1_21_port, 
      gi_matrix_1_23_port, gi_matrix_1_25_port, gi_matrix_1_27_port, 
      gi_matrix_1_29_port, gi_matrix_1_31_port, gi_matrix_2_7_port, 
      gi_matrix_2_11_port, gi_matrix_2_15_port, gi_matrix_2_19_port, 
      gi_matrix_2_23_port, gi_matrix_2_27_port, gi_matrix_2_31_port, 
      gi_matrix_3_15_port, gi_matrix_3_19_port, gi_matrix_3_23_port, 
      gi_matrix_3_27_port, gi_matrix_3_31_port, gi_matrix_4_31_port, 
      pi_matrix_0_1_port, pi_matrix_0_2_port, pi_matrix_0_3_port, 
      pi_matrix_0_4_port, pi_matrix_0_5_port, pi_matrix_0_6_port, 
      pi_matrix_0_7_port, pi_matrix_0_8_port, pi_matrix_0_9_port, 
      pi_matrix_0_10_port, pi_matrix_0_11_port, pi_matrix_0_12_port, 
      pi_matrix_0_13_port, pi_matrix_0_14_port, pi_matrix_0_15_port, 
      pi_matrix_0_16_port, pi_matrix_0_17_port, pi_matrix_0_18_port, 
      pi_matrix_0_19_port, pi_matrix_0_20_port, pi_matrix_0_21_port, 
      pi_matrix_0_22_port, pi_matrix_0_23_port, pi_matrix_0_24_port, 
      pi_matrix_0_25_port, pi_matrix_0_26_port, pi_matrix_0_27_port, 
      pi_matrix_0_28_port, pi_matrix_0_29_port, pi_matrix_0_30_port, 
      pi_matrix_0_31_port, pi_matrix_1_3_port, pi_matrix_1_5_port, 
      pi_matrix_1_7_port, pi_matrix_1_9_port, pi_matrix_1_11_port, 
      pi_matrix_1_13_port, pi_matrix_1_15_port, pi_matrix_1_17_port, 
      pi_matrix_1_19_port, pi_matrix_1_21_port, pi_matrix_1_23_port, 
      pi_matrix_1_25_port, pi_matrix_1_27_port, pi_matrix_1_29_port, 
      pi_matrix_1_31_port, pi_matrix_2_7_port, pi_matrix_2_11_port, 
      pi_matrix_2_15_port, pi_matrix_2_19_port, pi_matrix_2_23_port, 
      pi_matrix_2_27_port, pi_matrix_2_31_port, pi_matrix_3_15_port, 
      pi_matrix_3_19_port, pi_matrix_3_23_port, pi_matrix_3_27_port, 
      pi_matrix_3_31_port, pi_matrix_4_31_port : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   PG_0_0 : pgb_0 port map( ai => A(0), bi => B(0), p => p_pgb00_G00, g => 
                           g_pgb00_G00);
   G_0_0 : G_0 port map( Pik => p_pgb00_G00, Gik => g_pgb00_G00, Gdkj => Cin, 
                           Gij => gi_matrix_0_0_port);
   PG_i_1 : pgb_31 port map( ai => A(1), bi => B(1), p => pi_matrix_0_1_port, g
                           => gi_matrix_0_1_port);
   PG_i_2 : pgb_30 port map( ai => A(2), bi => B(2), p => pi_matrix_0_2_port, g
                           => gi_matrix_0_2_port);
   PG_i_3 : pgb_29 port map( ai => A(3), bi => B(3), p => pi_matrix_0_3_port, g
                           => gi_matrix_0_3_port);
   PG_i_4 : pgb_28 port map( ai => A(4), bi => B(4), p => pi_matrix_0_4_port, g
                           => gi_matrix_0_4_port);
   PG_i_5 : pgb_27 port map( ai => A(5), bi => B(5), p => pi_matrix_0_5_port, g
                           => gi_matrix_0_5_port);
   PG_i_6 : pgb_26 port map( ai => A(6), bi => B(6), p => pi_matrix_0_6_port, g
                           => gi_matrix_0_6_port);
   PG_i_7 : pgb_25 port map( ai => A(7), bi => B(7), p => pi_matrix_0_7_port, g
                           => gi_matrix_0_7_port);
   PG_i_8 : pgb_24 port map( ai => A(8), bi => B(8), p => pi_matrix_0_8_port, g
                           => gi_matrix_0_8_port);
   PG_i_9 : pgb_23 port map( ai => A(9), bi => B(9), p => pi_matrix_0_9_port, g
                           => gi_matrix_0_9_port);
   PG_i_10 : pgb_22 port map( ai => A(10), bi => B(10), p => 
                           pi_matrix_0_10_port, g => gi_matrix_0_10_port);
   PG_i_11 : pgb_21 port map( ai => A(11), bi => B(11), p => 
                           pi_matrix_0_11_port, g => gi_matrix_0_11_port);
   PG_i_12 : pgb_20 port map( ai => A(12), bi => B(12), p => 
                           pi_matrix_0_12_port, g => gi_matrix_0_12_port);
   PG_i_13 : pgb_19 port map( ai => A(13), bi => B(13), p => 
                           pi_matrix_0_13_port, g => gi_matrix_0_13_port);
   PG_i_14 : pgb_18 port map( ai => A(14), bi => B(14), p => 
                           pi_matrix_0_14_port, g => gi_matrix_0_14_port);
   PG_i_15 : pgb_17 port map( ai => A(15), bi => B(15), p => 
                           pi_matrix_0_15_port, g => gi_matrix_0_15_port);
   PG_i_16 : pgb_16 port map( ai => A(16), bi => B(16), p => 
                           pi_matrix_0_16_port, g => gi_matrix_0_16_port);
   PG_i_17 : pgb_15 port map( ai => A(17), bi => B(17), p => 
                           pi_matrix_0_17_port, g => gi_matrix_0_17_port);
   PG_i_18 : pgb_14 port map( ai => A(18), bi => B(18), p => 
                           pi_matrix_0_18_port, g => gi_matrix_0_18_port);
   PG_i_19 : pgb_13 port map( ai => A(19), bi => B(19), p => 
                           pi_matrix_0_19_port, g => gi_matrix_0_19_port);
   PG_i_20 : pgb_12 port map( ai => A(20), bi => B(20), p => 
                           pi_matrix_0_20_port, g => gi_matrix_0_20_port);
   PG_i_21 : pgb_11 port map( ai => A(21), bi => B(21), p => 
                           pi_matrix_0_21_port, g => gi_matrix_0_21_port);
   PG_i_22 : pgb_10 port map( ai => A(22), bi => B(22), p => 
                           pi_matrix_0_22_port, g => gi_matrix_0_22_port);
   PG_i_23 : pgb_9 port map( ai => A(23), bi => B(23), p => pi_matrix_0_23_port
                           , g => gi_matrix_0_23_port);
   PG_i_24 : pgb_8 port map( ai => A(24), bi => B(24), p => pi_matrix_0_24_port
                           , g => gi_matrix_0_24_port);
   PG_i_25 : pgb_7 port map( ai => A(25), bi => B(25), p => pi_matrix_0_25_port
                           , g => gi_matrix_0_25_port);
   PG_i_26 : pgb_6 port map( ai => A(26), bi => B(26), p => pi_matrix_0_26_port
                           , g => gi_matrix_0_26_port);
   PG_i_27 : pgb_5 port map( ai => A(27), bi => B(27), p => pi_matrix_0_27_port
                           , g => gi_matrix_0_27_port);
   PG_i_28 : pgb_4 port map( ai => A(28), bi => B(28), p => pi_matrix_0_28_port
                           , g => gi_matrix_0_28_port);
   PG_i_29 : pgb_3 port map( ai => A(29), bi => B(29), p => pi_matrix_0_29_port
                           , g => gi_matrix_0_29_port);
   PG_i_30 : pgb_2 port map( ai => A(30), bi => B(30), p => pi_matrix_0_30_port
                           , g => gi_matrix_0_30_port);
   PG_i_31 : pgb_1 port map( ai => A(31), bi => B(31), p => pi_matrix_0_31_port
                           , g => gi_matrix_0_31_port);
   INITIAL_PG_i_1_0 : PG_0 port map( Pik => pi_matrix_0_3_port, Pdkj => 
                           pi_matrix_0_2_port, Gik => gi_matrix_0_3_port, Gdkj 
                           => gi_matrix_0_2_port, Pij => pi_matrix_1_3_port, 
                           Gij => gi_matrix_1_3_port);
   INITIAL_G_i_1 : G_9 port map( Pik => pi_matrix_0_1_port, Gik => 
                           gi_matrix_0_1_port, Gdkj => gi_matrix_0_0_port, Gij 
                           => gi_matrix_1_1_port);
   INITIAL_G_i_2 : G_8 port map( Pik => pi_matrix_1_3_port, Gik => 
                           gi_matrix_1_3_port, Gdkj => gi_matrix_1_1_port, Gij 
                           => Co_0_port);
   PG_i_2_1_0 : PG_27 port map( Pik => pi_matrix_0_7_port, Pdkj => 
                           pi_matrix_0_6_port, Gik => gi_matrix_0_7_port, Gdkj 
                           => gi_matrix_0_6_port, Pij => pi_matrix_1_7_port, 
                           Gij => gi_matrix_1_7_port);
   PG_i_2_1_1 : PG_26 port map( Pik => pi_matrix_0_5_port, Pdkj => 
                           pi_matrix_0_4_port, Gik => gi_matrix_0_5_port, Gdkj 
                           => gi_matrix_0_4_port, Pij => pi_matrix_1_5_port, 
                           Gij => gi_matrix_1_5_port);
   PG_i_2_2_0 : PG_25 port map( Pik => pi_matrix_1_7_port, Pdkj => 
                           pi_matrix_1_5_port, Gik => gi_matrix_1_7_port, Gdkj 
                           => gi_matrix_1_5_port, Pij => pi_matrix_2_7_port, 
                           Gij => gi_matrix_2_7_port);
   FINAL_G_i_2 : G_7 port map( Pik => pi_matrix_2_7_port, Gik => 
                           gi_matrix_2_7_port, Gdkj => Co_0_port, Gij => 
                           Co_1_port);
   PG_i_3_1_0 : PG_24 port map( Pik => pi_matrix_0_11_port, Pdkj => 
                           pi_matrix_0_10_port, Gik => gi_matrix_0_11_port, 
                           Gdkj => gi_matrix_0_10_port, Pij => 
                           pi_matrix_1_11_port, Gij => gi_matrix_1_11_port);
   PG_i_3_1_1 : PG_23 port map( Pik => pi_matrix_0_9_port, Pdkj => 
                           pi_matrix_0_8_port, Gik => gi_matrix_0_9_port, Gdkj 
                           => gi_matrix_0_8_port, Pij => pi_matrix_1_9_port, 
                           Gij => gi_matrix_1_9_port);
   PG_i_3_2_0 : PG_22 port map( Pik => pi_matrix_1_11_port, Pdkj => 
                           pi_matrix_1_9_port, Gik => gi_matrix_1_11_port, Gdkj
                           => gi_matrix_1_9_port, Pij => pi_matrix_2_11_port, 
                           Gij => gi_matrix_2_11_port);
   FINAL_G_i_3 : G_6 port map( Pik => pi_matrix_2_11_port, Gik => 
                           gi_matrix_2_11_port, Gdkj => Co_1_port, Gij => 
                           Co_2_port);
   PG_i_4_1_0 : PG_21 port map( Pik => pi_matrix_0_15_port, Pdkj => 
                           pi_matrix_0_14_port, Gik => gi_matrix_0_15_port, 
                           Gdkj => gi_matrix_0_14_port, Pij => 
                           pi_matrix_1_15_port, Gij => gi_matrix_1_15_port);
   PG_i_4_1_1 : PG_20 port map( Pik => pi_matrix_0_13_port, Pdkj => 
                           pi_matrix_0_12_port, Gik => gi_matrix_0_13_port, 
                           Gdkj => gi_matrix_0_12_port, Pij => 
                           pi_matrix_1_13_port, Gij => gi_matrix_1_13_port);
   PG_i_4_2_0 : PG_19 port map( Pik => pi_matrix_1_15_port, Pdkj => 
                           pi_matrix_1_13_port, Gik => gi_matrix_1_15_port, 
                           Gdkj => gi_matrix_1_13_port, Pij => 
                           pi_matrix_2_15_port, Gij => gi_matrix_2_15_port);
   REMAINING_PG_i_4_2 : PG_18 port map( Pik => pi_matrix_2_15_port, Pdkj => 
                           pi_matrix_2_11_port, Gik => gi_matrix_2_15_port, 
                           Gdkj => gi_matrix_2_11_port, Pij => 
                           pi_matrix_3_15_port, Gij => gi_matrix_3_15_port);
   FINAL_G_i_4 : G_5 port map( Pik => pi_matrix_3_15_port, Gik => 
                           gi_matrix_3_15_port, Gdkj => Co_1_port, Gij => 
                           Co_3_port);
   PG_i_5_1_0 : PG_17 port map( Pik => pi_matrix_0_19_port, Pdkj => 
                           pi_matrix_0_18_port, Gik => gi_matrix_0_19_port, 
                           Gdkj => gi_matrix_0_18_port, Pij => 
                           pi_matrix_1_19_port, Gij => gi_matrix_1_19_port);
   PG_i_5_1_1 : PG_16 port map( Pik => pi_matrix_0_17_port, Pdkj => 
                           pi_matrix_0_16_port, Gik => gi_matrix_0_17_port, 
                           Gdkj => gi_matrix_0_16_port, Pij => 
                           pi_matrix_1_17_port, Gij => gi_matrix_1_17_port);
   PG_i_5_2_0 : PG_15 port map( Pik => pi_matrix_1_19_port, Pdkj => 
                           pi_matrix_1_17_port, Gik => gi_matrix_1_19_port, 
                           Gdkj => gi_matrix_1_17_port, Pij => 
                           pi_matrix_2_19_port, Gij => gi_matrix_2_19_port);
   REMAINING_PG_i_5_2 : PG_14 port map( Pik => pi_matrix_2_19_port, Pdkj => 
                           pi_matrix_2_15_port, Gik => gi_matrix_2_19_port, 
                           Gdkj => gi_matrix_2_15_port, Pij => 
                           pi_matrix_3_19_port, Gij => gi_matrix_3_19_port);
   FINAL_G_i_5 : G_4 port map( Pik => pi_matrix_3_19_port, Gik => 
                           gi_matrix_3_19_port, Gdkj => Co_3_port, Gij => 
                           Co_4_port);
   PG_i_6_1_0 : PG_13 port map( Pik => pi_matrix_0_23_port, Pdkj => 
                           pi_matrix_0_22_port, Gik => gi_matrix_0_23_port, 
                           Gdkj => gi_matrix_0_22_port, Pij => 
                           pi_matrix_1_23_port, Gij => gi_matrix_1_23_port);
   PG_i_6_1_1 : PG_12 port map( Pik => pi_matrix_0_21_port, Pdkj => 
                           pi_matrix_0_20_port, Gik => gi_matrix_0_21_port, 
                           Gdkj => gi_matrix_0_20_port, Pij => 
                           pi_matrix_1_21_port, Gij => gi_matrix_1_21_port);
   PG_i_6_2_0 : PG_11 port map( Pik => pi_matrix_1_23_port, Pdkj => 
                           pi_matrix_1_21_port, Gik => gi_matrix_1_23_port, 
                           Gdkj => gi_matrix_1_21_port, Pij => 
                           pi_matrix_2_23_port, Gij => gi_matrix_2_23_port);
   REMAINING_PG_i_6_2 : PG_10 port map( Pik => pi_matrix_2_23_port, Pdkj => 
                           pi_matrix_2_19_port, Gik => gi_matrix_2_23_port, 
                           Gdkj => gi_matrix_2_19_port, Pij => 
                           pi_matrix_3_23_port, Gij => gi_matrix_3_23_port);
   FINAL_G_i_6 : G_3 port map( Pik => pi_matrix_3_23_port, Gik => 
                           gi_matrix_3_23_port, Gdkj => Co_3_port, Gij => 
                           Co_5_port);
   PG_i_7_1_0 : PG_9 port map( Pik => pi_matrix_0_27_port, Pdkj => 
                           pi_matrix_0_26_port, Gik => gi_matrix_0_27_port, 
                           Gdkj => gi_matrix_0_26_port, Pij => 
                           pi_matrix_1_27_port, Gij => gi_matrix_1_27_port);
   PG_i_7_1_1 : PG_8 port map( Pik => pi_matrix_0_25_port, Pdkj => 
                           pi_matrix_0_24_port, Gik => gi_matrix_0_25_port, 
                           Gdkj => gi_matrix_0_24_port, Pij => 
                           pi_matrix_1_25_port, Gij => gi_matrix_1_25_port);
   PG_i_7_2_0 : PG_7 port map( Pik => pi_matrix_1_27_port, Pdkj => 
                           pi_matrix_1_25_port, Gik => gi_matrix_1_27_port, 
                           Gdkj => gi_matrix_1_25_port, Pij => 
                           pi_matrix_2_27_port, Gij => gi_matrix_2_27_port);
   REMAINING_PG_i_7_2 : PG_6 port map( Pik => pi_matrix_2_27_port, Pdkj => 
                           pi_matrix_2_23_port, Gik => gi_matrix_2_27_port, 
                           Gdkj => gi_matrix_2_23_port, Pij => 
                           pi_matrix_3_27_port, Gij => gi_matrix_3_27_port);
   FINAL_G_i_7 : G_2 port map( Pik => pi_matrix_3_27_port, Gik => 
                           gi_matrix_3_27_port, Gdkj => Co_3_port, Gij => 
                           Co_6_port);
   PG_i_8_1_0 : PG_5 port map( Pik => pi_matrix_0_31_port, Pdkj => 
                           pi_matrix_0_30_port, Gik => gi_matrix_0_31_port, 
                           Gdkj => gi_matrix_0_30_port, Pij => 
                           pi_matrix_1_31_port, Gij => gi_matrix_1_31_port);
   PG_i_8_1_1 : PG_4 port map( Pik => pi_matrix_0_29_port, Pdkj => 
                           pi_matrix_0_28_port, Gik => gi_matrix_0_29_port, 
                           Gdkj => gi_matrix_0_28_port, Pij => 
                           pi_matrix_1_29_port, Gij => gi_matrix_1_29_port);
   PG_i_8_2_0 : PG_3 port map( Pik => pi_matrix_1_31_port, Pdkj => 
                           pi_matrix_1_29_port, Gik => gi_matrix_1_31_port, 
                           Gdkj => gi_matrix_1_29_port, Pij => 
                           pi_matrix_2_31_port, Gij => gi_matrix_2_31_port);
   REMAINING_PG_i_8_2 : PG_2 port map( Pik => pi_matrix_2_31_port, Pdkj => 
                           pi_matrix_2_27_port, Gik => gi_matrix_2_31_port, 
                           Gdkj => gi_matrix_2_27_port, Pij => 
                           pi_matrix_3_31_port, Gij => gi_matrix_3_31_port);
   REMAINING_PG_i_8_3 : PG_1 port map( Pik => pi_matrix_3_31_port, Pdkj => 
                           pi_matrix_3_23_port, Gik => gi_matrix_3_31_port, 
                           Gdkj => gi_matrix_3_23_port, Pij => 
                           pi_matrix_4_31_port, Gij => gi_matrix_4_31_port);
   FINAL_G_i_8 : G_1 port map( Pik => pi_matrix_4_31_port, Gik => 
                           gi_matrix_4_31_port, Gdkj => Co_3_port, Gij => 
                           Co_7_port);

end SYN_structural_generic;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_adder_generic_NBIT32_NBIT_PER_BLOCK4.all;

entity adder_generic_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic;  S : out std_logic_vector (31 downto 0));

end adder_generic_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_add_struct of adder_generic_NBIT32_NBIT_PER_BLOCK4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GENERATOR_GENERIC_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CLA_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal carries_7_port, carries_6_port, carries_5_port, carries_4_port, 
      carries_3_port, carries_2_port, carries_1_port, xored_B_31_port, 
      xored_B_30_port, xored_B_29_port, xored_B_28_port, xored_B_27_port, 
      xored_B_26_port, xored_B_25_port, xored_B_24_port, xored_B_23_port, 
      xored_B_22_port, xored_B_21_port, xored_B_20_port, xored_B_19_port, 
      xored_B_18_port, xored_B_17_port, xored_B_16_port, xored_B_15_port, 
      xored_B_14_port, xored_B_13_port, xored_B_12_port, xored_B_11_port, 
      xored_B_10_port, xored_B_9_port, xored_B_8_port, xored_B_7_port, 
      xored_B_6_port, xored_B_5_port, xored_B_4_port, xored_B_3_port, 
      xored_B_2_port, xored_B_1_port, xored_B_0_port : std_logic;

begin
   
   carry : CLA_NBIT32_NBIT_PER_BLOCK4 port map( A(31) => A(31), A(30) => A(30),
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => xored_B_31_port, B(30) 
                           => xored_B_30_port, B(29) => xored_B_29_port, B(28) 
                           => xored_B_28_port, B(27) => xored_B_27_port, B(26) 
                           => xored_B_26_port, B(25) => xored_B_25_port, B(24) 
                           => xored_B_24_port, B(23) => xored_B_23_port, B(22) 
                           => xored_B_22_port, B(21) => xored_B_21_port, B(20) 
                           => xored_B_20_port, B(19) => xored_B_19_port, B(18) 
                           => xored_B_18_port, B(17) => xored_B_17_port, B(16) 
                           => xored_B_16_port, B(15) => xored_B_15_port, B(14) 
                           => xored_B_14_port, B(13) => xored_B_13_port, B(12) 
                           => xored_B_12_port, B(11) => xored_B_11_port, B(10) 
                           => xored_B_10_port, B(9) => xored_B_9_port, B(8) => 
                           xored_B_8_port, B(7) => xored_B_7_port, B(6) => 
                           xored_B_6_port, B(5) => xored_B_5_port, B(4) => 
                           xored_B_4_port, B(3) => xored_B_3_port, B(2) => 
                           xored_B_2_port, B(1) => xored_B_1_port, B(0) => 
                           xored_B_0_port, Cin => Cin, Co(7) => Cout, Co(6) => 
                           carries_7_port, Co(5) => carries_6_port, Co(4) => 
                           carries_5_port, Co(3) => carries_4_port, Co(2) => 
                           carries_3_port, Co(1) => carries_2_port, Co(0) => 
                           carries_1_port);
   sum : SUM_GENERATOR_GENERIC_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => 
                           A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => xored_B_31_port, B(30) => xored_B_30_port, 
                           B(29) => xored_B_29_port, B(28) => xored_B_28_port, 
                           B(27) => xored_B_27_port, B(26) => xored_B_26_port, 
                           B(25) => xored_B_25_port, B(24) => xored_B_24_port, 
                           B(23) => xored_B_23_port, B(22) => xored_B_22_port, 
                           B(21) => xored_B_21_port, B(20) => xored_B_20_port, 
                           B(19) => xored_B_19_port, B(18) => xored_B_18_port, 
                           B(17) => xored_B_17_port, B(16) => xored_B_16_port, 
                           B(15) => xored_B_15_port, B(14) => xored_B_14_port, 
                           B(13) => xored_B_13_port, B(12) => xored_B_12_port, 
                           B(11) => xored_B_11_port, B(10) => xored_B_10_port, 
                           B(9) => xored_B_9_port, B(8) => xored_B_8_port, B(7)
                           => xored_B_7_port, B(6) => xored_B_6_port, B(5) => 
                           xored_B_5_port, B(4) => xored_B_4_port, B(3) => 
                           xored_B_3_port, B(2) => xored_B_2_port, B(1) => 
                           xored_B_1_port, B(0) => xored_B_0_port, Ci(7) => 
                           carries_7_port, Ci(6) => carries_6_port, Ci(5) => 
                           carries_5_port, Ci(4) => carries_4_port, Ci(3) => 
                           carries_3_port, Ci(2) => carries_2_port, Ci(1) => 
                           carries_1_port, Ci(0) => Cin, S(31) => S(31), S(30) 
                           => S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));
   U33 : XOR2_X1 port map( A => Cin, B => B(9), Z => xored_B_9_port);
   U34 : XOR2_X1 port map( A => Cin, B => B(8), Z => xored_B_8_port);
   U35 : XOR2_X1 port map( A => Cin, B => B(7), Z => xored_B_7_port);
   U36 : XOR2_X1 port map( A => Cin, B => B(6), Z => xored_B_6_port);
   U37 : XOR2_X1 port map( A => Cin, B => B(5), Z => xored_B_5_port);
   U38 : XOR2_X1 port map( A => Cin, B => B(4), Z => xored_B_4_port);
   U39 : XOR2_X1 port map( A => Cin, B => B(3), Z => xored_B_3_port);
   U40 : XOR2_X1 port map( A => Cin, B => B(31), Z => xored_B_31_port);
   U41 : XOR2_X1 port map( A => Cin, B => B(30), Z => xored_B_30_port);
   U42 : XOR2_X1 port map( A => Cin, B => B(2), Z => xored_B_2_port);
   U43 : XOR2_X1 port map( A => Cin, B => B(29), Z => xored_B_29_port);
   U44 : XOR2_X1 port map( A => Cin, B => B(28), Z => xored_B_28_port);
   U45 : XOR2_X1 port map( A => Cin, B => B(27), Z => xored_B_27_port);
   U46 : XOR2_X1 port map( A => Cin, B => B(26), Z => xored_B_26_port);
   U47 : XOR2_X1 port map( A => Cin, B => B(25), Z => xored_B_25_port);
   U48 : XOR2_X1 port map( A => Cin, B => B(24), Z => xored_B_24_port);
   U49 : XOR2_X1 port map( A => Cin, B => B(23), Z => xored_B_23_port);
   U50 : XOR2_X1 port map( A => Cin, B => B(22), Z => xored_B_22_port);
   U51 : XOR2_X1 port map( A => Cin, B => B(21), Z => xored_B_21_port);
   U52 : XOR2_X1 port map( A => Cin, B => B(20), Z => xored_B_20_port);
   U53 : XOR2_X1 port map( A => Cin, B => B(1), Z => xored_B_1_port);
   U54 : XOR2_X1 port map( A => Cin, B => B(19), Z => xored_B_19_port);
   U55 : XOR2_X1 port map( A => Cin, B => B(18), Z => xored_B_18_port);
   U56 : XOR2_X1 port map( A => Cin, B => B(17), Z => xored_B_17_port);
   U57 : XOR2_X1 port map( A => Cin, B => B(16), Z => xored_B_16_port);
   U58 : XOR2_X1 port map( A => Cin, B => B(15), Z => xored_B_15_port);
   U59 : XOR2_X1 port map( A => Cin, B => B(14), Z => xored_B_14_port);
   U60 : XOR2_X1 port map( A => Cin, B => B(13), Z => xored_B_13_port);
   U61 : XOR2_X1 port map( A => Cin, B => B(12), Z => xored_B_12_port);
   U62 : XOR2_X1 port map( A => Cin, B => B(11), Z => xored_B_11_port);
   U63 : XOR2_X1 port map( A => Cin, B => B(10), Z => xored_B_10_port);
   U64 : XOR2_X1 port map( A => Cin, B => B(0), Z => xored_B_0_port);

end SYN_add_struct;
