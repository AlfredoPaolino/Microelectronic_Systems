
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_WRF_generic_M8_N8_F8_DATA_BIT32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_WRF_generic_M8_N8_F8_DATA_BIT32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_generic_M8_N8_F8_DATA_BIT32.all;

entity physicalRF_M8_N8_F8_DATA_BIT32 is

   port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADDR_WR, ADDR_RD1, 
         ADDR_RD2 : in std_logic_vector (7 downto 0);  DATA_IN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end physicalRF_M8_N8_F8_DATA_BIT32;

architecture SYN_beh of physicalRF_M8_N8_F8_DATA_BIT32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
      n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, 
      n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, 
      n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, 
      n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, 
      n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, 
      n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, 
      n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004
      , n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
      n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, 
      n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, 
      n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, 
      n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, 
      n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, 
      n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, 
      n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, 
      n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, 
      n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, 
      n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, 
      n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, 
      n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, 
      n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, 
      n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, 
      n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, 
      n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, 
      n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, 
      n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, 
      n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, 
      n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, 
      n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, 
      n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, 
      n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, 
      n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, 
      n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, 
      n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, 
      n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, 
      n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, 
      n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, 
      n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, 
      n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, 
      n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, 
      n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, 
      n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, 
      n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, 
      n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, 
      n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, 
      n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, 
      n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, 
      n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, 
      n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, 
      n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, 
      n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, 
      n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, 
      n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, 
      n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, 
      n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, 
      n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, 
      n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, 
      n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, 
      n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, 
      n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, 
      n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, 
      n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, 
      n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, 
      n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, 
      n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, 
      n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, 
      n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, 
      n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, 
      n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, 
      n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, 
      n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, 
      n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, 
      n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, 
      n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, 
      n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, 
      n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, 
      n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, 
      n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, 
      n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, 
      n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, 
      n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, 
      n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, 
      n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, 
      n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, 
      n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, 
      n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, 
      n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, 
      n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, 
      n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, 
      n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, 
      n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, 
      n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, 
      n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, 
      n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, 
      n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, 
      n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, 
      n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, 
      n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, 
      n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, 
      n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, 
      n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, 
      n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, 
      n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, 
      n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, 
      n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, 
      n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, 
      n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, 
      n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, 
      n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, 
      n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, 
      n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, 
      n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, 
      n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, 
      n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, 
      n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, 
      n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, 
      n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, 
      n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, 
      n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, 
      n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, 
      n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, 
      n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, 
      n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, 
      n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, 
      n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, 
      n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, 
      n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, 
      n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, 
      n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, 
      n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, 
      n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, 
      n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, 
      n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, 
      n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, 
      n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, 
      n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, 
      n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, 
      n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, 
      n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, 
      n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, 
      n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, 
      n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, 
      n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, 
      n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, 
      n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, 
      n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, 
      n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, 
      n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, 
      n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, 
      n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, 
      n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, 
      n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, 
      n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, 
      n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, 
      n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, 
      n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, 
      n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, 
      n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, 
      n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, 
      n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, 
      n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, 
      n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, 
      n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, 
      n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, 
      n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, 
      n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, 
      n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, 
      n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, 
      n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, 
      n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, 
      n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, 
      n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, 
      n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, 
      n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, 
      n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, 
      n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, 
      n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, 
      n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, 
      n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, 
      n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, 
      n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, 
      n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, 
      n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, 
      n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, 
      n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, 
      n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, 
      n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, 
      n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, 
      n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, 
      n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, 
      n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, 
      n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, 
      n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, 
      n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, 
      n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, 
      n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, 
      n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, 
      n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, 
      n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, 
      n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, 
      n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, 
      n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, 
      n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, 
      n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, 
      n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, 
      n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, 
      n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, 
      n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, 
      n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, 
      n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, 
      n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, 
      n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, 
      n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, 
      n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, 
      n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, 
      n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, 
      n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, 
      n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, 
      n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, 
      n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, 
      n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, 
      n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, 
      n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, 
      n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, 
      n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, 
      n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, 
      n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, 
      n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, 
      n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, 
      n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, 
      n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, 
      n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, 
      n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, 
      n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, 
      n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, 
      n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, 
      n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, 
      n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, 
      n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, 
      n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, 
      n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, 
      n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, 
      n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, 
      n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, 
      n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, 
      n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, 
      n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, 
      n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, 
      n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, 
      n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, 
      n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, 
      n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, 
      n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, 
      n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, 
      n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, 
      n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, 
      n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, 
      n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, 
      n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, 
      n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, 
      n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, 
      n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, 
      n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, 
      n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, 
      n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, 
      n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, 
      n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, 
      n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, 
      n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, 
      n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, 
      n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, 
      n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, 
      n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, 
      n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, 
      n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, 
      n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, 
      n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, 
      n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, 
      n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, 
      n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, 
      n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, 
      n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, 
      n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, 
      n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, 
      n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, 
      n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, 
      n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, 
      n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, 
      n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, 
      n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, 
      n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, 
      n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, 
      n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, 
      n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, 
      n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, 
      n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, 
      n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, 
      n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, 
      n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, 
      n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, 
      n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, 
      n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, 
      n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, 
      n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, 
      n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, 
      n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, 
      n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, 
      n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, 
      n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, 
      n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, 
      n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, 
      n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, 
      n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, 
      n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, 
      n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, 
      n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, 
      n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, 
      n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, 
      n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, 
      n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, 
      n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, 
      n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, 
      n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, 
      n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, 
      n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, 
      n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, 
      n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, 
      n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, 
      n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, 
      n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, 
      n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, 
      n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, 
      n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, 
      n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, 
      n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, 
      n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, 
      n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, 
      n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, 
      n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, 
      n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, 
      n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, 
      n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, 
      n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, 
      n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, 
      n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, 
      n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, 
      n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, 
      n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, 
      n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, 
      n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, 
      n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, 
      n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, 
      n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, 
      n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, 
      n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, 
      n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, 
      n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, 
      n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, 
      n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, 
      n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, 
      n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, 
      n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, 
      n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, 
      n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, 
      n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, 
      n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, 
      n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, 
      n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, 
      n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, 
      n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, 
      n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, 
      n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, 
      n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, 
      n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, 
      n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, 
      n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, 
      n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, 
      n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, 
      n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, 
      n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, 
      n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, 
      n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, 
      n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, 
      n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, 
      n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, 
      n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, 
      n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, 
      n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, 
      n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, 
      n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, 
      n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, 
      n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, 
      n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, 
      n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, 
      n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, 
      n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, 
      n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, 
      n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, 
      n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, 
      n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, 
      n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, 
      n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, 
      n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, 
      n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, 
      n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, 
      n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, 
      n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, 
      n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, 
      n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, 
      n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, 
      n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, 
      n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, 
      n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, 
      n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, 
      n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, 
      n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, 
      n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, 
      n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, 
      n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, 
      n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, 
      n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, 
      n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, 
      n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, 
      n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, 
      n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, 
      n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, 
      n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, 
      n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, 
      n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, 
      n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, 
      n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, 
      n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, 
      n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, 
      n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, 
      n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, 
      n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, 
      n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, 
      n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, 
      n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, 
      n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, 
      n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, 
      n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, 
      n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, 
      n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, 
      n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, 
      n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, 
      n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, 
      n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, 
      n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, 
      n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, 
      n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, 
      n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, 
      n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, 
      n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, 
      n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, 
      n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, 
      n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, 
      n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, 
      n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, 
      n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, 
      n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, 
      n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, 
      n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, 
      n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, 
      n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, 
      n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, 
      n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, 
      n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, 
      n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, 
      n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, 
      n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, 
      n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, 
      n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, 
      n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, 
      n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, 
      n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, 
      n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, 
      n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, 
      n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, 
      n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, 
      n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, 
      n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, 
      n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, 
      n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, 
      n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, 
      n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, 
      n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, 
      n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, 
      n14334, n14335, n14336, n14337, n14338, n14339, n14340, n50932, n50933, 
      n50934, n50935, n50936, n50937, n50938, n50939, n50964, n50965, n50966, 
      n50967, n50968, n50969, n50970, n50971, n51600, n51601, n51602, n51603, 
      n51604, n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612, 
      n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620, n51621, 
      n51622, n51623, n51624, n51625, n51626, n51627, n51628, n51629, n51630, 
      n51631, n51632, n51633, n51634, n51635, n51636, n51637, n51638, n51639, 
      n51640, n51641, n51642, n51643, n51644, n51645, n51646, n51647, n51648, 
      n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51664, n51665, 
      n51666, n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674, 
      n51675, n51676, n51677, n51678, n51679, n51712, n51713, n51714, n51715, 
      n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724, 
      n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733, 
      n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742, 
      n51743, n51760, n51761, n51762, n51763, n51764, n51765, n51766, n51767, 
      n51768, n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776, 
      n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51808, n51809, 
      n51810, n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818, 
      n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826, n52160, 
      n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168, n52169, 
      n52170, n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178, 
      n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187, 
      n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196, 
      n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204, n52205, 
      n52206, n52207, n52236, n52237, n52238, n52239, n52240, n52241, n52242, 
      n52243, n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275, 
      n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316, 
      n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324, n52325, 
      n52326, n52327, n52328, n52329, n52330, n52331, n52351, n52352, n52353, 
      n52354, n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362, 
      n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371, 
      n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380, 
      n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388, n52389, 
      n52390, n52496, n52497, n52498, n52499, n52500, n52501, n52502, n52503, 
      n52504, n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512, 
      n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520, n52521, 
      n52522, n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530, 
      n52531, n52532, n52533, n52534, n52535, n52584, n52585, n52586, n52587, 
      n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, 
      n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, 
      n52606, n52607, n52656, n52657, n52658, n52659, n52660, n52661, n52662, 
      n52663, n52664, n52665, n52666, n52667, n52668, n52669, n52670, n52671, 
      n52672, n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52728, 
      n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736, n52737, 
      n52738, n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746, 
      n52747, n52748, n52749, n52750, n52751, n52760, n52761, n52762, n52763, 
      n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772, 
      n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780, n52781, 
      n52782, n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790, 
      n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798, n52799, 
      n52800, n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52856, 
      n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864, n52865, 
      n52866, n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874, 
      n52875, n52876, n52877, n52878, n52879, n52928, n52929, n52930, n52931, 
      n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940, 
      n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948, n52949, 
      n52950, n52951, n52952, n52953, n52954, n52955, n52956, n52957, n52958, 
      n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966, n52967, 
      n52968, n52969, n52970, n52971, n52972, n52973, n52974, n52975, n52976, 
      n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984, n52985, 
      n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994, 
      n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002, n53003, 
      n53028, n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036, 
      n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044, n53045, 
      n53046, n53047, n53048, n53049, n53050, n53051, n53124, n53125, n53126, 
      n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134, n53135, 
      n53136, n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144, 
      n53145, n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153, 
      n53154, n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162, 
      n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171, 
      n53172, n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180, 
      n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188, n53189, 
      n53190, n53191, n53192, n53193, n53194, n53195, n53244, n53245, n53246, 
      n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254, n53255, 
      n53256, n53257, n53356, n53357, n53358, n53359, n53360, n53361, n53362, 
      n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371, 
      n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380, 
      n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389, 
      n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398, 
      n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406, n53407, 
      n53408, n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416, 
      n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425, 
      n53426, n53427, n53476, n53477, n53478, n53479, n53480, n53481, n53482, 
      n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490, n53491, 
      n53492, n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53548, 
      n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556, n53557, 
      n53558, n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566, 
      n53567, n53568, n53569, n53570, n53571, n53572, n53573, n53574, n53575, 
      n53576, n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53632, 
      n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641, 
      n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650, 
      n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659, 
      n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668, 
      n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677, 
      n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686, 
      n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694, n53695, 
      n53696, n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704, 
      n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713, 
      n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722, 
      n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731, 
      n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740, 
      n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748, n53749, 
      n53750, n53751, n53916, n53917, n53918, n53919, n53920, n53921, n53922, 
      n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930, n53931, 
      n53932, n53933, n53934, n53935, n53936, n53937, n53938, n53939, n53940, 
      n53941, n53942, n53943, n53944, n53945, n53946, n53947, n53948, n53949, 
      n53950, n53951, n53952, n53953, n53954, n53955, n53956, n53957, n53958, 
      n53959, n53960, n53961, n53962, n53963, n53964, n53965, n53966, n53967, 
      n53968, n53969, n53970, n53971, n53972, n53973, n53974, n53975, n53976, 
      n53977, n53978, n53979, n53980, n53981, n53982, n53983, n53984, n53985, 
      n53986, n53987, n54156, n54157, n54158, n54159, n54160, n54161, n54162, 
      n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170, n54171, 
      n54172, n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180, 
      n54181, n54182, n54183, n54184, n54185, n54186, n54187, n54188, n54189, 
      n54190, n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198, 
      n54199, n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207, 
      n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216, 
      n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225, 
      n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234, 
      n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243, 
      n54244, n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252, 
      n54253, n54254, n54255, n54256, n54257, n54258, n54259, n54260, n54261, 
      n54262, n54263, n54264, n54265, n54266, n54267, n54268, n54269, n54270, 
      n54271, n54272, n54273, n54274, n54275, n54324, n54325, n54326, n54327, 
      n54328, n54329, n54330, n54331, n54332, n54333, n54334, n54335, n54336, 
      n54337, n54338, n54339, n54340, n54341, n54342, n54343, n54344, n54345, 
      n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354, 
      n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362, n54363, 
      n54364, n54365, n54366, n54367, n54368, n54369, n54370, n54371, n54372, 
      n54373, n54374, n54375, n54376, n54377, n54378, n54379, n54380, n54381, 
      n54382, n54383, n54384, n54385, n54386, n54387, n54388, n54389, n54390, 
      n54391, n54392, n54393, n54394, n54395, n54396, n54397, n54398, n54399, 
      n54400, n54401, n54402, n54403, n54404, n54405, n54406, n54407, n54408, 
      n54409, n54410, n54411, n54412, n54413, n54414, n54415, n54416, n54417, 
      n54418, n54419, n54444, n54445, n54446, n54447, n54448, n54449, n54450, 
      n54451, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
      n351, n352, n353, n354, n355, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n519, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, 
      n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
      n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
      n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
      n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
      n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, 
      n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
      n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, 
      n758, n759, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, 
      n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, 
      n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, 
      n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, 
      n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, 
      n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, 
      n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, 
      n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, 
      n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
      n970, n971, n996, n997, n998, n999, n1518, n1567, n1568, n1569, n1570, 
      n1571, n1572, n1573, n1574, n1639, n1640, n1641, n1642, n1643, n1644, 
      n1645, n1646, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
      n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
      n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
      n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3099, n3100, 
      n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, 
      n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, 
      n3121, n3122, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, 
      n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, 
      n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, 
      n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, 
      n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, 
      n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, 
      n9341, n9342, n9343, n9344, n9345, n9346, n9603, n9604, n9605, n9606, 
      n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, 
      n9617, n9618, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, 
      n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, 
      n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, 
      n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, 
      n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, 
      n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, 
      n9805, n9806, n9807, n9808, n9809, n9810, n15171, n15172, n15173, n15174,
      n15175, n15176, n15177, n15203, n15204, n15205, n15206, n15207, n15208, 
      n15209, n15210, n15299, n15300, n15301, n15302, n15303, n15304, n15305, 
      n15306, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, 
      n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486, n54487, 
      n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496, 
      n54497, n54498, n54499, n54500, n54501, n54502, n54504, n54505, n54506, 
      n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514, n54515, 
      n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523, n54524, 
      n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532, n54533, 
      n54534, n54535, n54543, n54544, n54545, n54546, n54547, n54548, n54549, 
      n54550, n54551, n54552, n54553, n54558, n54563, n54564, n54570, n54571, 
      n54572, n54573, n54574, n54575, n54623, n54624, n54625, n54626, n54627, 
      n54628, n54629, n54630, n54631, n54632, n54633, n54634, n54635, n54636, 
      n54637, n54638, n54639, n54640, n54641, n54642, n54643, n54644, n54645, 
      n54646, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n452, n474, 
      n475, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n776, n777, n778, n779, n780, 
      n781, n782, n783, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
      n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, 
      n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, 
      n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, 
      n861, n862, n863, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
      n1583, n1584, n1585, n1586, n1587, n1588, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2075, n2076, n2077, n2078, n2213, n2214, 
      n2215, n2216, n2217, n2218, n2219, n2220, n2235, n2236, n2237, n2238, 
      n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, 
      n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, 
      n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, 
      n2269, n2270, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2439, n2440, n2441, n2442, n2443, n2444, 
      n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, 
      n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2483, n2484, 
      n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
      n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, 
      n2505, n2506, n2507, n2508, n2509, n2510, n2645, n2646, n2647, n2648, 
      n2649, n2650, n2651, n2909, n2910, n2911, n2912, n2913, n2914, n2915, 
      n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n3409, 
      n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, 
      n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, 
      n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, 
      n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
      n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3621, n3622, n3623, 
      n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, 
      n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, 
      n3644, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, 
      n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, 
      n3986, n3987, n3988, n3989, n3990, n15363, n15364, n15365, n15366, n15367
      , n15368, n15369, n15370, n15411, n15412, n15413, n15414, n15415, n15416,
      n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, 
      n15426, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, 
      n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, 
      n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, 
      n15493, n15494, n15495, n15496, n15497, n15498, n15520, n15521, n15522, 
      n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, 
      n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15601, n15602, 
      n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15707, 
      n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, 
      n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15803, n15804, 
      n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, 
      n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, 
      n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, 
      n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, 
      n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, 
      n15850, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, 
      n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, 
      n498, n499, n560, n561, n562, n563, n564, n565, n566, n567, n760, n761, 
      n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
      n774, n775, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, 
      n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, 
      n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n972, n973, 
      n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, 
      n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n1000, n1001,
      n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, 
      n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, 
      n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, 
      n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, 
      n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, 
      n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, 
      n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
      n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, 
      n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, 
      n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, 
      n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, 
      n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, 
      n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
      n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, 
      n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, 
      n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, 
      n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, 
      n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, 
      n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, 
      n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, 
      n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, 
      n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, 
      n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
      n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, 
      n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, 
      n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, 
      n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, 
      n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, 
      n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, 
      n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
      n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, 
      n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, 
      n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, 
      n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, 
      n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, 
      n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, 
      n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, 
      n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
      n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
      n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
      n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
      n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
      n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, 
      n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, 
      n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, 
      n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, 
      n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
      n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, 
      n1512, n1513, n1514, n1515, n1516, n1517, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1589, n1590, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, 
      n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, 
      n1665, n1666, n1667, n1668, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
      n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1813, n1814, n1815, 
      n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
      n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, 
      n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, 
      n1846, n1847, n1848, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
      n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
      n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2221, n2222, n2223, n2224, 
      n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, 
      n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
      n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
      n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2436, n2437, n2438, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2511, n2512, n2513, n2514, 
      n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
      n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
      n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, 
      n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, 
      n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, 
      n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, 
      n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, 
      n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, 
      n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, 
      n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
      n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, 
      n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, 
      n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, 
      n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, 
      n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, 
      n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2701, n2702, n2703, 
      n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
      n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
      n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
      n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
      n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
      n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, 
      n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, 
      n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
      n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2839, n2840, n2841, 
      n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, 
      n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, 
      n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, 
      n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
      n2882, n2883, n2884, n2885, n2886, n2907, n2908, n2925, n2926, n2927, 
      n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, 
      n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, 
      n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, 
      n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, 
      n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, 
      n2978, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, 
      n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, 
      n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, 
      n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, 
      n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, 
      n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, 
      n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, 
      n3096, n3097, n3098, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
      n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, 
      n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, 
      n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, 
      n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, 
      n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
      n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, 
      n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
      n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
      n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
      n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, 
      n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, 
      n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, 
      n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, 
      n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
      n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
      n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, 
      n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, 
      n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, 
      n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, 
      n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, 
      n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, 
      n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, 
      n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, 
      n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, 
      n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, 
      n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, 
      n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3457, 
      n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, 
      n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, 
      n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, 
      n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, 
      n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, 
      n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, 
      n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, 
      n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, 
      n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, 
      n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, 
      n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, 
      n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, 
      n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, 
      n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, 
      n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, 
      n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, 
      n3618, n3619, n3620, n3645, n3646, n3647, n3648, n3649, n3650, n3651, 
      n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, 
      n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, 
      n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, 
      n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, 
      n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, 
      n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, 
      n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, 
      n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, 
      n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
      n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, 
      n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, 
      n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, 
      n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, 
      n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, 
      n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, 
      n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, 
      n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, 
      n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, 
      n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, 
      n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, 
      n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, 
      n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, 
      n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, 
      n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, 
      n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, 
      n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, 
      n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3927, n3928, n3929, 
      n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, 
      n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, 
      n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, 
      n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3991, n3992, n3993, 
      n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, 
      n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, 
      n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, 
      n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, 
      n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, 
      n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, 
      n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, 
      n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, 
      n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, 
      n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, 
      n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, 
      n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, 
      n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, 
      n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, 
      n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, 
      n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, 
      n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, 
      n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
      n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, 
      n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, 
      n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, 
      n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
      n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, 
      n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, 
      n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, 
      n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
      n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, 
      n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, 
      n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, 
      n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
      n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
      n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, 
      n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, 
      n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
      n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, 
      n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, 
      n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
      n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, 
      n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, 
      n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, 
      n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, 
      n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
      n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, 
      n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, 
      n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, 
      n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, 
      n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, 
      n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, 
      n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, 
      n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, 
      n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, 
      n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, 
      n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, 
      n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, 
      n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, 
      n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
      n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, 
      n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, 
      n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, 
      n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, 
      n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, 
      n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, 
      n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, 
      n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, 
      n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, 
      n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
      n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, 
      n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, 
      n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, 
      n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, 
      n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, 
      n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, 
      n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, 
      n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
      n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, 
      n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, 
      n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, 
      n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, 
      n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, 
      n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, 
      n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5276, n5277, 
      n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5287, n5288, n5289, 
      n5290, n5293, n5297, n5300, n5306, n5307, n5308, n5309, n5313, n5314, 
      n5315, n5316, n5319, n5321, n5322, n5324, n5325, n5326, n5327, n5331, 
      n5333, n5334, n5335, n5338, n5339, n5342, n5343, n5346, n5347, n5348, 
      n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, 
      n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, 
      n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, 
      n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, 
      n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, 
      n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, 
      n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, 
      n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, 
      n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, 
      n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, 
      n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, 
      n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, 
      n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, 
      n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, 
      n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, 
      n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, 
      n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, 
      n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, 
      n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, 
      n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, 
      n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, 
      n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, 
      n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, 
      n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, 
      n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, 
      n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, 
      n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, 
      n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, 
      n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, 
      n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, 
      n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, 
      n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, 
      n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, 
      n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, 
      n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, 
      n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, 
      n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, 
      n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, 
      n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, 
      n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, 
      n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, 
      n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, 
      n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, 
      n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, 
      n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, 
      n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, 
      n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, 
      n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, 
      n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, 
      n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, 
      n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, 
      n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, 
      n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, 
      n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, 
      n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, 
      n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, 
      n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, 
      n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, 
      n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, 
      n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, 
      n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, 
      n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, 
      n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, 
      n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, 
      n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, 
      n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, 
      n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6018, n6019, 
      n6021, n6022, n6023, n6025, n6026, n6027, n6028, n6029, n6030, n6031, 
      n6032, n6033, n6034, n6035, n6037, n6038, n6039, n6040, n6041, n6042, 
      n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, 
      n6054, n6056, n6057, n6059, n6060, n6062, n6063, n6064, n6065, n6066, 
      n6067, n6068, n6069, n6070, n6071, n6073, n6074, n6075, n6076, n6078, 
      n6079, n6080, n6081, n6082, n6083, n6084, n6086, n6087, n6089, n6090, 
      n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, 
      n6102, n6103, n6104, n6105, n6107, n6108, n6109, n6110, n6111, n6112, 
      n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, 
      n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, 
      n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, 
      n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, 
      n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, 
      n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, 
      n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, 
      n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, 
      n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, 
      n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, 
      n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, 
      n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, 
      n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, 
      n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, 
      n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, 
      n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, 
      n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, 
      n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, 
      n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, 
      n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, 
      n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, 
      n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, 
      n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, 
      n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, 
      n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, 
      n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, 
      n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, 
      n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, 
      n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, 
      n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, 
      n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, 
      n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, 
      n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, 
      n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, 
      n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, 
      n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, 
      n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, 
      n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, 
      n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, 
      n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, 
      n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, 
      n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, 
      n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, 
      n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, 
      n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, 
      n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, 
      n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, 
      n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, 
      n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, 
      n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, 
      n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, 
      n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, 
      n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, 
      n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, 
      n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, 
      n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, 
      n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, 
      n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, 
      n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, 
      n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, 
      n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, 
      n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, 
      n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, 
      n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, 
      n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, 
      n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, 
      n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, 
      n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, 
      n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, 
      n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, 
      n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, 
      n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, 
      n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, 
      n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, 
      n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, 
      n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, 
      n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, 
      n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, 
      n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, 
      n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, 
      n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, 
      n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, 
      n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, 
      n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, 
      n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, 
      n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, 
      n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, 
      n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, 
      n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, 
      n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, 
      n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, 
      n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, 
      n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, 
      n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, 
      n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, 
      n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, 
      n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, 
      n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, 
      n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, 
      n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, 
      n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, 
      n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, 
      n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, 
      n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, 
      n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, 
      n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, 
      n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, 
      n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, 
      n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, 
      n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, 
      n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, 
      n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, 
      n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, 
      n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, 
      n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, 
      n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, 
      n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, 
      n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, 
      n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, 
      n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, 
      n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, 
      n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, 
      n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, 
      n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, 
      n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, 
      n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, 
      n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, 
      n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, 
      n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, 
      n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, 
      n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, 
      n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, 
      n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, 
      n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, 
      n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, 
      n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, 
      n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, 
      n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, 
      n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, 
      n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, 
      n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, 
      n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, 
      n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, 
      n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, 
      n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, 
      n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, 
      n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, 
      n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, 
      n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, 
      n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, 
      n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, 
      n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, 
      n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, 
      n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, 
      n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, 
      n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, 
      n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, 
      n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, 
      n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, 
      n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, 
      n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, 
      n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, 
      n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, 
      n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, 
      n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, 
      n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, 
      n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, 
      n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, 
      n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, 
      n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, 
      n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, 
      n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, 
      n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, 
      n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, 
      n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, 
      n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, 
      n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, 
      n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, 
      n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, 
      n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, 
      n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, 
      n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, 
      n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, 
      n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, 
      n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, 
      n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, 
      n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, 
      n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, 
      n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, 
      n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, 
      n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, 
      n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, 
      n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, 
      n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, 
      n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, 
      n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, 
      n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, 
      n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, 
      n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, 
      n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, 
      n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, 
      n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, 
      n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, 
      n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, 
      n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, 
      n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, 
      n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, 
      n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, 
      n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, 
      n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, 
      n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, 
      n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, 
      n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, 
      n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, 
      n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, 
      n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, 
      n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, 
      n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, 
      n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, 
      n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, 
      n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, 
      n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, 
      n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, 
      n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, 
      n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, 
      n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, 
      n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, 
      n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, 
      n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, 
      n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, 
      n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, 
      n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, 
      n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, 
      n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, 
      n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, 
      n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, 
      n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, 
      n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, 
      n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, 
      n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, 
      n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, 
      n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, 
      n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, 
      n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, 
      n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, 
      n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, 
      n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, 
      n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, 
      n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, 
      n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, 
      n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, 
      n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, 
      n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, 
      n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, 
      n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, 
      n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, 
      n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, 
      n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, 
      n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, 
      n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, 
      n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, 
      n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, 
      n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, 
      n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, 
      n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, 
      n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, 
      n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, 
      n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, 
      n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, 
      n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, 
      n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, 
      n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, 
      n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, 
      n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, 
      n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, 
      n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, 
      n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, 
      n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, 
      n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, 
      n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, 
      n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, 
      n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, 
      n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, 
      n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, 
      n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, 
      n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, 
      n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, 
      n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, 
      n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, 
      n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, 
      n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, 
      n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, 
      n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, 
      n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, 
      n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, 
      n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, 
      n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, 
      n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, 
      n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, 
      n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, 
      n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, 
      n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, 
      n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, 
      n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, 
      n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, 
      n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, 
      n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, 
      n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, 
      n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, 
      n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, 
      n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, 
      n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, 
      n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, 
      n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, 
      n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, 
      n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, 
      n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, 
      n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, 
      n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, 
      n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, 
      n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, 
      n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, 
      n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, 
      n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, 
      n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, 
      n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, 
      n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, 
      n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, 
      n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, 
      n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, 
      n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, 
      n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, 
      n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, 
      n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, 
      n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, 
      n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, 
      n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, 
      n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, 
      n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, 
      n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, 
      n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, 
      n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, 
      n9597, n9598, n9599, n9600, n9601, n9602, n9619, n9620, n9621, n9622, 
      n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, 
      n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, 
      n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, 
      n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, 
      n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, 
      n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, 
      n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, 
      n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, 
      n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, 
      n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, 
      n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, 
      n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, 
      n9743, n9744, n9745, n9746, n9811, n9812, n9813, n9814, n9815, n9816, 
      n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, 
      n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, 
      n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, 
      n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, 
      n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, 
      n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, 
      n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, 
      n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, 
      n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, 
      n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, 
      n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n14341, n14342, 
      n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, 
      n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, 
      n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, 
      n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, 
      n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, 
      n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, 
      n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, 
      n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, 
      n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, 
      n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, 
      n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, 
      n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, 
      n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, 
      n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, 
      n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, 
      n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, 
      n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, 
      n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, 
      n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, 
      n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, 
      n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, 
      n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, 
      n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, 
      n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, 
      n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, 
      n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, 
      n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, 
      n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, 
      n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, 
      n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, 
      n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, 
      n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, 
      n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, 
      n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, 
      n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, 
      n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, 
      n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, 
      n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, 
      n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, 
      n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, 
      n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, 
      n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, 
      n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, 
      n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, 
      n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, 
      n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, 
      n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, 
      n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, 
      n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, 
      n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, 
      n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, 
      n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, 
      n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, 
      n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, 
      n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, 
      n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, 
      n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, 
      n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, 
      n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, 
      n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, 
      n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, 
      n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, 
      n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, 
      n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, 
      n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, 
      n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, 
      n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, 
      n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, 
      n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, 
      n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, 
      n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, 
      n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, 
      n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, 
      n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, 
      n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, 
      n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, 
      n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, 
      n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, 
      n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, 
      n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, 
      n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, 
      n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, 
      n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, 
      n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, 
      n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, 
      n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, 
      n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, 
      n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, 
      n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, 
      n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, 
      n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, 
      n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, 
      n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, 
      n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, 
      n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15211, n15212, 
      n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, 
      n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, 
      n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, 
      n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, 
      n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, 
      n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, 
      n15267, n15268, n15269, n15270, n15279, n15280, n15281, n15282, n15283, 
      n15284, n15285, n15286, n15287, n15316, n15317, n15318, n15319, n15320, 
      n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, 
      n15330, n15343, n15380, n15381, n15382, n15383, n15384, n15385, n15386, 
      n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15427, 
      n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, 
      n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, 
      n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, 
      n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, 
      n15464, n15465, n15466, n15499, n15500, n15501, n15502, n15503, n15504, 
      n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, 
      n15514, n15515, n15516, n15517, n15518, n15519, n15587, n15588, n15589, 
      n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, 
      n15599, n15600, n15611, n15612, n15663, n15666, n15669, n15672, n15675, 
      n15678, n15681, n15684, n15685, n15688, n15691, n15694, n15697, n15700, 
      n15703, n15706, n15726, n15729, n15748, n15749, n15750, n15751, n15752, 
      n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, 
      n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, 
      n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, 
      n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, 
      n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, 
      n15798, n15799, n15800, n15801, n15802, n15851, n15852, n15853, n15854, 
      n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, 
      n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, 
      n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, 
      n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, 
      n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, 
      n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, 
      n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15918, n15919, 
      n15922, n15947, n15950, n15951, n15954, n15955, n15958, n15959, n15962, 
      n15963, n15966, n15967, n15970, n15971, n16100, n16101, n16102, n16103, 
      n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, 
      n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, 
      n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, 
      n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, 
      n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, 
      n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, 
      n16158, n16189, n16190, n16195, n16196, n16201, n16202, n16207, n16208, 
      n16231, n16232, n16237, n16238, n16243, n16244, n16249, n16250, n16255, 
      n16256, n16279, n16280, n16298, n16300, n16302, n16304, n16306, n16308, 
      n16320, n16322, n16324, n16326, n16328, n16330, n16332, n16334, n16341, 
      n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, 
      n16351, n16352, n16353, n16354, n16355, n16356, n16413, n16414, n16415, 
      n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, 
      n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, 
      n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, 
      n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, 
      n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, 
      n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, 
      n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, 
      n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, 
      n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, 
      n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, 
      n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, 
      n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, 
      n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, 
      n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, 
      n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, 
      n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, 
      n16560, n16561, n16562, n16563, n16588, n16589, n16590, n16591, n16592, 
      n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, 
      n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, 
      n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, 
      n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, 
      n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, 
      n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, 
      n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, 
      n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, 
      n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, 
      n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, 
      n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, 
      n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, 
      n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, 
      n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, 
      n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, 
      n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, 
      n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, 
      n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, 
      n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, 
      n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, 
      n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, 
      n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, 
      n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, 
      n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, 
      n16809, n16810, n16811, n16812, n16813, n16830, n16831, n16832, n16833, 
      n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, 
      n16843, n16844, n16845, n59635, n59636, n59637, n59638, n59639, n59640, 
      n59641, n59642, n59643, n59644, n59645, n59646, n59647, n59648, n59649, 
      n59650, n59651, n59652, n59653, n59654, n59655, n59656, n59657, n59658, 
      n59659, n59660, n59661, n59662, n59663, n59664, n59665, n59666, n59667, 
      n59668, n59669, n59670, n59671, n59672, n59673, n59674, n59675, n59676, 
      n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684, n59685, 
      n59686, n59687, n59688, n59689, n59690, n59691, n59692, n59693, n59694, 
      n59695, n59696, n59697, n59698, n59699, n59700, n59701, n59702, n59703, 
      n59704, n59705, n59706, n59707, n59708, n59709, n59710, n59711, n59712, 
      n59713, n59714, n59715, n59716, n59717, n59718, n59719, n59720, n59721, 
      n59722, n59723, n59724, n59725, n59726, n59727, n59728, n59729, n59730, 
      n59731, n59732, n59733, n59734, n59735, n59736, n59737, n59738, n59739, 
      n59740, n59741, n59742, n59743, n59744, n59745, n59746, n59747, n59748, 
      n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59756, n59757, 
      n59758, n59759, n59760, n59761, n59762, n59763, n59764, n59765, n59766, 
      n59767, n59768, n59769, n59770, n59771, n59772, n59773, n59774, n59775, 
      n59776, n59777, n59778, n59779, n59780, n59781, n59782, n59783, n59784, 
      n59785, n59786, n59787, n59788, n59789, n59790, n59791, n59792, n59793, 
      n59794, n59795, n59796, n59797, n59798, n59799, n59800, n59801, n59802, 
      n59803, n59804, n59805, n59806, n59807, n59808, n59809, n59810, n59811, 
      n59812, n59813, n59814, n59815, n59816, n59817, n59818, n59819, n59820, 
      n59821, n59822, n59823, n59824, n59825, n59826, n59827, n59828, n59829, 
      n59830, n59831, n59832, n59833, n59834, n59835, n59836, n59837, n59838, 
      n59839, n59840, n59841, n59842, n59843, n59844, n59845, n59846, n59847, 
      n59848, n59849, n59850, n59851, n59852, n59853, n59854, n59855, n59856, 
      n59857, n59858, n59859, n59860, n59861, n59862, n59863, n59864, n59865, 
      n59866, n59867, n59868, n59869, n59870, n59871, n59872, n59873, n59874, 
      n59875, n59876, n59877, n59878, n59879, n59880, n59881, n59882, n59883, 
      n59884, n59885, n59886, n59887, n59888, n59889, n59890, n59891, n59892, 
      n59893, n59894, n59895, n59896, n59897, n59898, n59899, n59900, n59901, 
      n59902, n59903, n59904, n59905, n59906, n59907, n59908, n59909, n59910, 
      n59911, n59912, n59913, n59914, n59915, n59916, n59917, n59918, n59919, 
      n59920, n59921, n59922, n59923, n59924, n59925, n59926, n59927, n59928, 
      n59929, n59930, n59931, n59932, n59933, n59934, n59935, n59936, n59937, 
      n59938, n59939, n59940, n59941, n59942, n59943, n59944, n59945, n59946, 
      n59947, n59948, n59949, n59950, n59951, n59952, n59953, n59954, n59955, 
      n59956, n59957, n59958, n59959, n59960, n59961, n59962, n59963, n59964, 
      n59965, n59966, n59967, n59968, n59969, n59970, n59971, n59972, n59973, 
      n59974, n59975, n59976, n59977, n59978, n59979, n59980, n59981, n59982, 
      n59983, n59984, n59985, n59986, n59987, n59988, n59989, n59990, n59991, 
      n59992, n59993, n59994, n59995, n59996, n59997, n59998, n59999, n60000, 
      n60001, n60002, n60003, n60004, n60005, n60006, n60007, n60008, n60009, 
      n60010, n60011, n60012, n60013, n60014, n60015, n60016, n60017, n60018, 
      n60019, n60020, n60021, n60022, n60023, n60024, n60025, n60026, n60027, 
      n60028, n60029, n60030, n60031, n60032, n60033, n60034, n60035, n60036, 
      n60037, n60038, n60039, n60040, n60041, n60042, n60043, n60044, n60045, 
      n60046, n60047, n60048, n60049, n60050, n60051, n60052, n60053, n60054, 
      n60055, n60056, n60057, n60058, n60059, n60060, n60061, n60062, n60063, 
      n60064, n60065, n60066, n60067, n60068, n60069, n60070, n60071, n60072, 
      n60073, n60074, n60075, n60076, n60077, n60078, n60079, n60080, n60081, 
      n60082, n60083, n60084, n60085, n60086, n60087, n60088, n60089, n60090, 
      n60091, n60092, n60093, n60094, n60095, n60096, n60097, n60098, n60099, 
      n60100, n60101, n60102, n60103, n60104, n60105, n60106, n60107, n60108, 
      n60109, n60110, n60111, n60112, n60113, n60114, n60115, n60116, n60117, 
      n60118, n60119, n60120, n60121, n60122, n60123, n60124, n60125, n60126, 
      n60127, n60128, n60129, n60130, n60131, n60132, n60133, n60134, n60135, 
      n60136, n60137, n60138, n60139, n60140, n60141, n60142, n60143, n60144, 
      n60145, n60146, n60147, n60148, n60149, n60150, n60151, n60152, n60153, 
      n60154, n60155, n60156, n60157, n60158, n60159, n60160, n60161, n60162, 
      n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170, n60171, 
      n60172, n60173, n60174, n60175, n60176, n60177, n60178, n60179, n60180, 
      n60181, n60182, n60183, n60184, n60185, n60186, n60187, n60188, n60189, 
      n60190, n60191, n60192, n60193, n60194, n60195, n60196, n60197, n60198, 
      n60199, n60200, n60201, n60202, n60203, n60204, n60205, n60206, n60207, 
      n60208, n60209, n60210, n60211, n60212, n60213, n60214, n60215, n60216, 
      n60217, n60218, n60219, n60220, n60221, n60222, n60223, n60224, n60225, 
      n60226, n60227, n60228, n60229, n60230, n60231, n60232, n60233, n60234, 
      n60235, n60236, n60237, n60238, n60239, n60240, n60241, n60242, n60243, 
      n60244, n60245, n60246, n60247, n60248, n60249, n60250, n60251, n60252, 
      n60253, n60254, n60255, n60256, n60257, n60258, n60259, n60260, n60261, 
      n60262, n60263, n60264, n60265, n60266, n60267, n60268, n60269, n60270, 
      n60271, n60272, n60273, n60274, n60275, n60276, n60277, n60278, n60279, 
      n60280, n60281, n60282, n60283, n60284, n60285, n60286, n60287, n60288, 
      n60289, n60290, n60291, n60292, n60293, n60294, n60295, n60296, n60297, 
      n60298, n60299, n60300, n60301, n60302, n60303, n60304, n60305, n60306, 
      n60307, n60308, n60309, n60310, n60311, n60312, n60313, n60314, n60315, 
      n60316, n60317, n60318, n60319, n60320, n60321, n60322, n60323, n60324, 
      n60325, n60326, n60327, n60328, n60329, n60330, n60331, n60332, n60333, 
      n60334, n60335, n60336, n60337, n60338, n60339, n60340, n60341, n60342, 
      n60343, n60344, n60345, n60346, n60347, n60348, n60349, n60350, n60351, 
      n60352, n60353, n60354, n60355, n60356, n60357, n60358, n60359, n60360, 
      n60361, n60362, n60363, n60364, n60365, n60366, n60367, n60368, n60369, 
      n60370, n60371, n60372, n60373, n60374, n60375, n60376, n60377, n60378, 
      n60379, n60380, n60381, n60382, n60383, n60384, n60385, n60386, n60387, 
      n60388, n60389, n60390, n60391, n60392, n60393, n60394, n60395, n60396, 
      n60397, n60398, n60399, n60400, n60401, n60402, n60403, n60404, n60405, 
      n60406, n60407, n60408, n60409, n60410, n60411, n60412, n60413, n60414, 
      n60415, n60416, n60417, n60418, n60419, n60420, n60421, n60422, n60423, 
      n60424, n60425, n60426, n60427, n60428, n60429, n60430, n60431, n60432, 
      n60433, n60434, n60435, n60436, n60437, n60438, n60439, n60440, n60441, 
      n60442, n60443, n60444, n60445, n60446, n60447, n60448, n60449, n60450, 
      n60451, n60452, n60453, n60454, n60455, n60456, n60457, n60458, n60459, 
      n60460, n60461, n60462, n60463, n60464, n60465, n60466, n60467, n60468, 
      n60469, n60470, n60471, n60472, n60473, n60474, n60475, n60476, n60477, 
      n60478, n60479, n60480, n60481, n60482, n60483, n60484, n60485, n60486, 
      n60487, n60488, n60489, n60490, n60491, n60492, n60493, n60494, n60495, 
      n60496, n60497, n60498, n60499, n60500, n60501, n60502, n60503, n60504, 
      n60505, n60506, n60507, n60508, n60509, n60510, n60511, n60512, n60513, 
      n60514, n60515, n60516, n60517, n60518, n60519, n60520, n60521, n60522, 
      n60523, n60524, n60525, n60526, n60527, n60528, n60529, n60530, n60531, 
      n60532, n60533, n60534, n60535, n60536, n60537, n60538, n60539, n60540, 
      n60541, n60542, n60543, n60544, n60545, n60546, n60547, n60548, n60549, 
      n60550, n60551, n60552, n60553, n60554, n60555, n60556, n60557, n60558, 
      n60559, n60560, n60561, n60562, n60563, n60564, n60565, n60566, n60567, 
      n60568, n60569, n60570, n60571, n60572, n60573, n60574, n60575, n60576, 
      n60577, n60578, n60579, n60580, n60581, n60582, n60583, n60584, n60585, 
      n60586, n60587, n60588, n60589, n60590, n60591, n60592, n60593, n60594, 
      n60595, n60596, n60597, n60598, n60599, n60600, n60601, n60602, n60603, 
      n60604, n60605, n60606, n60607, n60608, n60609, n60610, n60611, n60612, 
      n60613, n60614, n60615, n60616, n60617, n60618, n60619, n60620, n60621, 
      n60622, n60623, n60624, n60625, n60626, n60627, n60628, n60629, n60630, 
      n60631, n60632, n60633, n60634, n60635, n60636, n60637, n60638, n60639, 
      n60640, n60641, n60642, n60643, n60644, n60645, n60646, n60647, n60648, 
      n60649, n60650, n60651, n60652, n60653, n60654, n60655, n60656, n60657, 
      n60658, n60659, n60660, n60661, n60662, n60663, n60664, n60665, n60666, 
      n60667, n60668, n60669, n60670, n60671, n60672, n60673, n60674, n60675, 
      n60676, n60677, n60678, n60679, n60680, n60681, n60682, n60683, n60684, 
      n60685, n60686, n60687, n60688, n60689, n60690, n60691, n60692, n60693, 
      n60694, n60695, n60696, n60697, n60698, n60699, n60700, n60701, n60702, 
      n60703, n60704, n60705, n60706, n60707, n60708, n60709, n60710, n60711, 
      n60712, n60713, n60714, n60715, n60716, n60717, n60718, n60719, n60720, 
      n60721, n60722, n60723, n60724, n60725, n60726, n60727, n60728, n60729, 
      n60730, n60731, n60732, n60733, n60734, n60735, n60736, n60737, n60738, 
      n60739, n60740, n60741, n60742, n60743, n60744, n60745, n60746, n60747, 
      n60748, n60749, n60750, n60751, n60752, n60753, n60754, n60755, n60756, 
      n60757, n60758, n60759, n60760, n60761, n60762, n60763, n60764, n60765, 
      n60766, n60767, n60768, n60769, n60770, n60771, n60772, n60773, n60774, 
      n60775, n60776, n60777, n60778, n60779, n60780, n60781, n60782, n60783, 
      n60784, n60785, n60786, n60787, n60788, n60789, n60790, n60791, n60792, 
      n60793, n60794, n60795, n60796, n60797, n60798, n60799, n60800, n60801, 
      n60802, n60803, n60804, n60805, n60806, n60807, n60808, n60809, n60810, 
      n60811, n60812, n60813, n60814, n60815, n60816, n60817, n60818, n60819, 
      n60820, n60821, n60822, n60823, n60824, n60825, n60826, n60827, n60828, 
      n60829, n60830, n60831, n60832, n60833, n60834, n60835, n60836, n60837, 
      n60838, n60839, n60840, n60841, n60842, n60843, n60844, n60845, n60846, 
      n60847, n60848, n60849, n60850, n60851, n60852, n60853, n60854, n60855, 
      n60856, n60857, n60858, n60859, n60860, n60861, n60862, n60863, n60864, 
      n60865, n60866, n60867, n60868, n60869, n60870, n60871, n60872, n60873, 
      n60874, n60875, n60876, n60877, n60878, n60879, n60880, n60881, n60882, 
      n60883, n60884, n60885, n60886, n60887, n60888, n60889, n60890, n60891, 
      n60892, n60893, n60894, n60895, n60896, n60897, n60898, n60899, n60900, 
      n60901, n60902, n60903, n60904, n60905, n60906, n60907, n60908, n60909, 
      n60910, n60911, n60912, n60913, n60914, n60915, n60916, n60917, n60918, 
      n60919, n60920, n60921, n60922, n60923, n60924, n60925, n60926, n60927, 
      n60928, n60929, n60930, n60931, n60932, n60933, n60934, n60935, n60936, 
      n60937, n60938, n60939, n60940, n60941, n60942, n60943, n60944, n60945, 
      n60946, n60947, n60948, n60949, n60950, n60951, n60952, n60953, n60954, 
      n60955, n60956, n60957, n60958, n60959, n60960, n60961, n60962, n60963, 
      n60964, n60965, n60966, n60967, n60968, n60969, n60970, n60971, n60972, 
      n60973, n60974, n60975, n60976, n60977, n60978, n60979, n60980, n60981, 
      n60982, n60983, n60984, n60985, n60986, n60987, n60988, n60989, n60990, 
      n60991, n60992, n60993, n60994, n60995, n60996, n60997, n60998, n60999, 
      n61000, n61001, n61002, n61003, n61004, n61005, n61006, n61007, n61008, 
      n61009, n61010, n61011, n61012, n61013, n61014, n61015, n61016, n61017, 
      n61018, n61019, n61020, n61021, n61022, n61023, n61024, n61025, n61026, 
      n61027, n61028, n61029, n61030, n61031, n61032, n61033, n61034, n61035, 
      n61036, n61037, n61038, n61039, n61040, n61041, n61042, n61043, n61044, 
      n61045, n61046, n61047, n61048, n61049, n61050, n61051, n61052, n61053, 
      n61054, n61055, n61056, n61057, n61058, n61059, n61060, n61061, n61062, 
      n61063, n61064, n61065, n61066, n61067, n61068, n61069, n61070, n61071, 
      n61072, n61073, n61074, n61075, n61076, n61077, n61078, n61079, n61080, 
      n61081, n61082, n61083, n61084, n61085, n61086, n61087, n61088, n61089, 
      n61090, n61091, n61092, n61093, n61094, n61095, n61096, n61097, n61098, 
      n61099, n61100, n61101, n61102, n61103, n61104, n61105, n61106, n61107, 
      n61108, n61109, n61110, n61111, n61112, n61113, n61114, n61115, n61116, 
      n61117, n61118, n61119, n61120, n61121, n61122, n61123, n61124, n61125, 
      n61126, n61127, n61128, n61129, n61130, n61131, n61132, n61133, n61134, 
      n61135, n61136, n61137, n61138, n61139, n61140, n61141, n61142, n61143, 
      n61144, n61145, n61146, n61147, n61148, n61149, n61150, n61151, n61152, 
      n61153, n61154, n61155, n61156, n61157, n61158, n61159, n61160, n61161, 
      n61162, n61163, n61164, n61165, n61166, n61167, n61168, n61169, n61170, 
      n61171, n61172, n61173, n61174, n61175, n61176, n61177, n61178, n61179, 
      n61180, n61181, n61182, n61183, n61184, n61185, n61186, n61187, n61188, 
      n61189, n61190, n61191, n61192, n61193, n61194, n61195, n61196, n61197, 
      n61198, n61199, n61200, n61201, n61202, n61203, n61204, n61205, n61206, 
      n61207, n61208, n61209, n61210, n61211, n61212, n61213, n61214, n61215, 
      n61216, n61217, n61218, n61219, n61220, n61221, n61222, n61223, n61224, 
      n61225, n61226, n61227, n61228, n61229, n61230, n61231, n61232, n61233, 
      n61234, n61235, n61236, n61237, n61238, n61239, n61240, n61241, n61242, 
      n61243, n61244, n61245, n61246, n61247, n61248, n61249, n61250, n61251, 
      n61252, n61253, n61254, n61255, n61256, n61257, n61258, n61259, n61260, 
      n61261, n61262, n61263, n61264, n61265, n61266, n61267, n61268, n61269, 
      n61270, n61271, n61272, n61273, n61274, n61275, n61276, n61277, n61278, 
      n61279, n61280, n61281, n61282, n61283, n61284, n61285, n61286, n61287, 
      n61288, n61289, n61290, n61291, n61292, n61293, n61294, n61295, n61296, 
      n61297, n61298, n61299, n61300, n61301, n61302, n61303, n61304, n61305, 
      n61306, n61307, n61308, n61309, n61310, n61311, n61312, n61313, n61314, 
      n61315, n61316, n61317, n61318, n61319, n61320, n61321, n61322, n61323, 
      n61324, n61325, n61326, n61327, n61328, n61329, n61330, n61331, n61332, 
      n61333, n61334, n61335, n61336, n61337, n61338, n61339, n61340, n61341, 
      n61342, n61343, n61344, n61345, n61346, n61347, n61348, n61349, n61350, 
      n61351, n61352, n61353, n61354, n61355, n61356, n61357, n61358, n61359, 
      n61360, n61361, n61362, n61363, n61364, n61365, n61366, n61367, n61368, 
      n61369, n61370, n61371, n61372, n61373, n61374, n61375, n61376, n61377, 
      n61378, n61379, n61380, n61381, n61382, n61383, n61384, n61385, n61386, 
      n61387, n61388, n61389, n61390, n61391, n61392, n61393, n61394, n61395, 
      n61396, n61397, n61398, n61399, n61400, n61401, n61402, n61403, n61404, 
      n61405, n61406, n61407, n61408, n61409, n61410, n61411, n61412, n61413, 
      n61414, n61415, n61416, n61417, n61418, n61419, n61420, n61421, n61422, 
      n61423, n61424, n61425, n61426, n61427, n61428, n61429, n61430, n61431, 
      n61432, n61433, n61434, n61435, n61436, n61437, n61438, n61439, n61440, 
      n61441, n61442, n61443, n61444, n61445, n61446, n61447, n61448, n61449, 
      n61450, n61451, n61452, n61453, n61454, n61455, n61456, n61457, n61458, 
      n61459, n61460, n61461, n61462, n61463, n61464, n61465, n61466, n61467, 
      n61468, n61469, n61470, n61471, n61472, n61473, n61474, n61475, n61476, 
      n61477, n61478, n61479, n61480, n61481, n61482, n61483, n61484, n61485, 
      n61486, n61487, n61488, n61489, n61490, n61491, n61492, n61493, n61494, 
      n61495, n61496, n61497, n61498, n61499, n61500, n61501, n61502, n61503, 
      n61504, n61505, n61506, n61507, n61508, n61509, n61510, n61511, n61512, 
      n61513, n61514, n61515, n61516, n61517, n61518, n61519, n61520, n61521, 
      n61522, n61523, n61524, n61525, n61526, n61527, n61528, n61529, n61530, 
      n61531, n61532, n61533, n61534, n61535, n61536, n61537, n61538, n61539, 
      n61540, n61541, n61542, n61543, n61544, n61545, n61546, n61547, n61548, 
      n61549, n61550, n61551, n61552, n61553, n61554, n61555, n61556, n61557, 
      n61558, n61559, n61560, n61561, n61562, n61563, n61564, n61565, n61566, 
      n61567, n61568, n61569, n61570, n61571, n61572, n61573, n61574, n61575, 
      n61576, n61577, n61578, n61579, n61580, n61581, n61582, n61583, n61584, 
      n61585, n61586, n61587, n61588, n61589, n61590, n61591, n61592, n61593, 
      n61594, n61595, n61596, n61597, n61598, n61599, n61600, n61601, n61602, 
      n61603, n61604, n61605, n61606, n61607, n61608, n61609, n61610, n61611, 
      n61612, n61613, n61614, n61615, n61616, n61617, n61618, n61619, n61620, 
      n61621, n61622, n61623, n61624, n61625, n61626, n61627, n61628, n61629, 
      n61630, n61631, n61632, n61633, n61634, n61635, n61636, n61637, n61638, 
      n61639, n61640, n61641, n61642, n61643, n61644, n61645, n61646, n61647, 
      n61648, n61649, n61650, n61651, n61652, n61653, n61654, n61655, n61656, 
      n61657, n61658, n61659, n61660, n61661, n61662, n61663, n61664, n61665, 
      n61666, n61667, n61668, n61669, n61670, n61671, n61672, n61673, n61674, 
      n61675, n61676, n61677, n61678, n61679, n61680, n61681, n61682, n61683, 
      n61684, n61685, n61686, n61687, n61688, n61689, n61690, n61691, n61692, 
      n61693, n61694, n61695, n61696, n61697, n61698, n61699, n61700, n61701, 
      n61702, n61703, n61704, n61705, n61706, n61707, n61708, n61709, n61710, 
      n61711, n61712, n61713, n61714, n61715, n61716, n61717, n61718, n61719, 
      n61720, n61721, n61722, n61723, n61724, n61725, n61726, n61727, n61728, 
      n61729, n61730, n61731, n61732, n61733, n61734, n61735, n61736, n61737, 
      n61738, n61739, n61740, n61741, n61742, n61743, n61744, n61745, n61746, 
      n61747, n61748, n61749, n61750, n61751, n61752, n61753, n61754, n61755, 
      n61756, n61757, n61758, n61759, n61760, n61761, n61762, n61763, n61764, 
      n61765, n61766, n61767, n61768, n61769, n61770, n61771, n61772, n61773, 
      n61774, n61775, n61776, n61777, n61778, n61779, n61780, n61781, n61782, 
      n61783, n61784, n61785, n61786, n61787, n61788, n61789, n61790, n61791, 
      n61792, n61793, n61794, n61795, n61796, n61797, n61798, n61799, n61800, 
      n61801, n61802, n61803, n61804, n61805, n61806, n61807, n61808, n61809, 
      n61810, n61811, n61812, n61813, n61814, n61815, n61816, n61817, n61818, 
      n61819, n61820, n61821, n61822, n61823, n61824, n61825, n61826, n61827, 
      n61828, n61829, n61830, n61831, n61832, n61833, n61834, n61835, n61836, 
      n61837, n61838, n61839, n61840, n61841, n61842, n61843, n61844, n61845, 
      n61846, n61847, n61848, n61849, n61850, n61851, n61852, n61853, n61854, 
      n61855, n61856, n61857, n61858, n61859, n61860, n61861, n61862, n61863, 
      n61864, n61865, n61866, n61867, n61868, n61869, n61870, n61871, n61872, 
      n61873, n61874, n61875, n61876, n61877, n61878, n61879, n61880, n61881, 
      n61882, n61883, n61884, n61885, n61886, n61887, n61888, n61889, n61890, 
      n61891, n61892, n61893, n61894, n61895, n61896, n61897, n61898, n61899, 
      n61900, n61901, n61902, n61903, n61904, n61905, n61906, n61907, n61908, 
      n61909, n61910, n61911, n61912, n61913, n61914, n61915, n61916, n61917, 
      n61918, n61919, n61920, n61921, n61922, n61923, n61924, n61925, n61926, 
      n61927, n61928, n61929, n61930, n61931, n61932, n61933, n61934, n61935, 
      n61936, n61937, n61938, n61939, n61940, n61941, n61942, n61943, n61944, 
      n61945, n61946, n61947, n61948, n61949, n61950, n61951, n61952, n61953, 
      n61954, n61955, n61956, n61957, n61958, n61959, n61960, n61961, n61962, 
      n61963, n61964, n61965, n61966, n61967, n61968, n61969, n61970, n61971, 
      n61972, n61973, n61974, n61975, n61976, n61977, n61978, n61979, n61980, 
      n61981, n61982, n61983, n61984, n61985, n61986, n61987, n61988, n61989, 
      n61990, n61991, n61992, n61993, n61994, n61995, n61996, n61997, n61998, 
      n61999, n62000, n62001, n62002, n62003, n62004, n62005, n62006, n62007, 
      n62008, n62009, n62010, n62011, n62012, n62013, n62014, n62015, n62016, 
      n62017, n62018, n62019, n62020, n62021, n62022, n62023, n62024, n62025, 
      n62026, n62027, n62028, n62029, n62030, n62031, n62032, n62033, n62034, 
      n62035, n62036, n62037, n62038, n62039, n62040, n62041, n62042, n62043, 
      n62044, n62045, n62046, n62047, n62048, n62049, n62050, n62051, n62052, 
      n62053, n62054, n62055, n62056, n62057, n62058, n62059, n62060, n62061, 
      n62062, n62063, n62064, n62065, n62066, n62067, n62068, n62069, n62070, 
      n62071, n62072, n62073, n62074, n62075, n62076, n62077, n62078, n62079, 
      n62080, n62081, n62082, n62083, n62084, n62085, n62086, n62087, n62088, 
      n62089, n62090, n62091, n62092, n62093, n62094, n62095, n62096, n62097, 
      n62098, n62099, n62100, n62101, n62102, n62103, n62104, n62105, n62106, 
      n62107, n62108, n62109, n62110, n62111, n62112, n62113, n62114, n62115, 
      n62116, n62117, n62118, n62119, n62120, n62121, n62122, n62123, n62124, 
      n62125, n62126, n62127, n62128, n62129, n62130, n62131, n62132, n62133, 
      n62134, n62135, n62136, n62137, n62138, n62139, n62140, n62141, n62142, 
      n62143, n62144, n62145, n62146, n62147, n62148, n62149, n62150, n62151, 
      n62152, n62153, n62154, n62155, n62156, n62157, n62158, n62159, n62160, 
      n62161, n62162, n62163, n62164, n62165, n62166, n62167, n62168, n62169, 
      n62170, n62171, n62172, n62173, n62174, n62175, n62176, n62177, n62178, 
      n62179, n62180, n62181, n62182, n62183, n62184, n62185, n62186, n62187, 
      n62188, n62189, n62190, n62191, n62192, n62193, n62194, n62195, n62196, 
      n62197, n62198, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, 
      n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, 
      n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, 
      n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, 
      n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, 
      n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, 
      n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, 
      n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, 
      n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, 
      n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, 
      n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, 
      n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, 
      n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, 
      n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, 
      n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, 
      n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, 
      n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, 
      n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, 
      n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, 
      n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, 
      n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, 
      n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, 
      n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, 
      n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, 
      n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, 
      n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, 
      n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, 
      n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, 
      n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, 
      n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, 
      n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, 
      n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, 
      n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, 
      n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, 
      n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, 
      n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, 
      n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, 
      n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, 
      n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, 
      n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, 
      n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, 
      n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, 
      n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, 
      n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, 
      n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, 
      n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, 
      n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, 
      n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, 
      n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, 
      n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, 
      n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, 
      n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, 
      n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, 
      n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, 
      n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, 
      n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, 
      n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, 
      n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, 
      n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, 
      n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, 
      n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, 
      n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, 
      n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, 
      n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, 
      n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, 
      n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, 
      n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, 
      n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, 
      n_2276, n_2277, n_2278, n_2279, n_2280, n_2281 : std_logic;

begin
   
   REGS_reg_94_23_inst : DFF_X1 port map( D => n11324, CK => CLK, Q => n59736, 
                           QN => n2645);
   REGS_reg_94_22_inst : DFF_X1 port map( D => n11323, CK => CLK, Q => n59735, 
                           QN => n2646);
   REGS_reg_94_21_inst : DFF_X1 port map( D => n11322, CK => CLK, Q => n59734, 
                           QN => n2647);
   REGS_reg_94_20_inst : DFF_X1 port map( D => n11321, CK => CLK, Q => n59733, 
                           QN => n2648);
   REGS_reg_94_19_inst : DFF_X1 port map( D => n11320, CK => CLK, Q => n59732, 
                           QN => n2649);
   REGS_reg_94_18_inst : DFF_X1 port map( D => n11319, CK => CLK, Q => n59731, 
                           QN => n2650);
   REGS_reg_94_17_inst : DFF_X1 port map( D => n11318, CK => CLK, Q => n59730, 
                           QN => n2651);
   REGS_reg_93_4_inst : DFF_X1 port map( D => n11337, CK => CLK, Q => n59693, 
                           QN => n160);
   REGS_reg_93_3_inst : DFF_X1 port map( D => n11336, CK => CLK, Q => n59692, 
                           QN => n161);
   REGS_reg_93_2_inst : DFF_X1 port map( D => n11335, CK => CLK, Q => n59691, 
                           QN => n162);
   REGS_reg_93_1_inst : DFF_X1 port map( D => n11334, CK => CLK, Q => n59690, 
                           QN => n163);
   REGS_reg_93_0_inst : DFF_X1 port map( D => n11333, CK => CLK, Q => n59689, 
                           QN => n164);
   REGS_reg_92_23_inst : DFF_X1 port map( D => n11388, CK => CLK, Q => n59709, 
                           QN => n165);
   REGS_reg_92_22_inst : DFF_X1 port map( D => n11387, CK => CLK, Q => n59708, 
                           QN => n166);
   REGS_reg_92_21_inst : DFF_X1 port map( D => n11386, CK => CLK, Q => n59707, 
                           QN => n167);
   REGS_reg_92_20_inst : DFF_X1 port map( D => n11385, CK => CLK, Q => n59706, 
                           QN => n168);
   REGS_reg_92_19_inst : DFF_X1 port map( D => n11384, CK => CLK, Q => n59705, 
                           QN => n169);
   REGS_reg_92_18_inst : DFF_X1 port map( D => n11383, CK => CLK, Q => n59704, 
                           QN => n170);
   REGS_reg_92_17_inst : DFF_X1 port map( D => n11382, CK => CLK, Q => n59703, 
                           QN => n171);
   REGS_reg_92_16_inst : DFF_X1 port map( D => n11381, CK => CLK, Q => n59702, 
                           QN => n172);
   REGS_reg_92_15_inst : DFF_X1 port map( D => n11380, CK => CLK, Q => n59701, 
                           QN => n173);
   REGS_reg_92_14_inst : DFF_X1 port map( D => n11379, CK => CLK, Q => n59700, 
                           QN => n174);
   REGS_reg_92_13_inst : DFF_X1 port map( D => n11378, CK => CLK, Q => n59699, 
                           QN => n175);
   REGS_reg_92_12_inst : DFF_X1 port map( D => n11377, CK => CLK, Q => n59698, 
                           QN => n176);
   REGS_reg_92_11_inst : DFF_X1 port map( D => n11376, CK => CLK, Q => n59697, 
                           QN => n177);
   REGS_reg_92_10_inst : DFF_X1 port map( D => n11375, CK => CLK, Q => n59696, 
                           QN => n178);
   REGS_reg_92_9_inst : DFF_X1 port map( D => n11374, CK => CLK, Q => n59695, 
                           QN => n179);
   REGS_reg_92_8_inst : DFF_X1 port map( D => n11373, CK => CLK, Q => n59694, 
                           QN => n180);
   REGS_reg_92_7_inst : DFF_X1 port map( D => n11372, CK => CLK, Q => n59717, 
                           QN => n181);
   REGS_reg_92_6_inst : DFF_X1 port map( D => n11371, CK => CLK, Q => n59716, 
                           QN => n182);
   REGS_reg_92_5_inst : DFF_X1 port map( D => n11370, CK => CLK, Q => n59715, 
                           QN => n183);
   REGS_reg_92_4_inst : DFF_X1 port map( D => n11369, CK => CLK, Q => n59714, 
                           QN => n184);
   REGS_reg_92_3_inst : DFF_X1 port map( D => n11368, CK => CLK, Q => n59713, 
                           QN => n185);
   REGS_reg_92_2_inst : DFF_X1 port map( D => n11367, CK => CLK, Q => n59712, 
                           QN => n186);
   REGS_reg_92_1_inst : DFF_X1 port map( D => n11366, CK => CLK, Q => n59711, 
                           QN => n187);
   REGS_reg_92_0_inst : DFF_X1 port map( D => n11365, CK => CLK, Q => n59710, 
                           QN => n188);
   REGS_reg_91_23_inst : DFF_X1 port map( D => n11420, CK => CLK, Q => n59664, 
                           QN => n189);
   REGS_reg_91_22_inst : DFF_X1 port map( D => n11419, CK => CLK, Q => n59663, 
                           QN => n190);
   REGS_reg_91_21_inst : DFF_X1 port map( D => n11418, CK => CLK, Q => n59662, 
                           QN => n191);
   REGS_reg_91_20_inst : DFF_X1 port map( D => n11417, CK => CLK, Q => n59661, 
                           QN => n192);
   REGS_reg_91_19_inst : DFF_X1 port map( D => n11416, CK => CLK, Q => n59660, 
                           QN => n193);
   REGS_reg_91_18_inst : DFF_X1 port map( D => n11415, CK => CLK, Q => n59659, 
                           QN => n194);
   REGS_reg_91_17_inst : DFF_X1 port map( D => n11414, CK => CLK, Q => n59658, 
                           QN => n195);
   REGS_reg_91_16_inst : DFF_X1 port map( D => n11413, CK => CLK, Q => n59657, 
                           QN => n196);
   REGS_reg_91_15_inst : DFF_X1 port map( D => n11412, CK => CLK, Q => n59656, 
                           QN => n197);
   REGS_reg_91_14_inst : DFF_X1 port map( D => n11411, CK => CLK, Q => n59655, 
                           QN => n198);
   REGS_reg_91_13_inst : DFF_X1 port map( D => n11410, CK => CLK, Q => n59654, 
                           QN => n199);
   REGS_reg_91_12_inst : DFF_X1 port map( D => n11409, CK => CLK, Q => n59653, 
                           QN => n200);
   REGS_reg_91_11_inst : DFF_X1 port map( D => n11408, CK => CLK, Q => n59652, 
                           QN => n201);
   REGS_reg_91_10_inst : DFF_X1 port map( D => n11407, CK => CLK, Q => n59651, 
                           QN => n202);
   REGS_reg_91_9_inst : DFF_X1 port map( D => n11406, CK => CLK, Q => n59650, 
                           QN => n203);
   REGS_reg_91_8_inst : DFF_X1 port map( D => n11405, CK => CLK, Q => n59649, 
                           QN => n204);
   REGS_reg_91_7_inst : DFF_X1 port map( D => n11404, CK => CLK, Q => n59672, 
                           QN => n205);
   REGS_reg_91_6_inst : DFF_X1 port map( D => n11403, CK => CLK, Q => n59671, 
                           QN => n206);
   REGS_reg_91_5_inst : DFF_X1 port map( D => n11402, CK => CLK, Q => n59670, 
                           QN => n207);
   REGS_reg_91_4_inst : DFF_X1 port map( D => n11401, CK => CLK, Q => n59669, 
                           QN => n208);
   REGS_reg_91_3_inst : DFF_X1 port map( D => n11400, CK => CLK, Q => n59668, 
                           QN => n209);
   REGS_reg_91_2_inst : DFF_X1 port map( D => n11399, CK => CLK, Q => n59667, 
                           QN => n210);
   REGS_reg_91_1_inst : DFF_X1 port map( D => n11398, CK => CLK, Q => n59666, 
                           QN => n211);
   REGS_reg_91_0_inst : DFF_X1 port map( D => n11397, CK => CLK, Q => n59665, 
                           QN => n212);
   REGS_reg_66_11_inst : DFF_X1 port map( D => n12208, CK => CLK, Q => n59721, 
                           QN => n80);
   REGS_reg_66_10_inst : DFF_X1 port map( D => n12207, CK => CLK, Q => n59720, 
                           QN => n81);
   REGS_reg_66_9_inst : DFF_X1 port map( D => n12206, CK => CLK, Q => n59719, 
                           QN => n82);
   REGS_reg_66_8_inst : DFF_X1 port map( D => n12205, CK => CLK, Q => n59718, 
                           QN => n83);
   REGS_reg_66_7_inst : DFF_X1 port map( D => n12204, CK => CLK, Q => n59729, 
                           QN => n84);
   REGS_reg_66_6_inst : DFF_X1 port map( D => n12203, CK => CLK, Q => n59728, 
                           QN => n85);
   REGS_reg_66_5_inst : DFF_X1 port map( D => n12202, CK => CLK, Q => n59727, 
                           QN => n86);
   REGS_reg_66_4_inst : DFF_X1 port map( D => n12201, CK => CLK, Q => n59726, 
                           QN => n87);
   REGS_reg_66_3_inst : DFF_X1 port map( D => n12200, CK => CLK, Q => n59725, 
                           QN => n88);
   REGS_reg_66_2_inst : DFF_X1 port map( D => n12199, CK => CLK, Q => n59724, 
                           QN => n89);
   REGS_reg_66_1_inst : DFF_X1 port map( D => n12198, CK => CLK, Q => n59723, 
                           QN => n90);
   REGS_reg_66_0_inst : DFF_X1 port map( D => n12197, CK => CLK, Q => n59722, 
                           QN => n91);
   REGS_reg_64_23_inst : DFF_X1 port map( D => n12284, CK => CLK, Q => n_1000, 
                           QN => n413);
   REGS_reg_64_22_inst : DFF_X1 port map( D => n12283, CK => CLK, Q => n_1001, 
                           QN => n414);
   REGS_reg_64_21_inst : DFF_X1 port map( D => n12282, CK => CLK, Q => n_1002, 
                           QN => n415);
   REGS_reg_64_20_inst : DFF_X1 port map( D => n12281, CK => CLK, Q => n_1003, 
                           QN => n416);
   REGS_reg_64_19_inst : DFF_X1 port map( D => n12280, CK => CLK, Q => n_1004, 
                           QN => n417);
   REGS_reg_64_18_inst : DFF_X1 port map( D => n12279, CK => CLK, Q => n_1005, 
                           QN => n418);
   REGS_reg_64_17_inst : DFF_X1 port map( D => n12278, CK => CLK, Q => n_1006, 
                           QN => n419);
   REGS_reg_64_16_inst : DFF_X1 port map( D => n12277, CK => CLK, Q => n_1007, 
                           QN => n420);
   REGS_reg_64_15_inst : DFF_X1 port map( D => n12276, CK => CLK, Q => n_1008, 
                           QN => n421);
   REGS_reg_64_14_inst : DFF_X1 port map( D => n12275, CK => CLK, Q => n_1009, 
                           QN => n422);
   REGS_reg_64_13_inst : DFF_X1 port map( D => n12274, CK => CLK, Q => n_1010, 
                           QN => n423);
   REGS_reg_64_12_inst : DFF_X1 port map( D => n12273, CK => CLK, Q => n_1011, 
                           QN => n424);
   REGS_reg_64_11_inst : DFF_X1 port map( D => n12272, CK => CLK, Q => n_1012, 
                           QN => n425);
   REGS_reg_64_10_inst : DFF_X1 port map( D => n12271, CK => CLK, Q => n_1013, 
                           QN => n426);
   REGS_reg_64_9_inst : DFF_X1 port map( D => n12270, CK => CLK, Q => n_1014, 
                           QN => n427);
   REGS_reg_64_8_inst : DFF_X1 port map( D => n12269, CK => CLK, Q => n_1015, 
                           QN => n428);
   REGS_reg_64_7_inst : DFF_X1 port map( D => n12268, CK => CLK, Q => n_1016, 
                           QN => n429);
   REGS_reg_64_6_inst : DFF_X1 port map( D => n12267, CK => CLK, Q => n_1017, 
                           QN => n430);
   REGS_reg_64_5_inst : DFF_X1 port map( D => n12266, CK => CLK, Q => n_1018, 
                           QN => n431);
   REGS_reg_64_4_inst : DFF_X1 port map( D => n12265, CK => CLK, Q => n_1019, 
                           QN => n432);
   REGS_reg_64_3_inst : DFF_X1 port map( D => n12264, CK => CLK, Q => n_1020, 
                           QN => n433);
   REGS_reg_64_2_inst : DFF_X1 port map( D => n12263, CK => CLK, Q => n_1021, 
                           QN => n434);
   REGS_reg_64_1_inst : DFF_X1 port map( D => n12262, CK => CLK, Q => n_1022, 
                           QN => n435);
   REGS_reg_64_0_inst : DFF_X1 port map( D => n12261, CK => CLK, Q => n_1023, 
                           QN => n452);
   REGS_reg_1_9_inst : DFF_X1 port map( D => n14286, CK => CLK, Q => n_1024, QN
                           => n2240);
   REGS_reg_1_8_inst : DFF_X1 port map( D => n14285, CK => CLK, Q => n_1025, QN
                           => n2241);
   REGS_reg_1_7_inst : DFF_X1 port map( D => n14284, CK => CLK, Q => n_1026, QN
                           => n2242);
   REGS_reg_1_6_inst : DFF_X1 port map( D => n14283, CK => CLK, Q => n_1027, QN
                           => n2243);
   REGS_reg_1_5_inst : DFF_X1 port map( D => n14282, CK => CLK, Q => n_1028, QN
                           => n2244);
   REGS_reg_1_4_inst : DFF_X1 port map( D => n14281, CK => CLK, Q => n_1029, QN
                           => n2245);
   REGS_reg_1_3_inst : DFF_X1 port map( D => n14280, CK => CLK, Q => n_1030, QN
                           => n2246);
   REGS_reg_1_2_inst : DFF_X1 port map( D => n14279, CK => CLK, Q => n_1031, QN
                           => n2247);
   REGS_reg_1_1_inst : DFF_X1 port map( D => n14278, CK => CLK, Q => n_1032, QN
                           => n2248);
   REGS_reg_1_0_inst : DFF_X1 port map( D => n14277, CK => CLK, Q => n_1033, QN
                           => n2076);
   REGS_reg_0_23_inst : DFF_X1 port map( D => n14332, CK => CLK, Q => n_1034, 
                           QN => n2249);
   REGS_reg_0_22_inst : DFF_X1 port map( D => n14331, CK => CLK, Q => n_1035, 
                           QN => n2250);
   REGS_reg_0_21_inst : DFF_X1 port map( D => n14330, CK => CLK, Q => n_1036, 
                           QN => n2251);
   REGS_reg_0_20_inst : DFF_X1 port map( D => n14329, CK => CLK, Q => n_1037, 
                           QN => n2252);
   REGS_reg_0_19_inst : DFF_X1 port map( D => n14328, CK => CLK, Q => n_1038, 
                           QN => n2253);
   REGS_reg_0_18_inst : DFF_X1 port map( D => n14327, CK => CLK, Q => n_1039, 
                           QN => n2254);
   REGS_reg_0_17_inst : DFF_X1 port map( D => n14326, CK => CLK, Q => n_1040, 
                           QN => n2255);
   REGS_reg_0_16_inst : DFF_X1 port map( D => n14325, CK => CLK, Q => n_1041, 
                           QN => n2256);
   REGS_reg_0_15_inst : DFF_X1 port map( D => n14324, CK => CLK, Q => n_1042, 
                           QN => n2257);
   REGS_reg_0_14_inst : DFF_X1 port map( D => n14323, CK => CLK, Q => n_1043, 
                           QN => n2258);
   REGS_reg_0_13_inst : DFF_X1 port map( D => n14322, CK => CLK, Q => n_1044, 
                           QN => n2259);
   REGS_reg_0_12_inst : DFF_X1 port map( D => n14321, CK => CLK, Q => n_1045, 
                           QN => n2260);
   REGS_reg_0_11_inst : DFF_X1 port map( D => n14320, CK => CLK, Q => n_1046, 
                           QN => n2077);
   REGS_reg_0_10_inst : DFF_X1 port map( D => n14319, CK => CLK, Q => n_1047, 
                           QN => n2261);
   REGS_reg_0_9_inst : DFF_X1 port map( D => n14318, CK => CLK, Q => n_1048, QN
                           => n2262);
   REGS_reg_0_8_inst : DFF_X1 port map( D => n14317, CK => CLK, Q => n_1049, QN
                           => n2263);
   REGS_reg_0_7_inst : DFF_X1 port map( D => n14316, CK => CLK, Q => n_1050, QN
                           => n2264);
   REGS_reg_0_6_inst : DFF_X1 port map( D => n14315, CK => CLK, Q => n_1051, QN
                           => n2265);
   REGS_reg_0_5_inst : DFF_X1 port map( D => n14314, CK => CLK, Q => n_1052, QN
                           => n2266);
   REGS_reg_0_4_inst : DFF_X1 port map( D => n14313, CK => CLK, Q => n_1053, QN
                           => n2267);
   REGS_reg_0_3_inst : DFF_X1 port map( D => n14312, CK => CLK, Q => n_1054, QN
                           => n2268);
   REGS_reg_0_2_inst : DFF_X1 port map( D => n14311, CK => CLK, Q => n_1055, QN
                           => n2269);
   REGS_reg_0_1_inst : DFF_X1 port map( D => n14310, CK => CLK, Q => n_1056, QN
                           => n2270);
   REGS_reg_0_0_inst : DFF_X1 port map( D => n14309, CK => CLK, Q => n_1057, QN
                           => n2078);
   REGS_reg_120_23_inst : DFF_X1 port map( D => n10492, CK => CLK, Q => n_1058,
                           QN => n2343);
   REGS_reg_120_22_inst : DFF_X1 port map( D => n10491, CK => CLK, Q => n_1059,
                           QN => n2344);
   REGS_reg_120_21_inst : DFF_X1 port map( D => n10490, CK => CLK, Q => n_1060,
                           QN => n2345);
   REGS_reg_120_20_inst : DFF_X1 port map( D => n10489, CK => CLK, Q => n_1061,
                           QN => n2346);
   REGS_reg_120_19_inst : DFF_X1 port map( D => n10488, CK => CLK, Q => n_1062,
                           QN => n2347);
   REGS_reg_120_18_inst : DFF_X1 port map( D => n10487, CK => CLK, Q => n_1063,
                           QN => n2348);
   REGS_reg_120_17_inst : DFF_X1 port map( D => n10486, CK => CLK, Q => n_1064,
                           QN => n2349);
   REGS_reg_120_16_inst : DFF_X1 port map( D => n10485, CK => CLK, Q => n_1065,
                           QN => n2350);
   REGS_reg_120_15_inst : DFF_X1 port map( D => n10484, CK => CLK, Q => n_1066,
                           QN => n2351);
   REGS_reg_120_14_inst : DFF_X1 port map( D => n10483, CK => CLK, Q => n_1067,
                           QN => n2352);
   REGS_reg_120_13_inst : DFF_X1 port map( D => n10482, CK => CLK, Q => n_1068,
                           QN => n2353);
   REGS_reg_120_12_inst : DFF_X1 port map( D => n10481, CK => CLK, Q => n_1069,
                           QN => n2354);
   REGS_reg_120_11_inst : DFF_X1 port map( D => n10480, CK => CLK, Q => n_1070,
                           QN => n2355);
   REGS_reg_120_10_inst : DFF_X1 port map( D => n10479, CK => CLK, Q => n_1071,
                           QN => n2356);
   REGS_reg_120_9_inst : DFF_X1 port map( D => n10478, CK => CLK, Q => n_1072, 
                           QN => n2357);
   REGS_reg_120_8_inst : DFF_X1 port map( D => n10477, CK => CLK, Q => n_1073, 
                           QN => n2358);
   REGS_reg_120_7_inst : DFF_X1 port map( D => n10476, CK => CLK, Q => n_1074, 
                           QN => n2359);
   REGS_reg_120_6_inst : DFF_X1 port map( D => n10475, CK => CLK, Q => n_1075, 
                           QN => n2360);
   REGS_reg_120_5_inst : DFF_X1 port map( D => n10474, CK => CLK, Q => n_1076, 
                           QN => n2361);
   REGS_reg_120_4_inst : DFF_X1 port map( D => n10473, CK => CLK, Q => n_1077, 
                           QN => n2362);
   REGS_reg_120_3_inst : DFF_X1 port map( D => n10472, CK => CLK, Q => n_1078, 
                           QN => n2363);
   REGS_reg_120_2_inst : DFF_X1 port map( D => n10471, CK => CLK, Q => n_1079, 
                           QN => n2364);
   REGS_reg_120_1_inst : DFF_X1 port map( D => n10470, CK => CLK, Q => n_1080, 
                           QN => n2365);
   REGS_reg_120_0_inst : DFF_X1 port map( D => n10469, CK => CLK, Q => n_1081, 
                           QN => n2366);
   REGS_reg_119_23_inst : DFF_X1 port map( D => n10524, CK => CLK, Q => n_1082,
                           QN => n2367);
   REGS_reg_119_22_inst : DFF_X1 port map( D => n10523, CK => CLK, Q => n_1083,
                           QN => n2368);
   REGS_reg_119_21_inst : DFF_X1 port map( D => n10522, CK => CLK, Q => n_1084,
                           QN => n2369);
   REGS_reg_119_20_inst : DFF_X1 port map( D => n10521, CK => CLK, Q => n_1085,
                           QN => n2370);
   REGS_reg_119_19_inst : DFF_X1 port map( D => n10520, CK => CLK, Q => n_1086,
                           QN => n2371);
   REGS_reg_119_18_inst : DFF_X1 port map( D => n10519, CK => CLK, Q => n_1087,
                           QN => n2372);
   REGS_reg_119_17_inst : DFF_X1 port map( D => n10518, CK => CLK, Q => n_1088,
                           QN => n2373);
   REGS_reg_119_16_inst : DFF_X1 port map( D => n10517, CK => CLK, Q => n_1089,
                           QN => n2374);
   REGS_reg_119_15_inst : DFF_X1 port map( D => n10516, CK => CLK, Q => n_1090,
                           QN => n2375);
   REGS_reg_119_14_inst : DFF_X1 port map( D => n10515, CK => CLK, Q => n_1091,
                           QN => n2376);
   REGS_reg_119_13_inst : DFF_X1 port map( D => n10514, CK => CLK, Q => n_1092,
                           QN => n2377);
   REGS_reg_119_12_inst : DFF_X1 port map( D => n10513, CK => CLK, Q => n_1093,
                           QN => n2378);
   REGS_reg_119_11_inst : DFF_X1 port map( D => n10512, CK => CLK, Q => n_1094,
                           QN => n2379);
   REGS_reg_119_10_inst : DFF_X1 port map( D => n10511, CK => CLK, Q => n_1095,
                           QN => n2380);
   REGS_reg_119_9_inst : DFF_X1 port map( D => n10510, CK => CLK, Q => n_1096, 
                           QN => n2381);
   REGS_reg_119_8_inst : DFF_X1 port map( D => n10509, CK => CLK, Q => n_1097, 
                           QN => n2382);
   REGS_reg_119_7_inst : DFF_X1 port map( D => n10508, CK => CLK, Q => n_1098, 
                           QN => n2383);
   REGS_reg_119_6_inst : DFF_X1 port map( D => n10507, CK => CLK, Q => n_1099, 
                           QN => n2384);
   REGS_reg_119_5_inst : DFF_X1 port map( D => n10506, CK => CLK, Q => n_1100, 
                           QN => n2385);
   REGS_reg_119_4_inst : DFF_X1 port map( D => n10505, CK => CLK, Q => n_1101, 
                           QN => n2386);
   REGS_reg_119_3_inst : DFF_X1 port map( D => n10504, CK => CLK, Q => n_1102, 
                           QN => n2387);
   REGS_reg_119_2_inst : DFF_X1 port map( D => n10503, CK => CLK, Q => n_1103, 
                           QN => n2388);
   REGS_reg_119_1_inst : DFF_X1 port map( D => n10502, CK => CLK, Q => n_1104, 
                           QN => n2389);
   REGS_reg_119_0_inst : DFF_X1 port map( D => n10501, CK => CLK, Q => n_1105, 
                           QN => n2390);
   REGS_reg_109_23_inst : DFF_X1 port map( D => n10844, CK => CLK, Q => n_1106,
                           QN => n2487);
   REGS_reg_109_22_inst : DFF_X1 port map( D => n10843, CK => CLK, Q => n_1107,
                           QN => n2488);
   REGS_reg_109_21_inst : DFF_X1 port map( D => n10842, CK => CLK, Q => n_1108,
                           QN => n2489);
   REGS_reg_109_20_inst : DFF_X1 port map( D => n10841, CK => CLK, Q => n_1109,
                           QN => n2490);
   REGS_reg_109_19_inst : DFF_X1 port map( D => n10840, CK => CLK, Q => n_1110,
                           QN => n2491);
   REGS_reg_109_18_inst : DFF_X1 port map( D => n10839, CK => CLK, Q => n_1111,
                           QN => n2492);
   REGS_reg_109_17_inst : DFF_X1 port map( D => n10838, CK => CLK, Q => n_1112,
                           QN => n2493);
   REGS_reg_109_16_inst : DFF_X1 port map( D => n10837, CK => CLK, Q => n_1113,
                           QN => n2494);
   REGS_reg_109_15_inst : DFF_X1 port map( D => n10836, CK => CLK, Q => n_1114,
                           QN => n2495);
   REGS_reg_109_14_inst : DFF_X1 port map( D => n10835, CK => CLK, Q => n_1115,
                           QN => n2496);
   REGS_reg_109_13_inst : DFF_X1 port map( D => n10834, CK => CLK, Q => n_1116,
                           QN => n2497);
   REGS_reg_109_12_inst : DFF_X1 port map( D => n10833, CK => CLK, Q => n_1117,
                           QN => n2498);
   REGS_reg_109_11_inst : DFF_X1 port map( D => n10832, CK => CLK, Q => n_1118,
                           QN => n2499);
   REGS_reg_109_10_inst : DFF_X1 port map( D => n10831, CK => CLK, Q => n_1119,
                           QN => n2500);
   REGS_reg_109_9_inst : DFF_X1 port map( D => n10830, CK => CLK, Q => n_1120, 
                           QN => n2501);
   REGS_reg_109_8_inst : DFF_X1 port map( D => n10829, CK => CLK, Q => n_1121, 
                           QN => n2502);
   REGS_reg_109_7_inst : DFF_X1 port map( D => n10828, CK => CLK, Q => n_1122, 
                           QN => n2503);
   REGS_reg_109_6_inst : DFF_X1 port map( D => n10827, CK => CLK, Q => n_1123, 
                           QN => n2504);
   REGS_reg_109_5_inst : DFF_X1 port map( D => n10826, CK => CLK, Q => n_1124, 
                           QN => n2505);
   REGS_reg_109_4_inst : DFF_X1 port map( D => n10825, CK => CLK, Q => n_1125, 
                           QN => n2506);
   REGS_reg_109_3_inst : DFF_X1 port map( D => n10824, CK => CLK, Q => n_1126, 
                           QN => n2507);
   REGS_reg_109_2_inst : DFF_X1 port map( D => n10823, CK => CLK, Q => n_1127, 
                           QN => n2508);
   REGS_reg_109_1_inst : DFF_X1 port map( D => n10822, CK => CLK, Q => n_1128, 
                           QN => n2509);
   REGS_reg_109_0_inst : DFF_X1 port map( D => n10821, CK => CLK, Q => n_1129, 
                           QN => n2510);
   REGS_reg_108_23_inst : DFF_X1 port map( D => n10876, CK => CLK, Q => n_1130,
                           QN => n3967);
   REGS_reg_108_22_inst : DFF_X1 port map( D => n10875, CK => CLK, Q => n_1131,
                           QN => n3968);
   REGS_reg_108_21_inst : DFF_X1 port map( D => n10874, CK => CLK, Q => n_1132,
                           QN => n3969);
   REGS_reg_108_20_inst : DFF_X1 port map( D => n10873, CK => CLK, Q => n_1133,
                           QN => n3970);
   REGS_reg_108_19_inst : DFF_X1 port map( D => n10872, CK => CLK, Q => n_1134,
                           QN => n3971);
   REGS_reg_108_18_inst : DFF_X1 port map( D => n10871, CK => CLK, Q => n_1135,
                           QN => n3972);
   REGS_reg_108_17_inst : DFF_X1 port map( D => n10870, CK => CLK, Q => n_1136,
                           QN => n3973);
   REGS_reg_108_16_inst : DFF_X1 port map( D => n10869, CK => CLK, Q => n_1137,
                           QN => n3974);
   REGS_reg_108_15_inst : DFF_X1 port map( D => n10868, CK => CLK, Q => n_1138,
                           QN => n3975);
   REGS_reg_108_14_inst : DFF_X1 port map( D => n10867, CK => CLK, Q => n_1139,
                           QN => n3976);
   REGS_reg_108_13_inst : DFF_X1 port map( D => n10866, CK => CLK, Q => n_1140,
                           QN => n3977);
   REGS_reg_108_12_inst : DFF_X1 port map( D => n10865, CK => CLK, Q => n_1141,
                           QN => n3978);
   REGS_reg_108_11_inst : DFF_X1 port map( D => n10864, CK => CLK, Q => n_1142,
                           QN => n3979);
   REGS_reg_108_10_inst : DFF_X1 port map( D => n10863, CK => CLK, Q => n_1143,
                           QN => n3980);
   REGS_reg_108_9_inst : DFF_X1 port map( D => n10862, CK => CLK, Q => n_1144, 
                           QN => n3981);
   REGS_reg_108_8_inst : DFF_X1 port map( D => n10861, CK => CLK, Q => n_1145, 
                           QN => n3982);
   REGS_reg_108_7_inst : DFF_X1 port map( D => n10860, CK => CLK, Q => n_1146, 
                           QN => n3983);
   REGS_reg_108_6_inst : DFF_X1 port map( D => n10859, CK => CLK, Q => n_1147, 
                           QN => n3984);
   REGS_reg_108_5_inst : DFF_X1 port map( D => n10858, CK => CLK, Q => n_1148, 
                           QN => n3985);
   REGS_reg_108_4_inst : DFF_X1 port map( D => n10857, CK => CLK, Q => n_1149, 
                           QN => n3986);
   REGS_reg_108_3_inst : DFF_X1 port map( D => n10856, CK => CLK, Q => n_1150, 
                           QN => n3987);
   REGS_reg_108_2_inst : DFF_X1 port map( D => n10855, CK => CLK, Q => n_1151, 
                           QN => n3988);
   REGS_reg_108_1_inst : DFF_X1 port map( D => n10854, CK => CLK, Q => n_1152, 
                           QN => n3989);
   REGS_reg_108_0_inst : DFF_X1 port map( D => n10853, CK => CLK, Q => n_1153, 
                           QN => n3990);
   REGS_reg_134_10_inst : DFF_X1 port map( D => n10031, CK => CLK, Q => n59675,
                           QN => n92);
   REGS_reg_134_9_inst : DFF_X1 port map( D => n10030, CK => CLK, Q => n59674, 
                           QN => n93);
   REGS_reg_134_8_inst : DFF_X1 port map( D => n10029, CK => CLK, Q => n59673, 
                           QN => n94);
   REGS_reg_134_7_inst : DFF_X1 port map( D => n10028, CK => CLK, Q => n59680, 
                           QN => n95);
   REGS_reg_134_6_inst : DFF_X1 port map( D => n10027, CK => CLK, Q => n59679, 
                           QN => n96);
   REGS_reg_134_5_inst : DFF_X1 port map( D => n10026, CK => CLK, Q => n59678, 
                           QN => n97);
   REGS_reg_134_4_inst : DFF_X1 port map( D => n10025, CK => CLK, Q => n59677, 
                           QN => n98);
   REGS_reg_134_3_inst : DFF_X1 port map( D => n10024, CK => CLK, Q => n59676, 
                           QN => n99);
   REGS_reg_134_11_inst : DFF_X1 port map( D => n10032, CK => CLK, Q => n59681,
                           QN => n54444);
   REGS_reg_134_18_inst : DFF_X1 port map( D => n10039, CK => CLK, Q => n59687,
                           QN => n54445);
   REGS_reg_134_17_inst : DFF_X1 port map( D => n10038, CK => CLK, Q => n59686,
                           QN => n54446);
   REGS_reg_134_16_inst : DFF_X1 port map( D => n10037, CK => CLK, Q => n59685,
                           QN => n54447);
   REGS_reg_134_15_inst : DFF_X1 port map( D => n10036, CK => CLK, Q => n59684,
                           QN => n54448);
   REGS_reg_134_14_inst : DFF_X1 port map( D => n10035, CK => CLK, Q => n59683,
                           QN => n54449);
   REGS_reg_134_13_inst : DFF_X1 port map( D => n10034, CK => CLK, Q => n59682,
                           QN => n54450);
   REGS_reg_134_12_inst : DFF_X1 port map( D => n10033, CK => CLK, Q => n59688,
                           QN => n54451);
   OUT1_reg_0_inst : DFF_X1 port map( D => n9957, CK => CLK, Q => OUT1(0), QN 
                           => n9314);
   REGS_reg_133_31_inst : DFF_X1 port map( D => n10084, CK => CLK, Q => n52236,
                           QN => n1);
   REGS_reg_133_30_inst : DFF_X1 port map( D => n10083, CK => CLK, Q => n52237,
                           QN => n2);
   REGS_reg_133_29_inst : DFF_X1 port map( D => n10082, CK => CLK, Q => n52238,
                           QN => n3);
   REGS_reg_132_31_inst : DFF_X1 port map( D => n10116, CK => CLK, Q => n_1154,
                           QN => n4);
   REGS_reg_132_30_inst : DFF_X1 port map( D => n10115, CK => CLK, Q => n_1155,
                           QN => n5);
   REGS_reg_132_29_inst : DFF_X1 port map( D => n10114, CK => CLK, Q => n_1156,
                           QN => n6);
   REGS_reg_132_28_inst : DFF_X1 port map( D => n10113, CK => CLK, Q => n_1157,
                           QN => n7);
   REGS_reg_132_27_inst : DFF_X1 port map( D => n10112, CK => CLK, Q => n_1158,
                           QN => n8);
   REGS_reg_132_26_inst : DFF_X1 port map( D => n10111, CK => CLK, Q => n_1159,
                           QN => n9);
   REGS_reg_132_25_inst : DFF_X1 port map( D => n10110, CK => CLK, Q => n_1160,
                           QN => n10);
   REGS_reg_132_24_inst : DFF_X1 port map( D => n10109, CK => CLK, Q => n_1161,
                           QN => n11);
   REGS_reg_131_31_inst : DFF_X1 port map( D => n10148, CK => CLK, Q => n_1162,
                           QN => n12);
   REGS_reg_131_30_inst : DFF_X1 port map( D => n10147, CK => CLK, Q => n_1163,
                           QN => n13);
   REGS_reg_131_29_inst : DFF_X1 port map( D => n10146, CK => CLK, Q => n_1164,
                           QN => n14);
   REGS_reg_131_28_inst : DFF_X1 port map( D => n10145, CK => CLK, Q => n_1165,
                           QN => n15);
   REGS_reg_131_27_inst : DFF_X1 port map( D => n10144, CK => CLK, Q => n_1166,
                           QN => n16);
   REGS_reg_131_26_inst : DFF_X1 port map( D => n10143, CK => CLK, Q => n_1167,
                           QN => n17);
   REGS_reg_131_25_inst : DFF_X1 port map( D => n10142, CK => CLK, Q => n_1168,
                           QN => n18);
   REGS_reg_131_24_inst : DFF_X1 port map( D => n10141, CK => CLK, Q => n_1169,
                           QN => n19);
   REGS_reg_130_31_inst : DFF_X1 port map( D => n10180, CK => CLK, Q => n_1170,
                           QN => n20);
   REGS_reg_130_30_inst : DFF_X1 port map( D => n10179, CK => CLK, Q => n_1171,
                           QN => n21);
   REGS_reg_130_29_inst : DFF_X1 port map( D => n10178, CK => CLK, Q => n_1172,
                           QN => n22);
   REGS_reg_130_28_inst : DFF_X1 port map( D => n10177, CK => CLK, Q => n_1173,
                           QN => n23);
   REGS_reg_130_27_inst : DFF_X1 port map( D => n10176, CK => CLK, Q => n_1174,
                           QN => n24);
   REGS_reg_130_26_inst : DFF_X1 port map( D => n10175, CK => CLK, Q => n_1175,
                           QN => n25);
   REGS_reg_130_25_inst : DFF_X1 port map( D => n10174, CK => CLK, Q => n_1176,
                           QN => n26);
   REGS_reg_130_24_inst : DFF_X1 port map( D => n10173, CK => CLK, Q => n_1177,
                           QN => n27);
   REGS_reg_129_31_inst : DFF_X1 port map( D => n10212, CK => CLK, Q => n_1178,
                           QN => n28);
   REGS_reg_129_30_inst : DFF_X1 port map( D => n10211, CK => CLK, Q => n_1179,
                           QN => n29);
   REGS_reg_129_29_inst : DFF_X1 port map( D => n10210, CK => CLK, Q => n_1180,
                           QN => n30);
   REGS_reg_129_28_inst : DFF_X1 port map( D => n10209, CK => CLK, Q => n_1181,
                           QN => n31);
   REGS_reg_129_27_inst : DFF_X1 port map( D => n10208, CK => CLK, Q => n_1182,
                           QN => n32);
   REGS_reg_129_26_inst : DFF_X1 port map( D => n10207, CK => CLK, Q => n_1183,
                           QN => n33);
   REGS_reg_129_25_inst : DFF_X1 port map( D => n10206, CK => CLK, Q => n_1184,
                           QN => n34);
   REGS_reg_129_24_inst : DFF_X1 port map( D => n10205, CK => CLK, Q => n_1185,
                           QN => n35);
   REGS_reg_128_31_inst : DFF_X1 port map( D => n10244, CK => CLK, Q => n16476,
                           QN => n3940);
   REGS_reg_128_30_inst : DFF_X1 port map( D => n10243, CK => CLK, Q => n16475,
                           QN => n3941);
   REGS_reg_128_29_inst : DFF_X1 port map( D => n10242, CK => CLK, Q => n16474,
                           QN => n3942);
   REGS_reg_128_28_inst : DFF_X1 port map( D => n10241, CK => CLK, Q => n16473,
                           QN => n3943);
   REGS_reg_128_27_inst : DFF_X1 port map( D => n10240, CK => CLK, Q => n16472,
                           QN => n3944);
   REGS_reg_128_26_inst : DFF_X1 port map( D => n10239, CK => CLK, Q => n16471,
                           QN => n3945);
   REGS_reg_128_25_inst : DFF_X1 port map( D => n10238, CK => CLK, Q => n16470,
                           QN => n3946);
   REGS_reg_128_24_inst : DFF_X1 port map( D => n10237, CK => CLK, Q => n16469,
                           QN => n3947);
   REGS_reg_62_31_inst : DFF_X1 port map( D => n12356, CK => CLK, Q => n506, QN
                           => n4180);
   REGS_reg_62_30_inst : DFF_X1 port map( D => n12355, CK => CLK, Q => n507, QN
                           => n4181);
   REGS_reg_62_29_inst : DFF_X1 port map( D => n12354, CK => CLK, Q => n508, QN
                           => n4182);
   REGS_reg_62_28_inst : DFF_X1 port map( D => n12353, CK => CLK, Q => n509, QN
                           => n4183);
   REGS_reg_62_27_inst : DFF_X1 port map( D => n12352, CK => CLK, Q => n510, QN
                           => n4184);
   REGS_reg_62_26_inst : DFF_X1 port map( D => n12351, CK => CLK, Q => n511, QN
                           => n4185);
   REGS_reg_62_25_inst : DFF_X1 port map( D => n12350, CK => CLK, Q => n512, QN
                           => n4186);
   REGS_reg_62_24_inst : DFF_X1 port map( D => n12349, CK => CLK, Q => n513, QN
                           => n4187);
   REGS_reg_61_31_inst : DFF_X1 port map( D => n12388, CK => CLK, Q => n514, QN
                           => n4188);
   REGS_reg_61_30_inst : DFF_X1 port map( D => n12387, CK => CLK, Q => n515, QN
                           => n4189);
   REGS_reg_61_29_inst : DFF_X1 port map( D => n12386, CK => CLK, Q => n516, QN
                           => n4190);
   REGS_reg_61_28_inst : DFF_X1 port map( D => n12385, CK => CLK, Q => n517, QN
                           => n4191);
   REGS_reg_61_27_inst : DFF_X1 port map( D => n12384, CK => CLK, Q => n518, QN
                           => n4192);
   REGS_reg_61_26_inst : DFF_X1 port map( D => n12383, CK => CLK, Q => n520, QN
                           => n4193);
   REGS_reg_61_25_inst : DFF_X1 port map( D => n12382, CK => CLK, Q => n521, QN
                           => n4194);
   REGS_reg_61_24_inst : DFF_X1 port map( D => n12381, CK => CLK, Q => n522, QN
                           => n4195);
   REGS_reg_60_31_inst : DFF_X1 port map( D => n12420, CK => CLK, Q => n52268, 
                           QN => n487);
   REGS_reg_60_30_inst : DFF_X1 port map( D => n12419, CK => CLK, Q => n52269, 
                           QN => n488);
   REGS_reg_60_29_inst : DFF_X1 port map( D => n12418, CK => CLK, Q => n52270, 
                           QN => n489);
   REGS_reg_60_28_inst : DFF_X1 port map( D => n12417, CK => CLK, Q => n52271, 
                           QN => n490);
   REGS_reg_60_27_inst : DFF_X1 port map( D => n12416, CK => CLK, Q => n52272, 
                           QN => n491);
   REGS_reg_60_26_inst : DFF_X1 port map( D => n12415, CK => CLK, Q => n52273, 
                           QN => n492);
   REGS_reg_60_25_inst : DFF_X1 port map( D => n12414, CK => CLK, Q => n52274, 
                           QN => n493);
   REGS_reg_60_24_inst : DFF_X1 port map( D => n12413, CK => CLK, Q => n52275, 
                           QN => n494);
   REGS_reg_59_31_inst : DFF_X1 port map( D => n12452, CK => CLK, Q => n_1186, 
                           QN => n495);
   REGS_reg_59_30_inst : DFF_X1 port map( D => n12451, CK => CLK, Q => n_1187, 
                           QN => n496);
   REGS_reg_59_29_inst : DFF_X1 port map( D => n12450, CK => CLK, Q => n_1188, 
                           QN => n497);
   REGS_reg_59_28_inst : DFF_X1 port map( D => n12449, CK => CLK, Q => n_1189, 
                           QN => n498);
   REGS_reg_59_27_inst : DFF_X1 port map( D => n12448, CK => CLK, Q => n_1190, 
                           QN => n499);
   REGS_reg_59_26_inst : DFF_X1 port map( D => n12447, CK => CLK, Q => n_1191, 
                           QN => n560);
   REGS_reg_59_25_inst : DFF_X1 port map( D => n12446, CK => CLK, Q => n_1192, 
                           QN => n561);
   REGS_reg_59_24_inst : DFF_X1 port map( D => n12445, CK => CLK, Q => n_1193, 
                           QN => n562);
   REGS_reg_58_31_inst : DFF_X1 port map( D => n12484, CK => CLK, Q => n15611, 
                           QN => n563);
   REGS_reg_58_30_inst : DFF_X1 port map( D => n12483, CK => CLK, Q => n15599, 
                           QN => n564);
   REGS_reg_58_29_inst : DFF_X1 port map( D => n12482, CK => CLK, Q => n15597, 
                           QN => n565);
   REGS_reg_58_28_inst : DFF_X1 port map( D => n12481, CK => CLK, Q => n15595, 
                           QN => n566);
   REGS_reg_58_27_inst : DFF_X1 port map( D => n12480, CK => CLK, Q => n15593, 
                           QN => n567);
   REGS_reg_58_26_inst : DFF_X1 port map( D => n12479, CK => CLK, Q => n15591, 
                           QN => n760);
   REGS_reg_58_25_inst : DFF_X1 port map( D => n12478, CK => CLK, Q => n15589, 
                           QN => n761);
   REGS_reg_58_24_inst : DFF_X1 port map( D => n12477, CK => CLK, Q => n15587, 
                           QN => n762);
   REGS_reg_57_31_inst : DFF_X1 port map( D => n12516, CK => CLK, Q => n15612, 
                           QN => n763);
   REGS_reg_57_30_inst : DFF_X1 port map( D => n12515, CK => CLK, Q => n15600, 
                           QN => n764);
   REGS_reg_57_29_inst : DFF_X1 port map( D => n12514, CK => CLK, Q => n15598, 
                           QN => n765);
   REGS_reg_57_28_inst : DFF_X1 port map( D => n12513, CK => CLK, Q => n15596, 
                           QN => n766);
   REGS_reg_57_27_inst : DFF_X1 port map( D => n12512, CK => CLK, Q => n15594, 
                           QN => n767);
   REGS_reg_57_26_inst : DFF_X1 port map( D => n12511, CK => CLK, Q => n15592, 
                           QN => n768);
   REGS_reg_57_25_inst : DFF_X1 port map( D => n12510, CK => CLK, Q => n15590, 
                           QN => n769);
   REGS_reg_57_24_inst : DFF_X1 port map( D => n12509, CK => CLK, Q => n15588, 
                           QN => n770);
   REGS_reg_56_31_inst : DFF_X1 port map( D => n12548, CK => CLK, Q => n523, QN
                           => n4196);
   REGS_reg_56_30_inst : DFF_X1 port map( D => n12547, CK => CLK, Q => n524, QN
                           => n4197);
   REGS_reg_56_29_inst : DFF_X1 port map( D => n12546, CK => CLK, Q => n525, QN
                           => n4198);
   REGS_reg_56_28_inst : DFF_X1 port map( D => n12545, CK => CLK, Q => n526, QN
                           => n4199);
   REGS_reg_56_27_inst : DFF_X1 port map( D => n12544, CK => CLK, Q => n527, QN
                           => n4200);
   REGS_reg_56_26_inst : DFF_X1 port map( D => n12543, CK => CLK, Q => n528, QN
                           => n4201);
   REGS_reg_56_25_inst : DFF_X1 port map( D => n12542, CK => CLK, Q => n529, QN
                           => n4202);
   REGS_reg_56_24_inst : DFF_X1 port map( D => n12541, CK => CLK, Q => n530, QN
                           => n4203);
   REGS_reg_55_31_inst : DFF_X1 port map( D => n12580, CK => CLK, Q => n531, QN
                           => n4204);
   REGS_reg_55_30_inst : DFF_X1 port map( D => n12579, CK => CLK, Q => n532, QN
                           => n4205);
   REGS_reg_55_29_inst : DFF_X1 port map( D => n12578, CK => CLK, Q => n533, QN
                           => n4206);
   REGS_reg_55_28_inst : DFF_X1 port map( D => n12577, CK => CLK, Q => n534, QN
                           => n4207);
   REGS_reg_55_27_inst : DFF_X1 port map( D => n12576, CK => CLK, Q => n535, QN
                           => n4208);
   REGS_reg_55_26_inst : DFF_X1 port map( D => n12575, CK => CLK, Q => n536, QN
                           => n4209);
   REGS_reg_55_25_inst : DFF_X1 port map( D => n12574, CK => CLK, Q => n537, QN
                           => n4210);
   REGS_reg_55_24_inst : DFF_X1 port map( D => n12573, CK => CLK, Q => n538, QN
                           => n4211);
   REGS_reg_53_31_inst : DFF_X1 port map( D => n12644, CK => CLK, Q => n547, QN
                           => n4212);
   REGS_reg_53_30_inst : DFF_X1 port map( D => n12643, CK => CLK, Q => n548, QN
                           => n4213);
   REGS_reg_53_29_inst : DFF_X1 port map( D => n12642, CK => CLK, Q => n549, QN
                           => n4214);
   REGS_reg_53_28_inst : DFF_X1 port map( D => n12641, CK => CLK, Q => n550, QN
                           => n4215);
   REGS_reg_53_27_inst : DFF_X1 port map( D => n12640, CK => CLK, Q => n551, QN
                           => n4216);
   REGS_reg_53_26_inst : DFF_X1 port map( D => n12639, CK => CLK, Q => n552, QN
                           => n4217);
   REGS_reg_53_25_inst : DFF_X1 port map( D => n12638, CK => CLK, Q => n553, QN
                           => n4218);
   REGS_reg_53_24_inst : DFF_X1 port map( D => n12637, CK => CLK, Q => n554, QN
                           => n4219);
   REGS_reg_52_31_inst : DFF_X1 port map( D => n12676, CK => CLK, Q => n_1194, 
                           QN => n787);
   REGS_reg_52_30_inst : DFF_X1 port map( D => n12675, CK => CLK, Q => n_1195, 
                           QN => n788);
   REGS_reg_52_29_inst : DFF_X1 port map( D => n12674, CK => CLK, Q => n_1196, 
                           QN => n789);
   REGS_reg_52_28_inst : DFF_X1 port map( D => n12673, CK => CLK, Q => n_1197, 
                           QN => n790);
   REGS_reg_52_27_inst : DFF_X1 port map( D => n12672, CK => CLK, Q => n_1198, 
                           QN => n791);
   REGS_reg_52_26_inst : DFF_X1 port map( D => n12671, CK => CLK, Q => n_1199, 
                           QN => n792);
   REGS_reg_52_25_inst : DFF_X1 port map( D => n12670, CK => CLK, Q => n_1200, 
                           QN => n793);
   REGS_reg_52_24_inst : DFF_X1 port map( D => n12669, CK => CLK, Q => n_1201, 
                           QN => n794);
   REGS_reg_51_31_inst : DFF_X1 port map( D => n12708, CK => CLK, Q => n_1202, 
                           QN => n795);
   REGS_reg_51_30_inst : DFF_X1 port map( D => n12707, CK => CLK, Q => n_1203, 
                           QN => n796);
   REGS_reg_51_29_inst : DFF_X1 port map( D => n12706, CK => CLK, Q => n_1204, 
                           QN => n797);
   REGS_reg_51_28_inst : DFF_X1 port map( D => n12705, CK => CLK, Q => n_1205, 
                           QN => n798);
   REGS_reg_51_27_inst : DFF_X1 port map( D => n12704, CK => CLK, Q => n_1206, 
                           QN => n799);
   REGS_reg_51_26_inst : DFF_X1 port map( D => n12703, CK => CLK, Q => n_1207, 
                           QN => n800);
   REGS_reg_51_25_inst : DFF_X1 port map( D => n12702, CK => CLK, Q => n_1208, 
                           QN => n801);
   REGS_reg_51_24_inst : DFF_X1 port map( D => n12701, CK => CLK, Q => n_1209, 
                           QN => n802);
   REGS_reg_50_31_inst : DFF_X1 port map( D => n12740, CK => CLK, Q => n52308, 
                           QN => n803);
   REGS_reg_50_30_inst : DFF_X1 port map( D => n12739, CK => CLK, Q => n52309, 
                           QN => n804);
   REGS_reg_50_29_inst : DFF_X1 port map( D => n12738, CK => CLK, Q => n52310, 
                           QN => n805);
   REGS_reg_50_28_inst : DFF_X1 port map( D => n12737, CK => CLK, Q => n52311, 
                           QN => n806);
   REGS_reg_50_27_inst : DFF_X1 port map( D => n12736, CK => CLK, Q => n52312, 
                           QN => n807);
   REGS_reg_50_26_inst : DFF_X1 port map( D => n12735, CK => CLK, Q => n52313, 
                           QN => n808);
   REGS_reg_50_25_inst : DFF_X1 port map( D => n12734, CK => CLK, Q => n52314, 
                           QN => n809);
   REGS_reg_50_24_inst : DFF_X1 port map( D => n12733, CK => CLK, Q => n52315, 
                           QN => n810);
   REGS_reg_49_31_inst : DFF_X1 port map( D => n12772, CK => CLK, Q => n52316, 
                           QN => n811);
   REGS_reg_49_30_inst : DFF_X1 port map( D => n12771, CK => CLK, Q => n52317, 
                           QN => n812);
   REGS_reg_49_29_inst : DFF_X1 port map( D => n12770, CK => CLK, Q => n52318, 
                           QN => n813);
   REGS_reg_49_28_inst : DFF_X1 port map( D => n12769, CK => CLK, Q => n52319, 
                           QN => n814);
   REGS_reg_49_27_inst : DFF_X1 port map( D => n12768, CK => CLK, Q => n52320, 
                           QN => n815);
   REGS_reg_49_26_inst : DFF_X1 port map( D => n12767, CK => CLK, Q => n52321, 
                           QN => n972);
   REGS_reg_49_25_inst : DFF_X1 port map( D => n12766, CK => CLK, Q => n52322, 
                           QN => n973);
   REGS_reg_49_24_inst : DFF_X1 port map( D => n12765, CK => CLK, Q => n52323, 
                           QN => n974);
   REGS_reg_48_31_inst : DFF_X1 port map( D => n12804, CK => CLK, Q => n52324, 
                           QN => n975);
   REGS_reg_48_30_inst : DFF_X1 port map( D => n12803, CK => CLK, Q => n52325, 
                           QN => n976);
   REGS_reg_48_29_inst : DFF_X1 port map( D => n12802, CK => CLK, Q => n52326, 
                           QN => n977);
   REGS_reg_48_28_inst : DFF_X1 port map( D => n12801, CK => CLK, Q => n52327, 
                           QN => n978);
   REGS_reg_48_27_inst : DFF_X1 port map( D => n12800, CK => CLK, Q => n52328, 
                           QN => n979);
   REGS_reg_48_26_inst : DFF_X1 port map( D => n12799, CK => CLK, Q => n52329, 
                           QN => n980);
   REGS_reg_48_25_inst : DFF_X1 port map( D => n12798, CK => CLK, Q => n52330, 
                           QN => n981);
   REGS_reg_48_24_inst : DFF_X1 port map( D => n12797, CK => CLK, Q => n52331, 
                           QN => n982);
   REGS_reg_47_31_inst : DFF_X1 port map( D => n12836, CK => CLK, Q => n16468, 
                           QN => n4220);
   REGS_reg_47_30_inst : DFF_X1 port map( D => n12835, CK => CLK, Q => n16467, 
                           QN => n4221);
   REGS_reg_47_29_inst : DFF_X1 port map( D => n12834, CK => CLK, Q => n16466, 
                           QN => n4222);
   REGS_reg_47_28_inst : DFF_X1 port map( D => n12833, CK => CLK, Q => n16465, 
                           QN => n4223);
   REGS_reg_47_27_inst : DFF_X1 port map( D => n12832, CK => CLK, Q => n16464, 
                           QN => n4224);
   REGS_reg_47_26_inst : DFF_X1 port map( D => n12831, CK => CLK, Q => n16463, 
                           QN => n4225);
   REGS_reg_47_25_inst : DFF_X1 port map( D => n12830, CK => CLK, Q => n16462, 
                           QN => n4226);
   REGS_reg_47_24_inst : DFF_X1 port map( D => n12829, CK => CLK, Q => n16461, 
                           QN => n4227);
   REGS_reg_46_31_inst : DFF_X1 port map( D => n12868, CK => CLK, Q => n16460, 
                           QN => n4228);
   REGS_reg_46_30_inst : DFF_X1 port map( D => n12867, CK => CLK, Q => n16459, 
                           QN => n4229);
   REGS_reg_46_29_inst : DFF_X1 port map( D => n12866, CK => CLK, Q => n16458, 
                           QN => n4230);
   REGS_reg_46_28_inst : DFF_X1 port map( D => n12865, CK => CLK, Q => n16457, 
                           QN => n4231);
   REGS_reg_46_27_inst : DFF_X1 port map( D => n12864, CK => CLK, Q => n16456, 
                           QN => n4232);
   REGS_reg_46_26_inst : DFF_X1 port map( D => n12863, CK => CLK, Q => n16455, 
                           QN => n4233);
   REGS_reg_46_25_inst : DFF_X1 port map( D => n12862, CK => CLK, Q => n16454, 
                           QN => n4234);
   REGS_reg_46_24_inst : DFF_X1 port map( D => n12861, CK => CLK, Q => n16453, 
                           QN => n4235);
   REGS_reg_45_31_inst : DFF_X1 port map( D => n12900, CK => CLK, Q => n_1210, 
                           QN => n983);
   REGS_reg_45_30_inst : DFF_X1 port map( D => n12899, CK => CLK, Q => n_1211, 
                           QN => n984);
   REGS_reg_45_29_inst : DFF_X1 port map( D => n12898, CK => CLK, Q => n_1212, 
                           QN => n985);
   REGS_reg_45_28_inst : DFF_X1 port map( D => n12897, CK => CLK, Q => n_1213, 
                           QN => n4236);
   REGS_reg_45_27_inst : DFF_X1 port map( D => n12896, CK => CLK, Q => n_1214, 
                           QN => n4237);
   REGS_reg_45_26_inst : DFF_X1 port map( D => n12895, CK => CLK, Q => n_1215, 
                           QN => n4238);
   REGS_reg_45_25_inst : DFF_X1 port map( D => n12894, CK => CLK, Q => n_1216, 
                           QN => n4239);
   REGS_reg_45_24_inst : DFF_X1 port map( D => n12893, CK => CLK, Q => n_1217, 
                           QN => n4240);
   REGS_reg_44_31_inst : DFF_X1 port map( D => n12932, CK => CLK, Q => n52351, 
                           QN => n986);
   REGS_reg_44_30_inst : DFF_X1 port map( D => n12931, CK => CLK, Q => n52352, 
                           QN => n987);
   REGS_reg_44_29_inst : DFF_X1 port map( D => n12930, CK => CLK, Q => n52353, 
                           QN => n988);
   REGS_reg_44_28_inst : DFF_X1 port map( D => n12929, CK => CLK, Q => n52354, 
                           QN => n989);
   REGS_reg_44_27_inst : DFF_X1 port map( D => n12928, CK => CLK, Q => n52355, 
                           QN => n990);
   REGS_reg_44_26_inst : DFF_X1 port map( D => n12927, CK => CLK, Q => n52356, 
                           QN => n991);
   REGS_reg_44_25_inst : DFF_X1 port map( D => n12926, CK => CLK, Q => n52357, 
                           QN => n992);
   REGS_reg_44_24_inst : DFF_X1 port map( D => n12925, CK => CLK, Q => n52358, 
                           QN => n993);
   REGS_reg_43_31_inst : DFF_X1 port map( D => n12964, CK => CLK, Q => n16452, 
                           QN => n4241);
   REGS_reg_43_30_inst : DFF_X1 port map( D => n12963, CK => CLK, Q => n16451, 
                           QN => n4242);
   REGS_reg_43_29_inst : DFF_X1 port map( D => n12962, CK => CLK, Q => n16450, 
                           QN => n4243);
   REGS_reg_43_28_inst : DFF_X1 port map( D => n12961, CK => CLK, Q => n16449, 
                           QN => n4244);
   REGS_reg_43_27_inst : DFF_X1 port map( D => n12960, CK => CLK, Q => n16448, 
                           QN => n4245);
   REGS_reg_43_26_inst : DFF_X1 port map( D => n12959, CK => CLK, Q => n16447, 
                           QN => n4246);
   REGS_reg_43_25_inst : DFF_X1 port map( D => n12958, CK => CLK, Q => n16446, 
                           QN => n4247);
   REGS_reg_43_24_inst : DFF_X1 port map( D => n12957, CK => CLK, Q => n16445, 
                           QN => n4248);
   REGS_reg_42_31_inst : DFF_X1 port map( D => n12996, CK => CLK, Q => n16444, 
                           QN => n4249);
   REGS_reg_42_30_inst : DFF_X1 port map( D => n12995, CK => CLK, Q => n16443, 
                           QN => n4250);
   REGS_reg_42_29_inst : DFF_X1 port map( D => n12994, CK => CLK, Q => n16442, 
                           QN => n4251);
   REGS_reg_42_28_inst : DFF_X1 port map( D => n12993, CK => CLK, Q => n16441, 
                           QN => n4252);
   REGS_reg_42_27_inst : DFF_X1 port map( D => n12992, CK => CLK, Q => n16440, 
                           QN => n4253);
   REGS_reg_42_26_inst : DFF_X1 port map( D => n12991, CK => CLK, Q => n16439, 
                           QN => n4254);
   REGS_reg_42_25_inst : DFF_X1 port map( D => n12990, CK => CLK, Q => n16438, 
                           QN => n4255);
   REGS_reg_42_24_inst : DFF_X1 port map( D => n12989, CK => CLK, Q => n16437, 
                           QN => n4256);
   REGS_reg_41_31_inst : DFF_X1 port map( D => n13028, CK => CLK, Q => n_1218, 
                           QN => n994);
   REGS_reg_41_30_inst : DFF_X1 port map( D => n13027, CK => CLK, Q => n_1219, 
                           QN => n995);
   REGS_reg_41_29_inst : DFF_X1 port map( D => n13026, CK => CLK, Q => n_1220, 
                           QN => n1000);
   REGS_reg_41_28_inst : DFF_X1 port map( D => n13025, CK => CLK, Q => n_1221, 
                           QN => n1001);
   REGS_reg_41_27_inst : DFF_X1 port map( D => n13024, CK => CLK, Q => n_1222, 
                           QN => n1002);
   REGS_reg_41_26_inst : DFF_X1 port map( D => n13023, CK => CLK, Q => n_1223, 
                           QN => n1003);
   REGS_reg_41_25_inst : DFF_X1 port map( D => n13022, CK => CLK, Q => n_1224, 
                           QN => n1004);
   REGS_reg_41_24_inst : DFF_X1 port map( D => n13021, CK => CLK, Q => n_1225, 
                           QN => n1005);
   REGS_reg_40_31_inst : DFF_X1 port map( D => n13060, CK => CLK, Q => n_1226, 
                           QN => n1006);
   REGS_reg_40_30_inst : DFF_X1 port map( D => n13059, CK => CLK, Q => n_1227, 
                           QN => n1007);
   REGS_reg_40_29_inst : DFF_X1 port map( D => n13058, CK => CLK, Q => n_1228, 
                           QN => n1008);
   REGS_reg_40_28_inst : DFF_X1 port map( D => n13057, CK => CLK, Q => n_1229, 
                           QN => n1009);
   REGS_reg_40_27_inst : DFF_X1 port map( D => n13056, CK => CLK, Q => n_1230, 
                           QN => n1010);
   REGS_reg_40_26_inst : DFF_X1 port map( D => n13055, CK => CLK, Q => n_1231, 
                           QN => n1011);
   REGS_reg_40_25_inst : DFF_X1 port map( D => n13054, CK => CLK, Q => n_1232, 
                           QN => n1012);
   REGS_reg_40_24_inst : DFF_X1 port map( D => n13053, CK => CLK, Q => n_1233, 
                           QN => n1013);
   REGS_reg_37_31_inst : DFF_X1 port map( D => n13156, CK => CLK, Q => n52359, 
                           QN => n1014);
   REGS_reg_37_30_inst : DFF_X1 port map( D => n13155, CK => CLK, Q => n52360, 
                           QN => n1015);
   REGS_reg_37_29_inst : DFF_X1 port map( D => n13154, CK => CLK, Q => n52361, 
                           QN => n1016);
   REGS_reg_37_28_inst : DFF_X1 port map( D => n13153, CK => CLK, Q => n52362, 
                           QN => n1017);
   REGS_reg_37_27_inst : DFF_X1 port map( D => n13152, CK => CLK, Q => n52363, 
                           QN => n1018);
   REGS_reg_37_26_inst : DFF_X1 port map( D => n13151, CK => CLK, Q => n52364, 
                           QN => n1019);
   REGS_reg_37_25_inst : DFF_X1 port map( D => n13150, CK => CLK, Q => n52365, 
                           QN => n1020);
   REGS_reg_37_24_inst : DFF_X1 port map( D => n13149, CK => CLK, Q => n52366, 
                           QN => n1021);
   REGS_reg_36_31_inst : DFF_X1 port map( D => n13188, CK => CLK, Q => n52367, 
                           QN => n1022);
   REGS_reg_36_30_inst : DFF_X1 port map( D => n13187, CK => CLK, Q => n52368, 
                           QN => n1023);
   REGS_reg_36_29_inst : DFF_X1 port map( D => n13186, CK => CLK, Q => n52369, 
                           QN => n1024);
   REGS_reg_36_28_inst : DFF_X1 port map( D => n13185, CK => CLK, Q => n52370, 
                           QN => n1025);
   REGS_reg_36_27_inst : DFF_X1 port map( D => n13184, CK => CLK, Q => n52371, 
                           QN => n1026);
   REGS_reg_36_26_inst : DFF_X1 port map( D => n13183, CK => CLK, Q => n52372, 
                           QN => n1027);
   REGS_reg_36_25_inst : DFF_X1 port map( D => n13182, CK => CLK, Q => n52373, 
                           QN => n1028);
   REGS_reg_36_24_inst : DFF_X1 port map( D => n13181, CK => CLK, Q => n52374, 
                           QN => n1029);
   REGS_reg_35_31_inst : DFF_X1 port map( D => n13220, CK => CLK, Q => n16845, 
                           QN => n4273);
   REGS_reg_35_30_inst : DFF_X1 port map( D => n13219, CK => CLK, Q => n16843, 
                           QN => n4274);
   REGS_reg_35_29_inst : DFF_X1 port map( D => n13218, CK => CLK, Q => n16841, 
                           QN => n4275);
   REGS_reg_35_28_inst : DFF_X1 port map( D => n13217, CK => CLK, Q => n16839, 
                           QN => n4276);
   REGS_reg_35_27_inst : DFF_X1 port map( D => n13216, CK => CLK, Q => n16837, 
                           QN => n4277);
   REGS_reg_35_26_inst : DFF_X1 port map( D => n13215, CK => CLK, Q => n16835, 
                           QN => n4278);
   REGS_reg_35_25_inst : DFF_X1 port map( D => n13214, CK => CLK, Q => n16833, 
                           QN => n4279);
   REGS_reg_35_24_inst : DFF_X1 port map( D => n13213, CK => CLK, Q => n16831, 
                           QN => n4280);
   REGS_reg_34_31_inst : DFF_X1 port map( D => n13252, CK => CLK, Q => n16844, 
                           QN => n4281);
   REGS_reg_34_30_inst : DFF_X1 port map( D => n13251, CK => CLK, Q => n16842, 
                           QN => n4282);
   REGS_reg_34_29_inst : DFF_X1 port map( D => n13250, CK => CLK, Q => n16840, 
                           QN => n4283);
   REGS_reg_34_28_inst : DFF_X1 port map( D => n13249, CK => CLK, Q => n16838, 
                           QN => n4284);
   REGS_reg_34_27_inst : DFF_X1 port map( D => n13248, CK => CLK, Q => n16836, 
                           QN => n4285);
   REGS_reg_34_26_inst : DFF_X1 port map( D => n13247, CK => CLK, Q => n16834, 
                           QN => n4286);
   REGS_reg_34_25_inst : DFF_X1 port map( D => n13246, CK => CLK, Q => n16832, 
                           QN => n4287);
   REGS_reg_34_24_inst : DFF_X1 port map( D => n13245, CK => CLK, Q => n16830, 
                           QN => n4288);
   REGS_reg_33_31_inst : DFF_X1 port map( D => n13284, CK => CLK, Q => n52375, 
                           QN => n1030);
   REGS_reg_33_30_inst : DFF_X1 port map( D => n13283, CK => CLK, Q => n52376, 
                           QN => n1031);
   REGS_reg_33_29_inst : DFF_X1 port map( D => n13282, CK => CLK, Q => n52377, 
                           QN => n1032);
   REGS_reg_33_28_inst : DFF_X1 port map( D => n13281, CK => CLK, Q => n52378, 
                           QN => n1033);
   REGS_reg_33_27_inst : DFF_X1 port map( D => n13280, CK => CLK, Q => n52379, 
                           QN => n1034);
   REGS_reg_33_26_inst : DFF_X1 port map( D => n13279, CK => CLK, Q => n52380, 
                           QN => n1035);
   REGS_reg_33_25_inst : DFF_X1 port map( D => n13278, CK => CLK, Q => n52381, 
                           QN => n1036);
   REGS_reg_33_24_inst : DFF_X1 port map( D => n13277, CK => CLK, Q => n52382, 
                           QN => n1037);
   REGS_reg_32_31_inst : DFF_X1 port map( D => n13316, CK => CLK, Q => n52383, 
                           QN => n1038);
   REGS_reg_32_30_inst : DFF_X1 port map( D => n13315, CK => CLK, Q => n52384, 
                           QN => n1039);
   REGS_reg_32_29_inst : DFF_X1 port map( D => n13314, CK => CLK, Q => n52385, 
                           QN => n1040);
   REGS_reg_32_28_inst : DFF_X1 port map( D => n13313, CK => CLK, Q => n52386, 
                           QN => n1041);
   REGS_reg_32_27_inst : DFF_X1 port map( D => n13312, CK => CLK, Q => n52387, 
                           QN => n1042);
   REGS_reg_32_26_inst : DFF_X1 port map( D => n13311, CK => CLK, Q => n52388, 
                           QN => n1043);
   REGS_reg_32_25_inst : DFF_X1 port map( D => n13310, CK => CLK, Q => n52389, 
                           QN => n1044);
   REGS_reg_32_24_inst : DFF_X1 port map( D => n13309, CK => CLK, Q => n52390, 
                           QN => n1045);
   REGS_reg_31_31_inst : DFF_X1 port map( D => n13348, CK => CLK, Q => n776, QN
                           => n3948);
   REGS_reg_31_30_inst : DFF_X1 port map( D => n13347, CK => CLK, Q => n777, QN
                           => n3949);
   REGS_reg_31_29_inst : DFF_X1 port map( D => n13346, CK => CLK, Q => n778, QN
                           => n3950);
   REGS_reg_31_28_inst : DFF_X1 port map( D => n13345, CK => CLK, Q => n779, QN
                           => n3951);
   REGS_reg_31_27_inst : DFF_X1 port map( D => n13344, CK => CLK, Q => n780, QN
                           => n3952);
   REGS_reg_31_26_inst : DFF_X1 port map( D => n13343, CK => CLK, Q => n781, QN
                           => n3953);
   REGS_reg_31_25_inst : DFF_X1 port map( D => n13342, CK => CLK, Q => n782, QN
                           => n3954);
   REGS_reg_31_24_inst : DFF_X1 port map( D => n13341, CK => CLK, Q => n783, QN
                           => n3955);
   REGS_reg_30_31_inst : DFF_X1 port map( D => n13380, CK => CLK, Q => n16158, 
                           QN => n36);
   REGS_reg_30_30_inst : DFF_X1 port map( D => n13379, CK => CLK, Q => n16156, 
                           QN => n37);
   REGS_reg_30_29_inst : DFF_X1 port map( D => n13378, CK => CLK, Q => n16154, 
                           QN => n38);
   REGS_reg_30_28_inst : DFF_X1 port map( D => n13377, CK => CLK, Q => n16152, 
                           QN => n39);
   REGS_reg_30_27_inst : DFF_X1 port map( D => n13376, CK => CLK, Q => n16150, 
                           QN => n40);
   REGS_reg_30_26_inst : DFF_X1 port map( D => n13375, CK => CLK, Q => n16148, 
                           QN => n41);
   REGS_reg_30_25_inst : DFF_X1 port map( D => n13374, CK => CLK, Q => n16146, 
                           QN => n42);
   REGS_reg_30_24_inst : DFF_X1 port map( D => n13373, CK => CLK, Q => n16144, 
                           QN => n43);
   REGS_reg_29_31_inst : DFF_X1 port map( D => n13412, CK => CLK, Q => n16157, 
                           QN => n44);
   REGS_reg_29_30_inst : DFF_X1 port map( D => n13411, CK => CLK, Q => n16155, 
                           QN => n45);
   REGS_reg_29_29_inst : DFF_X1 port map( D => n13410, CK => CLK, Q => n16153, 
                           QN => n46);
   REGS_reg_29_28_inst : DFF_X1 port map( D => n13409, CK => CLK, Q => n16151, 
                           QN => n47);
   REGS_reg_29_27_inst : DFF_X1 port map( D => n13408, CK => CLK, Q => n16149, 
                           QN => n48);
   REGS_reg_29_26_inst : DFF_X1 port map( D => n13407, CK => CLK, Q => n16147, 
                           QN => n49);
   REGS_reg_29_25_inst : DFF_X1 port map( D => n13406, CK => CLK, Q => n16145, 
                           QN => n50);
   REGS_reg_29_24_inst : DFF_X1 port map( D => n13405, CK => CLK, Q => n16143, 
                           QN => n51);
   REGS_reg_26_31_inst : DFF_X1 port map( D => n13508, CK => CLK, Q => n_1234, 
                           QN => n52);
   REGS_reg_26_30_inst : DFF_X1 port map( D => n13507, CK => CLK, Q => n_1235, 
                           QN => n53);
   REGS_reg_26_29_inst : DFF_X1 port map( D => n13506, CK => CLK, Q => n_1236, 
                           QN => n54);
   REGS_reg_26_28_inst : DFF_X1 port map( D => n13505, CK => CLK, Q => n_1237, 
                           QN => n55);
   REGS_reg_26_27_inst : DFF_X1 port map( D => n13504, CK => CLK, Q => n_1238, 
                           QN => n56);
   REGS_reg_26_26_inst : DFF_X1 port map( D => n13503, CK => CLK, Q => n_1239, 
                           QN => n57);
   REGS_reg_26_25_inst : DFF_X1 port map( D => n13502, CK => CLK, Q => n_1240, 
                           QN => n58);
   REGS_reg_26_24_inst : DFF_X1 port map( D => n13501, CK => CLK, Q => n_1241, 
                           QN => n59);
   REGS_reg_25_31_inst : DFF_X1 port map( D => n13540, CK => CLK, Q => n_1242, 
                           QN => n60);
   REGS_reg_25_30_inst : DFF_X1 port map( D => n13539, CK => CLK, Q => n_1243, 
                           QN => n61);
   REGS_reg_25_29_inst : DFF_X1 port map( D => n13538, CK => CLK, Q => n_1244, 
                           QN => n62);
   REGS_reg_25_28_inst : DFF_X1 port map( D => n13537, CK => CLK, Q => n_1245, 
                           QN => n63);
   REGS_reg_25_27_inst : DFF_X1 port map( D => n13536, CK => CLK, Q => n_1246, 
                           QN => n64);
   REGS_reg_25_26_inst : DFF_X1 port map( D => n13535, CK => CLK, Q => n_1247, 
                           QN => n65);
   REGS_reg_25_25_inst : DFF_X1 port map( D => n13534, CK => CLK, Q => n_1248, 
                           QN => n66);
   REGS_reg_25_24_inst : DFF_X1 port map( D => n13533, CK => CLK, Q => n_1249, 
                           QN => n67);
   REGS_reg_24_31_inst : DFF_X1 port map( D => n13572, CK => CLK, Q => n15970, 
                           QN => n68);
   REGS_reg_24_30_inst : DFF_X1 port map( D => n13571, CK => CLK, Q => n15966, 
                           QN => n69);
   REGS_reg_24_29_inst : DFF_X1 port map( D => n13570, CK => CLK, Q => n15962, 
                           QN => n70);
   REGS_reg_24_28_inst : DFF_X1 port map( D => n13569, CK => CLK, Q => n15958, 
                           QN => n71);
   REGS_reg_24_27_inst : DFF_X1 port map( D => n13568, CK => CLK, Q => n15954, 
                           QN => n72);
   REGS_reg_24_26_inst : DFF_X1 port map( D => n13567, CK => CLK, Q => n15950, 
                           QN => n73);
   REGS_reg_24_25_inst : DFF_X1 port map( D => n13566, CK => CLK, Q => n15922, 
                           QN => n74);
   REGS_reg_24_24_inst : DFF_X1 port map( D => n13565, CK => CLK, Q => n15918, 
                           QN => n75);
   REGS_reg_23_31_inst : DFF_X1 port map( D => n13604, CK => CLK, Q => n15971, 
                           QN => n76);
   REGS_reg_23_30_inst : DFF_X1 port map( D => n13603, CK => CLK, Q => n15967, 
                           QN => n77);
   REGS_reg_23_29_inst : DFF_X1 port map( D => n13602, CK => CLK, Q => n15963, 
                           QN => n78);
   REGS_reg_23_28_inst : DFF_X1 port map( D => n13601, CK => CLK, Q => n15959, 
                           QN => n79);
   REGS_reg_23_27_inst : DFF_X1 port map( D => n13600, CK => CLK, Q => n15955, 
                           QN => n100);
   REGS_reg_23_26_inst : DFF_X1 port map( D => n13599, CK => CLK, Q => n15951, 
                           QN => n101);
   REGS_reg_23_25_inst : DFF_X1 port map( D => n13598, CK => CLK, Q => n15947, 
                           QN => n102);
   REGS_reg_23_24_inst : DFF_X1 port map( D => n13597, CK => CLK, Q => n15919, 
                           QN => n103);
   REGS_reg_18_31_inst : DFF_X1 port map( D => n13764, CK => CLK, Q => n832, QN
                           => n3996);
   REGS_reg_18_30_inst : DFF_X1 port map( D => n13763, CK => CLK, Q => n833, QN
                           => n3997);
   REGS_reg_18_29_inst : DFF_X1 port map( D => n13762, CK => CLK, Q => n834, QN
                           => n3998);
   REGS_reg_18_28_inst : DFF_X1 port map( D => n13761, CK => CLK, Q => n835, QN
                           => n3999);
   REGS_reg_18_27_inst : DFF_X1 port map( D => n13760, CK => CLK, Q => n836, QN
                           => n4000);
   REGS_reg_18_26_inst : DFF_X1 port map( D => n13759, CK => CLK, Q => n837, QN
                           => n4001);
   REGS_reg_18_25_inst : DFF_X1 port map( D => n13758, CK => CLK, Q => n838, QN
                           => n4002);
   REGS_reg_18_24_inst : DFF_X1 port map( D => n13757, CK => CLK, Q => n839, QN
                           => n4003);
   REGS_reg_17_31_inst : DFF_X1 port map( D => n13796, CK => CLK, Q => n840, QN
                           => n4004);
   REGS_reg_17_30_inst : DFF_X1 port map( D => n13795, CK => CLK, Q => n841, QN
                           => n4005);
   REGS_reg_17_29_inst : DFF_X1 port map( D => n13794, CK => CLK, Q => n842, QN
                           => n4006);
   REGS_reg_17_28_inst : DFF_X1 port map( D => n13793, CK => CLK, Q => n843, QN
                           => n4007);
   REGS_reg_17_27_inst : DFF_X1 port map( D => n13792, CK => CLK, Q => n844, QN
                           => n4008);
   REGS_reg_17_26_inst : DFF_X1 port map( D => n13791, CK => CLK, Q => n845, QN
                           => n4009);
   REGS_reg_17_25_inst : DFF_X1 port map( D => n13790, CK => CLK, Q => n846, QN
                           => n4010);
   REGS_reg_17_24_inst : DFF_X1 port map( D => n13789, CK => CLK, Q => n847, QN
                           => n4011);
   REGS_reg_16_31_inst : DFF_X1 port map( D => n13828, CK => CLK, Q => n51600, 
                           QN => n128);
   REGS_reg_16_30_inst : DFF_X1 port map( D => n13827, CK => CLK, Q => n51601, 
                           QN => n129);
   REGS_reg_16_29_inst : DFF_X1 port map( D => n13826, CK => CLK, Q => n51602, 
                           QN => n130);
   REGS_reg_16_28_inst : DFF_X1 port map( D => n13825, CK => CLK, Q => n51603, 
                           QN => n131);
   REGS_reg_16_27_inst : DFF_X1 port map( D => n13824, CK => CLK, Q => n51604, 
                           QN => n132);
   REGS_reg_16_26_inst : DFF_X1 port map( D => n13823, CK => CLK, Q => n51605, 
                           QN => n133);
   REGS_reg_16_25_inst : DFF_X1 port map( D => n13822, CK => CLK, Q => n51606, 
                           QN => n134);
   REGS_reg_16_24_inst : DFF_X1 port map( D => n13821, CK => CLK, Q => n51607, 
                           QN => n135);
   REGS_reg_135_18_inst : DFF_X1 port map( D => n10007, CK => CLK, Q => n54534,
                           QN => n389);
   REGS_reg_135_17_inst : DFF_X1 port map( D => n10006, CK => CLK, Q => n54533,
                           QN => n390);
   REGS_reg_135_16_inst : DFF_X1 port map( D => n10005, CK => CLK, Q => n54532,
                           QN => n391);
   REGS_reg_135_15_inst : DFF_X1 port map( D => n10004, CK => CLK, Q => n54531,
                           QN => n392);
   REGS_reg_135_14_inst : DFF_X1 port map( D => n10003, CK => CLK, Q => n54530,
                           QN => n393);
   REGS_reg_135_13_inst : DFF_X1 port map( D => n10002, CK => CLK, Q => n54529,
                           QN => n394);
   REGS_reg_135_12_inst : DFF_X1 port map( D => n10001, CK => CLK, Q => n54528,
                           QN => n395);
   REGS_reg_135_11_inst : DFF_X1 port map( D => n10000, CK => CLK, Q => n54535,
                           QN => n396);
   REGS_reg_15_31_inst : DFF_X1 port map( D => n13860, CK => CLK, Q => n848, QN
                           => n4100);
   REGS_reg_15_30_inst : DFF_X1 port map( D => n13859, CK => CLK, Q => n849, QN
                           => n4101);
   REGS_reg_15_29_inst : DFF_X1 port map( D => n13858, CK => CLK, Q => n850, QN
                           => n4102);
   REGS_reg_15_28_inst : DFF_X1 port map( D => n13857, CK => CLK, Q => n851, QN
                           => n4103);
   REGS_reg_15_27_inst : DFF_X1 port map( D => n13856, CK => CLK, Q => n852, QN
                           => n4104);
   REGS_reg_15_26_inst : DFF_X1 port map( D => n13855, CK => CLK, Q => n853, QN
                           => n4105);
   REGS_reg_15_25_inst : DFF_X1 port map( D => n13854, CK => CLK, Q => n854, QN
                           => n4106);
   REGS_reg_15_24_inst : DFF_X1 port map( D => n13853, CK => CLK, Q => n855, QN
                           => n4107);
   REGS_reg_14_31_inst : DFF_X1 port map( D => n13892, CK => CLK, Q => n856, QN
                           => n4108);
   REGS_reg_14_30_inst : DFF_X1 port map( D => n13891, CK => CLK, Q => n857, QN
                           => n4109);
   REGS_reg_14_29_inst : DFF_X1 port map( D => n13890, CK => CLK, Q => n858, QN
                           => n4110);
   REGS_reg_14_28_inst : DFF_X1 port map( D => n13889, CK => CLK, Q => n859, QN
                           => n4111);
   REGS_reg_14_27_inst : DFF_X1 port map( D => n13888, CK => CLK, Q => n860, QN
                           => n4112);
   REGS_reg_14_26_inst : DFF_X1 port map( D => n13887, CK => CLK, Q => n861, QN
                           => n4113);
   REGS_reg_14_25_inst : DFF_X1 port map( D => n13886, CK => CLK, Q => n862, QN
                           => n4114);
   REGS_reg_14_24_inst : DFF_X1 port map( D => n13885, CK => CLK, Q => n863, QN
                           => n4115);
   REGS_reg_13_31_inst : DFF_X1 port map( D => n13924, CK => CLK, Q => n16436, 
                           QN => n4116);
   REGS_reg_13_30_inst : DFF_X1 port map( D => n13923, CK => CLK, Q => n16435, 
                           QN => n4117);
   REGS_reg_13_29_inst : DFF_X1 port map( D => n13922, CK => CLK, Q => n16434, 
                           QN => n4118);
   REGS_reg_13_28_inst : DFF_X1 port map( D => n13921, CK => CLK, Q => n16433, 
                           QN => n4119);
   REGS_reg_13_27_inst : DFF_X1 port map( D => n13920, CK => CLK, Q => n16432, 
                           QN => n4120);
   REGS_reg_13_26_inst : DFF_X1 port map( D => n13919, CK => CLK, Q => n16431, 
                           QN => n4121);
   REGS_reg_13_25_inst : DFF_X1 port map( D => n13918, CK => CLK, Q => n16430, 
                           QN => n4122);
   REGS_reg_13_24_inst : DFF_X1 port map( D => n13917, CK => CLK, Q => n16429, 
                           QN => n4123);
   REGS_reg_12_31_inst : DFF_X1 port map( D => n13956, CK => CLK, Q => n16428, 
                           QN => n4124);
   REGS_reg_12_30_inst : DFF_X1 port map( D => n13955, CK => CLK, Q => n16427, 
                           QN => n4125);
   REGS_reg_12_29_inst : DFF_X1 port map( D => n13954, CK => CLK, Q => n16426, 
                           QN => n4126);
   REGS_reg_12_28_inst : DFF_X1 port map( D => n13953, CK => CLK, Q => n16425, 
                           QN => n4127);
   REGS_reg_12_27_inst : DFF_X1 port map( D => n13952, CK => CLK, Q => n16424, 
                           QN => n4128);
   REGS_reg_12_26_inst : DFF_X1 port map( D => n13951, CK => CLK, Q => n16423, 
                           QN => n4129);
   REGS_reg_12_25_inst : DFF_X1 port map( D => n13950, CK => CLK, Q => n16422, 
                           QN => n4130);
   REGS_reg_12_24_inst : DFF_X1 port map( D => n13949, CK => CLK, Q => n16421, 
                           QN => n4131);
   REGS_reg_11_31_inst : DFF_X1 port map( D => n13988, CK => CLK, Q => n51608, 
                           QN => n405);
   REGS_reg_11_30_inst : DFF_X1 port map( D => n13987, CK => CLK, Q => n51609, 
                           QN => n406);
   REGS_reg_11_29_inst : DFF_X1 port map( D => n13986, CK => CLK, Q => n51610, 
                           QN => n407);
   REGS_reg_11_28_inst : DFF_X1 port map( D => n13985, CK => CLK, Q => n51611, 
                           QN => n408);
   REGS_reg_11_27_inst : DFF_X1 port map( D => n13984, CK => CLK, Q => n51612, 
                           QN => n409);
   REGS_reg_11_26_inst : DFF_X1 port map( D => n13983, CK => CLK, Q => n51613, 
                           QN => n410);
   REGS_reg_11_25_inst : DFF_X1 port map( D => n13982, CK => CLK, Q => n51614, 
                           QN => n411);
   REGS_reg_11_24_inst : DFF_X1 port map( D => n13981, CK => CLK, Q => n51615, 
                           QN => n412);
   REGS_reg_10_31_inst : DFF_X1 port map( D => n14020, CK => CLK, Q => n51616, 
                           QN => n453);
   REGS_reg_10_30_inst : DFF_X1 port map( D => n14019, CK => CLK, Q => n51617, 
                           QN => n454);
   REGS_reg_10_29_inst : DFF_X1 port map( D => n14018, CK => CLK, Q => n51618, 
                           QN => n455);
   REGS_reg_10_28_inst : DFF_X1 port map( D => n14017, CK => CLK, Q => n51619, 
                           QN => n456);
   REGS_reg_10_27_inst : DFF_X1 port map( D => n14016, CK => CLK, Q => n51620, 
                           QN => n457);
   REGS_reg_10_26_inst : DFF_X1 port map( D => n14015, CK => CLK, Q => n51621, 
                           QN => n458);
   REGS_reg_10_25_inst : DFF_X1 port map( D => n14014, CK => CLK, Q => n51622, 
                           QN => n459);
   REGS_reg_10_24_inst : DFF_X1 port map( D => n14013, CK => CLK, Q => n51623, 
                           QN => n460);
   REGS_reg_9_31_inst : DFF_X1 port map( D => n14052, CK => CLK, Q => n16420, 
                           QN => n4132);
   REGS_reg_9_30_inst : DFF_X1 port map( D => n14051, CK => CLK, Q => n16419, 
                           QN => n4133);
   REGS_reg_9_29_inst : DFF_X1 port map( D => n14050, CK => CLK, Q => n16418, 
                           QN => n4134);
   REGS_reg_9_28_inst : DFF_X1 port map( D => n14049, CK => CLK, Q => n16417, 
                           QN => n4135);
   REGS_reg_9_27_inst : DFF_X1 port map( D => n14048, CK => CLK, Q => n16416, 
                           QN => n4136);
   REGS_reg_9_26_inst : DFF_X1 port map( D => n14047, CK => CLK, Q => n16415, 
                           QN => n4137);
   REGS_reg_9_25_inst : DFF_X1 port map( D => n14046, CK => CLK, Q => n16414, 
                           QN => n4138);
   REGS_reg_9_24_inst : DFF_X1 port map( D => n14045, CK => CLK, Q => n16413, 
                           QN => n4139);
   REGS_reg_8_31_inst : DFF_X1 port map( D => n14084, CK => CLK, Q => n_1250, 
                           QN => n4140);
   REGS_reg_8_30_inst : DFF_X1 port map( D => n14083, CK => CLK, Q => n_1251, 
                           QN => n4141);
   REGS_reg_8_29_inst : DFF_X1 port map( D => n14082, CK => CLK, Q => n_1252, 
                           QN => n4142);
   REGS_reg_8_28_inst : DFF_X1 port map( D => n14081, CK => CLK, Q => n_1253, 
                           QN => n4143);
   REGS_reg_8_27_inst : DFF_X1 port map( D => n14080, CK => CLK, Q => n_1254, 
                           QN => n4144);
   REGS_reg_8_26_inst : DFF_X1 port map( D => n14079, CK => CLK, Q => n_1255, 
                           QN => n4145);
   REGS_reg_8_25_inst : DFF_X1 port map( D => n14078, CK => CLK, Q => n_1256, 
                           QN => n4146);
   REGS_reg_8_24_inst : DFF_X1 port map( D => n14077, CK => CLK, Q => n_1257, 
                           QN => n4147);
   REGS_reg_6_31_inst : DFF_X1 port map( D => n14148, CK => CLK, Q => n51624, 
                           QN => n461);
   REGS_reg_6_30_inst : DFF_X1 port map( D => n14147, CK => CLK, Q => n51625, 
                           QN => n462);
   REGS_reg_6_29_inst : DFF_X1 port map( D => n14146, CK => CLK, Q => n51626, 
                           QN => n463);
   REGS_reg_6_28_inst : DFF_X1 port map( D => n14145, CK => CLK, Q => n51627, 
                           QN => n464);
   REGS_reg_6_27_inst : DFF_X1 port map( D => n14144, CK => CLK, Q => n51628, 
                           QN => n465);
   REGS_reg_6_26_inst : DFF_X1 port map( D => n14143, CK => CLK, Q => n51629, 
                           QN => n466);
   REGS_reg_6_25_inst : DFF_X1 port map( D => n14142, CK => CLK, Q => n51630, 
                           QN => n467);
   REGS_reg_6_24_inst : DFF_X1 port map( D => n14141, CK => CLK, Q => n51631, 
                           QN => n468);
   REGS_reg_5_31_inst : DFF_X1 port map( D => n14180, CK => CLK, Q => n_1258, 
                           QN => n4148);
   REGS_reg_5_30_inst : DFF_X1 port map( D => n14179, CK => CLK, Q => n_1259, 
                           QN => n4149);
   REGS_reg_5_29_inst : DFF_X1 port map( D => n14178, CK => CLK, Q => n_1260, 
                           QN => n4150);
   REGS_reg_5_28_inst : DFF_X1 port map( D => n14177, CK => CLK, Q => n_1261, 
                           QN => n4151);
   REGS_reg_5_27_inst : DFF_X1 port map( D => n14176, CK => CLK, Q => n_1262, 
                           QN => n4152);
   REGS_reg_5_26_inst : DFF_X1 port map( D => n14175, CK => CLK, Q => n_1263, 
                           QN => n4153);
   REGS_reg_5_25_inst : DFF_X1 port map( D => n14174, CK => CLK, Q => n_1264, 
                           QN => n4154);
   REGS_reg_5_24_inst : DFF_X1 port map( D => n14173, CK => CLK, Q => n_1265, 
                           QN => n4155);
   REGS_reg_4_31_inst : DFF_X1 port map( D => n14212, CK => CLK, Q => n_1266, 
                           QN => n4156);
   REGS_reg_4_30_inst : DFF_X1 port map( D => n14211, CK => CLK, Q => n_1267, 
                           QN => n4157);
   REGS_reg_4_29_inst : DFF_X1 port map( D => n14210, CK => CLK, Q => n_1268, 
                           QN => n4158);
   REGS_reg_4_28_inst : DFF_X1 port map( D => n14209, CK => CLK, Q => n_1269, 
                           QN => n4159);
   REGS_reg_4_27_inst : DFF_X1 port map( D => n14208, CK => CLK, Q => n_1270, 
                           QN => n4160);
   REGS_reg_4_26_inst : DFF_X1 port map( D => n14207, CK => CLK, Q => n_1271, 
                           QN => n4161);
   REGS_reg_4_25_inst : DFF_X1 port map( D => n14206, CK => CLK, Q => n_1272, 
                           QN => n4162);
   REGS_reg_4_24_inst : DFF_X1 port map( D => n14205, CK => CLK, Q => n_1273, 
                           QN => n4163);
   REGS_reg_1_31_inst : DFF_X1 port map( D => n14308, CK => CLK, Q => n15426, 
                           QN => n469);
   REGS_reg_1_30_inst : DFF_X1 port map( D => n14307, CK => CLK, Q => n15425, 
                           QN => n470);
   REGS_reg_1_29_inst : DFF_X1 port map( D => n14306, CK => CLK, Q => n15424, 
                           QN => n471);
   REGS_reg_1_28_inst : DFF_X1 port map( D => n14305, CK => CLK, Q => n15423, 
                           QN => n472);
   REGS_reg_1_27_inst : DFF_X1 port map( D => n14304, CK => CLK, Q => n15422, 
                           QN => n473);
   REGS_reg_1_26_inst : DFF_X1 port map( D => n14303, CK => CLK, Q => n15421, 
                           QN => n476);
   REGS_reg_1_25_inst : DFF_X1 port map( D => n14302, CK => CLK, Q => n15420, 
                           QN => n477);
   REGS_reg_1_24_inst : DFF_X1 port map( D => n14301, CK => CLK, Q => n15419, 
                           QN => n478);
   REGS_reg_0_31_inst : DFF_X1 port map( D => n14340, CK => CLK, Q => n15418, 
                           QN => n479);
   REGS_reg_0_30_inst : DFF_X1 port map( D => n14339, CK => CLK, Q => n15417, 
                           QN => n480);
   REGS_reg_0_29_inst : DFF_X1 port map( D => n14338, CK => CLK, Q => n15416, 
                           QN => n481);
   REGS_reg_0_28_inst : DFF_X1 port map( D => n14337, CK => CLK, Q => n15415, 
                           QN => n482);
   REGS_reg_0_27_inst : DFF_X1 port map( D => n14336, CK => CLK, Q => n15414, 
                           QN => n483);
   REGS_reg_0_26_inst : DFF_X1 port map( D => n14335, CK => CLK, Q => n15413, 
                           QN => n484);
   REGS_reg_0_25_inst : DFF_X1 port map( D => n14334, CK => CLK, Q => n15412, 
                           QN => n485);
   REGS_reg_0_24_inst : DFF_X1 port map( D => n14333, CK => CLK, Q => n15411, 
                           QN => n486);
   REGS_reg_7_31_inst : DFF_X1 port map( D => n14116, CK => CLK, Q => n51648, 
                           QN => n397);
   REGS_reg_7_30_inst : DFF_X1 port map( D => n14115, CK => CLK, Q => n51649, 
                           QN => n398);
   REGS_reg_7_29_inst : DFF_X1 port map( D => n14114, CK => CLK, Q => n51650, 
                           QN => n399);
   REGS_reg_7_28_inst : DFF_X1 port map( D => n14113, CK => CLK, Q => n51651, 
                           QN => n400);
   REGS_reg_7_27_inst : DFF_X1 port map( D => n14112, CK => CLK, Q => n51652, 
                           QN => n401);
   REGS_reg_7_26_inst : DFF_X1 port map( D => n14111, CK => CLK, Q => n51653, 
                           QN => n402);
   REGS_reg_7_25_inst : DFF_X1 port map( D => n14110, CK => CLK, Q => n51654, 
                           QN => n403);
   REGS_reg_7_24_inst : DFF_X1 port map( D => n14109, CK => CLK, Q => n51655, 
                           QN => n404);
   REGS_reg_127_31_inst : DFF_X1 port map( D => n10276, CK => CLK, Q => n15672,
                           QN => n1046);
   REGS_reg_127_30_inst : DFF_X1 port map( D => n10275, CK => CLK, Q => n15669,
                           QN => n1047);
   REGS_reg_127_29_inst : DFF_X1 port map( D => n10274, CK => CLK, Q => n15666,
                           QN => n1048);
   REGS_reg_127_28_inst : DFF_X1 port map( D => n10273, CK => CLK, Q => n15663,
                           QN => n1049);
   REGS_reg_127_27_inst : DFF_X1 port map( D => n10272, CK => CLK, Q => n15684,
                           QN => n1050);
   REGS_reg_127_26_inst : DFF_X1 port map( D => n10271, CK => CLK, Q => n15681,
                           QN => n1051);
   REGS_reg_127_25_inst : DFF_X1 port map( D => n10270, CK => CLK, Q => n15678,
                           QN => n1052);
   REGS_reg_127_24_inst : DFF_X1 port map( D => n10269, CK => CLK, Q => n15675,
                           QN => n1053);
   REGS_reg_124_31_inst : DFF_X1 port map( D => n10372, CK => CLK, Q => n51664,
                           QN => n1054);
   REGS_reg_124_30_inst : DFF_X1 port map( D => n10371, CK => CLK, Q => n51665,
                           QN => n1055);
   REGS_reg_124_29_inst : DFF_X1 port map( D => n10370, CK => CLK, Q => n51666,
                           QN => n1056);
   REGS_reg_124_28_inst : DFF_X1 port map( D => n10369, CK => CLK, Q => n51667,
                           QN => n1057);
   REGS_reg_124_27_inst : DFF_X1 port map( D => n10368, CK => CLK, Q => n51668,
                           QN => n1058);
   REGS_reg_124_26_inst : DFF_X1 port map( D => n10367, CK => CLK, Q => n51669,
                           QN => n1059);
   REGS_reg_124_25_inst : DFF_X1 port map( D => n10366, CK => CLK, Q => n51670,
                           QN => n1060);
   REGS_reg_124_24_inst : DFF_X1 port map( D => n10365, CK => CLK, Q => n51671,
                           QN => n1061);
   REGS_reg_123_31_inst : DFF_X1 port map( D => n10404, CK => CLK, Q => n51672,
                           QN => n1062);
   REGS_reg_123_30_inst : DFF_X1 port map( D => n10403, CK => CLK, Q => n51673,
                           QN => n1063);
   REGS_reg_123_29_inst : DFF_X1 port map( D => n10402, CK => CLK, Q => n51674,
                           QN => n1064);
   REGS_reg_123_28_inst : DFF_X1 port map( D => n10401, CK => CLK, Q => n51675,
                           QN => n1065);
   REGS_reg_123_27_inst : DFF_X1 port map( D => n10400, CK => CLK, Q => n51676,
                           QN => n1066);
   REGS_reg_123_26_inst : DFF_X1 port map( D => n10399, CK => CLK, Q => n51677,
                           QN => n1067);
   REGS_reg_123_25_inst : DFF_X1 port map( D => n10398, CK => CLK, Q => n51678,
                           QN => n1068);
   REGS_reg_123_24_inst : DFF_X1 port map( D => n10397, CK => CLK, Q => n51679,
                           QN => n1069);
   REGS_reg_121_27_inst : DFF_X1 port map( D => n10464, CK => CLK, Q => n52508,
                           QN => n1070);
   REGS_reg_121_26_inst : DFF_X1 port map( D => n10463, CK => CLK, Q => n52509,
                           QN => n1071);
   REGS_reg_121_25_inst : DFF_X1 port map( D => n10462, CK => CLK, Q => n52510,
                           QN => n1072);
   REGS_reg_121_24_inst : DFF_X1 port map( D => n10461, CK => CLK, Q => n52511,
                           QN => n1073);
   REGS_reg_120_31_inst : DFF_X1 port map( D => n10500, CK => CLK, Q => n15498,
                           QN => n1074);
   REGS_reg_120_30_inst : DFF_X1 port map( D => n10499, CK => CLK, Q => n15497,
                           QN => n1075);
   REGS_reg_120_29_inst : DFF_X1 port map( D => n10498, CK => CLK, Q => n15496,
                           QN => n1076);
   REGS_reg_120_28_inst : DFF_X1 port map( D => n10497, CK => CLK, Q => n15495,
                           QN => n1077);
   REGS_reg_120_27_inst : DFF_X1 port map( D => n10496, CK => CLK, Q => n15494,
                           QN => n1078);
   REGS_reg_120_26_inst : DFF_X1 port map( D => n10495, CK => CLK, Q => n15493,
                           QN => n1079);
   REGS_reg_120_25_inst : DFF_X1 port map( D => n10494, CK => CLK, Q => n15492,
                           QN => n1080);
   REGS_reg_120_24_inst : DFF_X1 port map( D => n10493, CK => CLK, Q => n15491,
                           QN => n1081);
   REGS_reg_119_31_inst : DFF_X1 port map( D => n10532, CK => CLK, Q => n15490,
                           QN => n1082);
   REGS_reg_119_30_inst : DFF_X1 port map( D => n10531, CK => CLK, Q => n15489,
                           QN => n1083);
   REGS_reg_119_29_inst : DFF_X1 port map( D => n10530, CK => CLK, Q => n15488,
                           QN => n1084);
   REGS_reg_119_28_inst : DFF_X1 port map( D => n10529, CK => CLK, Q => n15487,
                           QN => n1085);
   REGS_reg_119_27_inst : DFF_X1 port map( D => n10528, CK => CLK, Q => n15486,
                           QN => n1086);
   REGS_reg_119_26_inst : DFF_X1 port map( D => n10527, CK => CLK, Q => n15485,
                           QN => n1087);
   REGS_reg_119_25_inst : DFF_X1 port map( D => n10526, CK => CLK, Q => n15484,
                           QN => n1088);
   REGS_reg_119_24_inst : DFF_X1 port map( D => n10525, CK => CLK, Q => n15483,
                           QN => n1089);
   REGS_reg_118_31_inst : DFF_X1 port map( D => n10564, CK => CLK, Q => n52512,
                           QN => n1090);
   REGS_reg_118_30_inst : DFF_X1 port map( D => n10563, CK => CLK, Q => n52513,
                           QN => n1091);
   REGS_reg_118_29_inst : DFF_X1 port map( D => n10562, CK => CLK, Q => n52514,
                           QN => n1092);
   REGS_reg_118_28_inst : DFF_X1 port map( D => n10561, CK => CLK, Q => n52515,
                           QN => n1093);
   REGS_reg_118_27_inst : DFF_X1 port map( D => n10560, CK => CLK, Q => n52516,
                           QN => n1094);
   REGS_reg_118_26_inst : DFF_X1 port map( D => n10559, CK => CLK, Q => n52517,
                           QN => n1095);
   REGS_reg_118_25_inst : DFF_X1 port map( D => n10558, CK => CLK, Q => n52518,
                           QN => n1096);
   REGS_reg_118_24_inst : DFF_X1 port map( D => n10557, CK => CLK, Q => n52519,
                           QN => n1097);
   REGS_reg_117_31_inst : DFF_X1 port map( D => n10596, CK => CLK, Q => n52520,
                           QN => n1098);
   REGS_reg_117_30_inst : DFF_X1 port map( D => n10595, CK => CLK, Q => n52521,
                           QN => n1099);
   REGS_reg_117_29_inst : DFF_X1 port map( D => n10594, CK => CLK, Q => n52522,
                           QN => n1100);
   REGS_reg_117_28_inst : DFF_X1 port map( D => n10593, CK => CLK, Q => n52523,
                           QN => n1101);
   REGS_reg_117_27_inst : DFF_X1 port map( D => n10592, CK => CLK, Q => n52524,
                           QN => n1102);
   REGS_reg_117_26_inst : DFF_X1 port map( D => n10591, CK => CLK, Q => n52525,
                           QN => n1103);
   REGS_reg_117_25_inst : DFF_X1 port map( D => n10590, CK => CLK, Q => n52526,
                           QN => n1104);
   REGS_reg_117_24_inst : DFF_X1 port map( D => n10589, CK => CLK, Q => n52527,
                           QN => n1105);
   REGS_reg_116_31_inst : DFF_X1 port map( D => n10628, CK => CLK, Q => n52528,
                           QN => n1106);
   REGS_reg_116_30_inst : DFF_X1 port map( D => n10627, CK => CLK, Q => n52529,
                           QN => n1107);
   REGS_reg_116_29_inst : DFF_X1 port map( D => n10626, CK => CLK, Q => n52530,
                           QN => n1108);
   REGS_reg_116_28_inst : DFF_X1 port map( D => n10625, CK => CLK, Q => n52531,
                           QN => n1109);
   REGS_reg_116_27_inst : DFF_X1 port map( D => n10624, CK => CLK, Q => n52532,
                           QN => n1110);
   REGS_reg_116_26_inst : DFF_X1 port map( D => n10623, CK => CLK, Q => n52533,
                           QN => n1111);
   REGS_reg_116_25_inst : DFF_X1 port map( D => n10622, CK => CLK, Q => n52534,
                           QN => n1112);
   REGS_reg_116_24_inst : DFF_X1 port map( D => n10621, CK => CLK, Q => n52535,
                           QN => n1113);
   REGS_reg_114_24_inst : DFF_X1 port map( D => n10685, CK => CLK, Q => n1518, 
                           QN => n1114);
   REGS_reg_113_31_inst : DFF_X1 port map( D => n10724, CK => CLK, Q => n_1274,
                           QN => n1115);
   REGS_reg_113_30_inst : DFF_X1 port map( D => n10723, CK => CLK, Q => n_1275,
                           QN => n1116);
   REGS_reg_113_29_inst : DFF_X1 port map( D => n10722, CK => CLK, Q => n_1276,
                           QN => n1117);
   REGS_reg_113_28_inst : DFF_X1 port map( D => n10721, CK => CLK, Q => n_1277,
                           QN => n1118);
   REGS_reg_113_27_inst : DFF_X1 port map( D => n10720, CK => CLK, Q => n_1278,
                           QN => n1119);
   REGS_reg_113_26_inst : DFF_X1 port map( D => n10719, CK => CLK, Q => n_1279,
                           QN => n1120);
   REGS_reg_113_25_inst : DFF_X1 port map( D => n10718, CK => CLK, Q => n_1280,
                           QN => n1121);
   REGS_reg_113_24_inst : DFF_X1 port map( D => n10717, CK => CLK, Q => n_1281,
                           QN => n1122);
   REGS_reg_112_31_inst : DFF_X1 port map( D => n10756, CK => CLK, Q => n_1282,
                           QN => n1123);
   REGS_reg_112_30_inst : DFF_X1 port map( D => n10755, CK => CLK, Q => n_1283,
                           QN => n1124);
   REGS_reg_112_29_inst : DFF_X1 port map( D => n10754, CK => CLK, Q => n_1284,
                           QN => n1125);
   REGS_reg_112_28_inst : DFF_X1 port map( D => n10753, CK => CLK, Q => n_1285,
                           QN => n1126);
   REGS_reg_112_27_inst : DFF_X1 port map( D => n10752, CK => CLK, Q => n_1286,
                           QN => n1127);
   REGS_reg_112_26_inst : DFF_X1 port map( D => n10751, CK => CLK, Q => n_1287,
                           QN => n1128);
   REGS_reg_112_25_inst : DFF_X1 port map( D => n10750, CK => CLK, Q => n_1288,
                           QN => n1129);
   REGS_reg_112_24_inst : DFF_X1 port map( D => n10749, CK => CLK, Q => n_1289,
                           QN => n1130);
   REGS_reg_111_31_inst : DFF_X1 port map( D => n10788, CK => CLK, Q => n340, 
                           QN => n1131);
   REGS_reg_111_30_inst : DFF_X1 port map( D => n10787, CK => CLK, Q => n341, 
                           QN => n1132);
   REGS_reg_111_29_inst : DFF_X1 port map( D => n10786, CK => CLK, Q => n342, 
                           QN => n1133);
   REGS_reg_111_28_inst : DFF_X1 port map( D => n10785, CK => CLK, Q => n343, 
                           QN => n1134);
   REGS_reg_111_27_inst : DFF_X1 port map( D => n10784, CK => CLK, Q => n344, 
                           QN => n1135);
   REGS_reg_111_26_inst : DFF_X1 port map( D => n10783, CK => CLK, Q => n345, 
                           QN => n1136);
   REGS_reg_111_25_inst : DFF_X1 port map( D => n10782, CK => CLK, Q => n346, 
                           QN => n1137);
   REGS_reg_111_24_inst : DFF_X1 port map( D => n10781, CK => CLK, Q => n347, 
                           QN => n1138);
   REGS_reg_110_31_inst : DFF_X1 port map( D => n10820, CK => CLK, Q => n348, 
                           QN => n1139);
   REGS_reg_110_30_inst : DFF_X1 port map( D => n10819, CK => CLK, Q => n349, 
                           QN => n1140);
   REGS_reg_110_29_inst : DFF_X1 port map( D => n10818, CK => CLK, Q => n350, 
                           QN => n1141);
   REGS_reg_110_28_inst : DFF_X1 port map( D => n10817, CK => CLK, Q => n351, 
                           QN => n1142);
   REGS_reg_110_27_inst : DFF_X1 port map( D => n10816, CK => CLK, Q => n352, 
                           QN => n1143);
   REGS_reg_110_26_inst : DFF_X1 port map( D => n10815, CK => CLK, Q => n353, 
                           QN => n1144);
   REGS_reg_110_25_inst : DFF_X1 port map( D => n10814, CK => CLK, Q => n354, 
                           QN => n1145);
   REGS_reg_110_24_inst : DFF_X1 port map( D => n10813, CK => CLK, Q => n355, 
                           QN => n1146);
   REGS_reg_109_31_inst : DFF_X1 port map( D => n10852, CK => CLK, Q => n_1290,
                           QN => n1147);
   REGS_reg_109_30_inst : DFF_X1 port map( D => n10851, CK => CLK, Q => n_1291,
                           QN => n1148);
   REGS_reg_109_29_inst : DFF_X1 port map( D => n10850, CK => CLK, Q => n_1292,
                           QN => n1149);
   REGS_reg_109_28_inst : DFF_X1 port map( D => n10849, CK => CLK, Q => n_1293,
                           QN => n1150);
   REGS_reg_109_27_inst : DFF_X1 port map( D => n10848, CK => CLK, Q => n_1294,
                           QN => n1151);
   REGS_reg_109_26_inst : DFF_X1 port map( D => n10847, CK => CLK, Q => n_1295,
                           QN => n1152);
   REGS_reg_109_25_inst : DFF_X1 port map( D => n10846, CK => CLK, Q => n_1296,
                           QN => n1153);
   REGS_reg_109_24_inst : DFF_X1 port map( D => n10845, CK => CLK, Q => n_1297,
                           QN => n1154);
   REGS_reg_108_31_inst : DFF_X1 port map( D => n10884, CK => CLK, Q => n_1298,
                           QN => n1155);
   REGS_reg_108_30_inst : DFF_X1 port map( D => n10883, CK => CLK, Q => n_1299,
                           QN => n1156);
   REGS_reg_108_29_inst : DFF_X1 port map( D => n10882, CK => CLK, Q => n_1300,
                           QN => n1157);
   REGS_reg_108_28_inst : DFF_X1 port map( D => n10881, CK => CLK, Q => n_1301,
                           QN => n1158);
   REGS_reg_108_27_inst : DFF_X1 port map( D => n10880, CK => CLK, Q => n_1302,
                           QN => n1159);
   REGS_reg_108_26_inst : DFF_X1 port map( D => n10879, CK => CLK, Q => n_1303,
                           QN => n1160);
   REGS_reg_108_25_inst : DFF_X1 port map( D => n10878, CK => CLK, Q => n_1304,
                           QN => n1161);
   REGS_reg_108_24_inst : DFF_X1 port map( D => n10877, CK => CLK, Q => n_1305,
                           QN => n1162);
   REGS_reg_107_31_inst : DFF_X1 port map( D => n10916, CK => CLK, Q => n15343,
                           QN => n1163);
   REGS_reg_107_30_inst : DFF_X1 port map( D => n10915, CK => CLK, Q => n15330,
                           QN => n1164);
   REGS_reg_107_29_inst : DFF_X1 port map( D => n10914, CK => CLK, Q => n15329,
                           QN => n1165);
   REGS_reg_107_28_inst : DFF_X1 port map( D => n10913, CK => CLK, Q => n15328,
                           QN => n1166);
   REGS_reg_107_27_inst : DFF_X1 port map( D => n10912, CK => CLK, Q => n15327,
                           QN => n1167);
   REGS_reg_107_26_inst : DFF_X1 port map( D => n10911, CK => CLK, Q => n15326,
                           QN => n1168);
   REGS_reg_107_25_inst : DFF_X1 port map( D => n10910, CK => CLK, Q => n15325,
                           QN => n1169);
   REGS_reg_107_24_inst : DFF_X1 port map( D => n10909, CK => CLK, Q => n15324,
                           QN => n1170);
   REGS_reg_106_31_inst : DFF_X1 port map( D => n10948, CK => CLK, Q => n15323,
                           QN => n1171);
   REGS_reg_106_30_inst : DFF_X1 port map( D => n10947, CK => CLK, Q => n15322,
                           QN => n1172);
   REGS_reg_106_29_inst : DFF_X1 port map( D => n10946, CK => CLK, Q => n15321,
                           QN => n1173);
   REGS_reg_106_28_inst : DFF_X1 port map( D => n10945, CK => CLK, Q => n15320,
                           QN => n1174);
   REGS_reg_106_27_inst : DFF_X1 port map( D => n10944, CK => CLK, Q => n15319,
                           QN => n1175);
   REGS_reg_106_26_inst : DFF_X1 port map( D => n10943, CK => CLK, Q => n15318,
                           QN => n1176);
   REGS_reg_106_25_inst : DFF_X1 port map( D => n10942, CK => CLK, Q => n15317,
                           QN => n1177);
   REGS_reg_106_24_inst : DFF_X1 port map( D => n10941, CK => CLK, Q => n15316,
                           QN => n1178);
   REGS_reg_105_31_inst : DFF_X1 port map( D => n10980, CK => CLK, Q => n_1306,
                           QN => n1179);
   REGS_reg_105_30_inst : DFF_X1 port map( D => n10979, CK => CLK, Q => n_1307,
                           QN => n1180);
   REGS_reg_105_29_inst : DFF_X1 port map( D => n10978, CK => CLK, Q => n_1308,
                           QN => n1181);
   REGS_reg_105_28_inst : DFF_X1 port map( D => n10977, CK => CLK, Q => n_1309,
                           QN => n1182);
   REGS_reg_105_27_inst : DFF_X1 port map( D => n10976, CK => CLK, Q => n_1310,
                           QN => n1183);
   REGS_reg_105_26_inst : DFF_X1 port map( D => n10975, CK => CLK, Q => n_1311,
                           QN => n1184);
   REGS_reg_105_25_inst : DFF_X1 port map( D => n10974, CK => CLK, Q => n_1312,
                           QN => n1185);
   REGS_reg_105_24_inst : DFF_X1 port map( D => n10973, CK => CLK, Q => n_1313,
                           QN => n1186);
   REGS_reg_104_31_inst : DFF_X1 port map( D => n11012, CK => CLK, Q => n_1314,
                           QN => n1187);
   REGS_reg_104_30_inst : DFF_X1 port map( D => n11011, CK => CLK, Q => n_1315,
                           QN => n1188);
   REGS_reg_104_29_inst : DFF_X1 port map( D => n11010, CK => CLK, Q => n_1316,
                           QN => n1189);
   REGS_reg_104_28_inst : DFF_X1 port map( D => n11009, CK => CLK, Q => n_1317,
                           QN => n1190);
   REGS_reg_104_27_inst : DFF_X1 port map( D => n11008, CK => CLK, Q => n_1318,
                           QN => n1191);
   REGS_reg_104_26_inst : DFF_X1 port map( D => n11007, CK => CLK, Q => n_1319,
                           QN => n1192);
   REGS_reg_104_25_inst : DFF_X1 port map( D => n11006, CK => CLK, Q => n_1320,
                           QN => n1193);
   REGS_reg_104_24_inst : DFF_X1 port map( D => n11005, CK => CLK, Q => n_1321,
                           QN => n1194);
   REGS_reg_103_31_inst : DFF_X1 port map( D => n11044, CK => CLK, Q => n372, 
                           QN => n1195);
   REGS_reg_103_30_inst : DFF_X1 port map( D => n11043, CK => CLK, Q => n373, 
                           QN => n1196);
   REGS_reg_103_29_inst : DFF_X1 port map( D => n11042, CK => CLK, Q => n374, 
                           QN => n1197);
   REGS_reg_103_28_inst : DFF_X1 port map( D => n11041, CK => CLK, Q => n375, 
                           QN => n1198);
   REGS_reg_103_27_inst : DFF_X1 port map( D => n11040, CK => CLK, Q => n376, 
                           QN => n1199);
   REGS_reg_103_26_inst : DFF_X1 port map( D => n11039, CK => CLK, Q => n377, 
                           QN => n1200);
   REGS_reg_103_25_inst : DFF_X1 port map( D => n11038, CK => CLK, Q => n378, 
                           QN => n1201);
   REGS_reg_103_24_inst : DFF_X1 port map( D => n11037, CK => CLK, Q => n379, 
                           QN => n1202);
   REGS_reg_102_31_inst : DFF_X1 port map( D => n11076, CK => CLK, Q => n380, 
                           QN => n1203);
   REGS_reg_102_30_inst : DFF_X1 port map( D => n11075, CK => CLK, Q => n381, 
                           QN => n1204);
   REGS_reg_102_29_inst : DFF_X1 port map( D => n11074, CK => CLK, Q => n382, 
                           QN => n1205);
   REGS_reg_102_28_inst : DFF_X1 port map( D => n11073, CK => CLK, Q => n383, 
                           QN => n1206);
   REGS_reg_102_27_inst : DFF_X1 port map( D => n11072, CK => CLK, Q => n384, 
                           QN => n1207);
   REGS_reg_102_26_inst : DFF_X1 port map( D => n11071, CK => CLK, Q => n385, 
                           QN => n1208);
   REGS_reg_102_25_inst : DFF_X1 port map( D => n11070, CK => CLK, Q => n386, 
                           QN => n1209);
   REGS_reg_102_24_inst : DFF_X1 port map( D => n11069, CK => CLK, Q => n387, 
                           QN => n1210);
   REGS_reg_101_31_inst : DFF_X1 port map( D => n11108, CK => CLK, Q => n52584,
                           QN => n1211);
   REGS_reg_101_30_inst : DFF_X1 port map( D => n11107, CK => CLK, Q => n52585,
                           QN => n1212);
   REGS_reg_101_29_inst : DFF_X1 port map( D => n11106, CK => CLK, Q => n52586,
                           QN => n1213);
   REGS_reg_101_28_inst : DFF_X1 port map( D => n11105, CK => CLK, Q => n52587,
                           QN => n1214);
   REGS_reg_101_27_inst : DFF_X1 port map( D => n11104, CK => CLK, Q => n52588,
                           QN => n1215);
   REGS_reg_101_26_inst : DFF_X1 port map( D => n11103, CK => CLK, Q => n52589,
                           QN => n1216);
   REGS_reg_101_25_inst : DFF_X1 port map( D => n11102, CK => CLK, Q => n52590,
                           QN => n1217);
   REGS_reg_101_24_inst : DFF_X1 port map( D => n11101, CK => CLK, Q => n52591,
                           QN => n1218);
   REGS_reg_100_31_inst : DFF_X1 port map( D => n11140, CK => CLK, Q => n52592,
                           QN => n1219);
   REGS_reg_100_30_inst : DFF_X1 port map( D => n11139, CK => CLK, Q => n52593,
                           QN => n1220);
   REGS_reg_100_29_inst : DFF_X1 port map( D => n11138, CK => CLK, Q => n52594,
                           QN => n1221);
   REGS_reg_100_28_inst : DFF_X1 port map( D => n11137, CK => CLK, Q => n52595,
                           QN => n1222);
   REGS_reg_100_27_inst : DFF_X1 port map( D => n11136, CK => CLK, Q => n52596,
                           QN => n1223);
   REGS_reg_100_26_inst : DFF_X1 port map( D => n11135, CK => CLK, Q => n52597,
                           QN => n1224);
   REGS_reg_100_25_inst : DFF_X1 port map( D => n11134, CK => CLK, Q => n52598,
                           QN => n1225);
   REGS_reg_100_24_inst : DFF_X1 port map( D => n11133, CK => CLK, Q => n52599,
                           QN => n1226);
   REGS_reg_99_31_inst : DFF_X1 port map( D => n11172, CK => CLK, Q => n52600, 
                           QN => n1227);
   REGS_reg_99_30_inst : DFF_X1 port map( D => n11171, CK => CLK, Q => n52601, 
                           QN => n1228);
   REGS_reg_99_29_inst : DFF_X1 port map( D => n11170, CK => CLK, Q => n52602, 
                           QN => n1229);
   REGS_reg_99_28_inst : DFF_X1 port map( D => n11169, CK => CLK, Q => n52603, 
                           QN => n1230);
   REGS_reg_99_27_inst : DFF_X1 port map( D => n11168, CK => CLK, Q => n52604, 
                           QN => n1231);
   REGS_reg_99_26_inst : DFF_X1 port map( D => n11167, CK => CLK, Q => n52605, 
                           QN => n1232);
   REGS_reg_99_25_inst : DFF_X1 port map( D => n11166, CK => CLK, Q => n52606, 
                           QN => n1233);
   REGS_reg_99_24_inst : DFF_X1 port map( D => n11165, CK => CLK, Q => n52607, 
                           QN => n1234);
   REGS_reg_98_31_inst : DFF_X1 port map( D => n11204, CK => CLK, Q => n_1322, 
                           QN => n1235);
   REGS_reg_98_30_inst : DFF_X1 port map( D => n11203, CK => CLK, Q => n_1323, 
                           QN => n1236);
   REGS_reg_98_29_inst : DFF_X1 port map( D => n11202, CK => CLK, Q => n_1324, 
                           QN => n1237);
   REGS_reg_98_28_inst : DFF_X1 port map( D => n11201, CK => CLK, Q => n_1325, 
                           QN => n1238);
   REGS_reg_98_27_inst : DFF_X1 port map( D => n11200, CK => CLK, Q => n_1326, 
                           QN => n1239);
   REGS_reg_98_26_inst : DFF_X1 port map( D => n11199, CK => CLK, Q => n_1327, 
                           QN => n1240);
   REGS_reg_98_25_inst : DFF_X1 port map( D => n11198, CK => CLK, Q => n_1328, 
                           QN => n1241);
   REGS_reg_98_24_inst : DFF_X1 port map( D => n11197, CK => CLK, Q => n_1329, 
                           QN => n1242);
   REGS_reg_97_31_inst : DFF_X1 port map( D => n11236, CK => CLK, Q => n1567, 
                           QN => n1243);
   REGS_reg_97_30_inst : DFF_X1 port map( D => n11235, CK => CLK, Q => n1568, 
                           QN => n1244);
   REGS_reg_97_29_inst : DFF_X1 port map( D => n11234, CK => CLK, Q => n1569, 
                           QN => n1245);
   REGS_reg_97_28_inst : DFF_X1 port map( D => n11233, CK => CLK, Q => n1570, 
                           QN => n1246);
   REGS_reg_97_27_inst : DFF_X1 port map( D => n11232, CK => CLK, Q => n1571, 
                           QN => n1247);
   REGS_reg_97_26_inst : DFF_X1 port map( D => n11231, CK => CLK, Q => n1572, 
                           QN => n1248);
   REGS_reg_97_25_inst : DFF_X1 port map( D => n11230, CK => CLK, Q => n1573, 
                           QN => n1249);
   REGS_reg_97_24_inst : DFF_X1 port map( D => n11229, CK => CLK, Q => n1574, 
                           QN => n1250);
   REGS_reg_96_31_inst : DFF_X1 port map( D => n11268, CK => CLK, Q => n50964, 
                           QN => n1251);
   REGS_reg_96_30_inst : DFF_X1 port map( D => n11267, CK => CLK, Q => n50965, 
                           QN => n1252);
   REGS_reg_96_29_inst : DFF_X1 port map( D => n11266, CK => CLK, Q => n50966, 
                           QN => n1253);
   REGS_reg_96_28_inst : DFF_X1 port map( D => n11265, CK => CLK, Q => n50967, 
                           QN => n1254);
   REGS_reg_96_27_inst : DFF_X1 port map( D => n11264, CK => CLK, Q => n50968, 
                           QN => n1255);
   REGS_reg_96_26_inst : DFF_X1 port map( D => n11263, CK => CLK, Q => n50969, 
                           QN => n1256);
   REGS_reg_96_25_inst : DFF_X1 port map( D => n11262, CK => CLK, Q => n50970, 
                           QN => n1257);
   REGS_reg_96_24_inst : DFF_X1 port map( D => n11261, CK => CLK, Q => n50971, 
                           QN => n1258);
   REGS_reg_95_31_inst : DFF_X1 port map( D => n11300, CK => CLK, Q => n50932, 
                           QN => n136);
   REGS_reg_95_30_inst : DFF_X1 port map( D => n11299, CK => CLK, Q => n50933, 
                           QN => n137);
   REGS_reg_95_29_inst : DFF_X1 port map( D => n11298, CK => CLK, Q => n50934, 
                           QN => n138);
   REGS_reg_95_28_inst : DFF_X1 port map( D => n11297, CK => CLK, Q => n50935, 
                           QN => n139);
   REGS_reg_95_27_inst : DFF_X1 port map( D => n11296, CK => CLK, Q => n50936, 
                           QN => n140);
   REGS_reg_95_26_inst : DFF_X1 port map( D => n11295, CK => CLK, Q => n50937, 
                           QN => n141);
   REGS_reg_95_25_inst : DFF_X1 port map( D => n11294, CK => CLK, Q => n50938, 
                           QN => n142);
   REGS_reg_95_24_inst : DFF_X1 port map( D => n11293, CK => CLK, Q => n50939, 
                           QN => n143);
   REGS_reg_94_31_inst : DFF_X1 port map( D => n11332, CK => CLK, Q => n15370, 
                           QN => n144);
   REGS_reg_94_30_inst : DFF_X1 port map( D => n11331, CK => CLK, Q => n15369, 
                           QN => n145);
   REGS_reg_94_29_inst : DFF_X1 port map( D => n11330, CK => CLK, Q => n15368, 
                           QN => n146);
   REGS_reg_94_28_inst : DFF_X1 port map( D => n11329, CK => CLK, Q => n15367, 
                           QN => n147);
   REGS_reg_94_27_inst : DFF_X1 port map( D => n11328, CK => CLK, Q => n15366, 
                           QN => n148);
   REGS_reg_94_26_inst : DFF_X1 port map( D => n11327, CK => CLK, Q => n15365, 
                           QN => n149);
   REGS_reg_94_25_inst : DFF_X1 port map( D => n11326, CK => CLK, Q => n15364, 
                           QN => n150);
   REGS_reg_94_24_inst : DFF_X1 port map( D => n11325, CK => CLK, Q => n15363, 
                           QN => n151);
   REGS_reg_93_31_inst : DFF_X1 port map( D => n11364, CK => CLK, Q => n_1330, 
                           QN => n152);
   REGS_reg_93_30_inst : DFF_X1 port map( D => n11363, CK => CLK, Q => n_1331, 
                           QN => n153);
   REGS_reg_93_29_inst : DFF_X1 port map( D => n11362, CK => CLK, Q => n_1332, 
                           QN => n154);
   REGS_reg_93_28_inst : DFF_X1 port map( D => n11361, CK => CLK, Q => n_1333, 
                           QN => n155);
   REGS_reg_93_27_inst : DFF_X1 port map( D => n11360, CK => CLK, Q => n_1334, 
                           QN => n156);
   REGS_reg_93_26_inst : DFF_X1 port map( D => n11359, CK => CLK, Q => n_1335, 
                           QN => n157);
   REGS_reg_93_25_inst : DFF_X1 port map( D => n11358, CK => CLK, Q => n_1336, 
                           QN => n158);
   REGS_reg_93_24_inst : DFF_X1 port map( D => n11357, CK => CLK, Q => n_1337, 
                           QN => n159);
   REGS_reg_92_31_inst : DFF_X1 port map( D => n11396, CK => CLK, Q => n15482, 
                           QN => n213);
   REGS_reg_92_30_inst : DFF_X1 port map( D => n11395, CK => CLK, Q => n15481, 
                           QN => n214);
   REGS_reg_92_29_inst : DFF_X1 port map( D => n11394, CK => CLK, Q => n15480, 
                           QN => n215);
   REGS_reg_92_28_inst : DFF_X1 port map( D => n11393, CK => CLK, Q => n15479, 
                           QN => n216);
   REGS_reg_92_27_inst : DFF_X1 port map( D => n11392, CK => CLK, Q => n15478, 
                           QN => n217);
   REGS_reg_92_26_inst : DFF_X1 port map( D => n11391, CK => CLK, Q => n15477, 
                           QN => n218);
   REGS_reg_92_25_inst : DFF_X1 port map( D => n11390, CK => CLK, Q => n15476, 
                           QN => n219);
   REGS_reg_92_24_inst : DFF_X1 port map( D => n11389, CK => CLK, Q => n15475, 
                           QN => n220);
   REGS_reg_91_31_inst : DFF_X1 port map( D => n11428, CK => CLK, Q => n15474, 
                           QN => n221);
   REGS_reg_91_30_inst : DFF_X1 port map( D => n11427, CK => CLK, Q => n15473, 
                           QN => n222);
   REGS_reg_91_29_inst : DFF_X1 port map( D => n11426, CK => CLK, Q => n15472, 
                           QN => n223);
   REGS_reg_91_28_inst : DFF_X1 port map( D => n11425, CK => CLK, Q => n15471, 
                           QN => n224);
   REGS_reg_91_27_inst : DFF_X1 port map( D => n11424, CK => CLK, Q => n15470, 
                           QN => n225);
   REGS_reg_91_26_inst : DFF_X1 port map( D => n11423, CK => CLK, Q => n15469, 
                           QN => n226);
   REGS_reg_91_25_inst : DFF_X1 port map( D => n11422, CK => CLK, Q => n15468, 
                           QN => n227);
   REGS_reg_91_24_inst : DFF_X1 port map( D => n11421, CK => CLK, Q => n15467, 
                           QN => n228);
   REGS_reg_90_31_inst : DFF_X1 port map( D => n11460, CK => CLK, Q => n_1338, 
                           QN => n4012);
   REGS_reg_90_30_inst : DFF_X1 port map( D => n11459, CK => CLK, Q => n_1339, 
                           QN => n4013);
   REGS_reg_90_29_inst : DFF_X1 port map( D => n11458, CK => CLK, Q => n_1340, 
                           QN => n4014);
   REGS_reg_90_28_inst : DFF_X1 port map( D => n11457, CK => CLK, Q => n_1341, 
                           QN => n4015);
   REGS_reg_90_27_inst : DFF_X1 port map( D => n11456, CK => CLK, Q => n_1342, 
                           QN => n4016);
   REGS_reg_90_26_inst : DFF_X1 port map( D => n11455, CK => CLK, Q => n_1343, 
                           QN => n4017);
   REGS_reg_90_25_inst : DFF_X1 port map( D => n11454, CK => CLK, Q => n_1344, 
                           QN => n4018);
   REGS_reg_90_24_inst : DFF_X1 port map( D => n11453, CK => CLK, Q => n_1345, 
                           QN => n4019);
   REGS_reg_89_31_inst : DFF_X1 port map( D => n11492, CK => CLK, Q => n_1346, 
                           QN => n4020);
   REGS_reg_89_30_inst : DFF_X1 port map( D => n11491, CK => CLK, Q => n_1347, 
                           QN => n4021);
   REGS_reg_89_29_inst : DFF_X1 port map( D => n11490, CK => CLK, Q => n_1348, 
                           QN => n4022);
   REGS_reg_89_28_inst : DFF_X1 port map( D => n11489, CK => CLK, Q => n_1349, 
                           QN => n4023);
   REGS_reg_89_27_inst : DFF_X1 port map( D => n11488, CK => CLK, Q => n_1350, 
                           QN => n4024);
   REGS_reg_89_26_inst : DFF_X1 port map( D => n11487, CK => CLK, Q => n_1351, 
                           QN => n4025);
   REGS_reg_89_25_inst : DFF_X1 port map( D => n11486, CK => CLK, Q => n_1352, 
                           QN => n4026);
   REGS_reg_89_24_inst : DFF_X1 port map( D => n11485, CK => CLK, Q => n_1353, 
                           QN => n4027);
   REGS_reg_88_31_inst : DFF_X1 port map( D => n11524, CK => CLK, Q => n51712, 
                           QN => n229);
   REGS_reg_88_30_inst : DFF_X1 port map( D => n11523, CK => CLK, Q => n51713, 
                           QN => n230);
   REGS_reg_88_29_inst : DFF_X1 port map( D => n11522, CK => CLK, Q => n51714, 
                           QN => n231);
   REGS_reg_88_28_inst : DFF_X1 port map( D => n11521, CK => CLK, Q => n51715, 
                           QN => n232);
   REGS_reg_88_27_inst : DFF_X1 port map( D => n11520, CK => CLK, Q => n51716, 
                           QN => n233);
   REGS_reg_88_26_inst : DFF_X1 port map( D => n11519, CK => CLK, Q => n51717, 
                           QN => n234);
   REGS_reg_88_25_inst : DFF_X1 port map( D => n11518, CK => CLK, Q => n51718, 
                           QN => n235);
   REGS_reg_88_24_inst : DFF_X1 port map( D => n11517, CK => CLK, Q => n51719, 
                           QN => n236);
   REGS_reg_87_31_inst : DFF_X1 port map( D => n11556, CK => CLK, Q => n51720, 
                           QN => n237);
   REGS_reg_87_30_inst : DFF_X1 port map( D => n11555, CK => CLK, Q => n51721, 
                           QN => n238);
   REGS_reg_87_29_inst : DFF_X1 port map( D => n11554, CK => CLK, Q => n51722, 
                           QN => n239);
   REGS_reg_87_28_inst : DFF_X1 port map( D => n11553, CK => CLK, Q => n51723, 
                           QN => n240);
   REGS_reg_87_27_inst : DFF_X1 port map( D => n11552, CK => CLK, Q => n51724, 
                           QN => n241);
   REGS_reg_87_26_inst : DFF_X1 port map( D => n11551, CK => CLK, Q => n51725, 
                           QN => n242);
   REGS_reg_87_25_inst : DFF_X1 port map( D => n11550, CK => CLK, Q => n51726, 
                           QN => n243);
   REGS_reg_87_24_inst : DFF_X1 port map( D => n11549, CK => CLK, Q => n51727, 
                           QN => n244);
   REGS_reg_86_31_inst : DFF_X1 port map( D => n11588, CK => CLK, Q => n_1354, 
                           QN => n245);
   REGS_reg_86_30_inst : DFF_X1 port map( D => n11587, CK => CLK, Q => n_1355, 
                           QN => n246);
   REGS_reg_86_29_inst : DFF_X1 port map( D => n11586, CK => CLK, Q => n_1356, 
                           QN => n247);
   REGS_reg_86_28_inst : DFF_X1 port map( D => n11585, CK => CLK, Q => n_1357, 
                           QN => n248);
   REGS_reg_86_27_inst : DFF_X1 port map( D => n11584, CK => CLK, Q => n_1358, 
                           QN => n249);
   REGS_reg_86_26_inst : DFF_X1 port map( D => n11583, CK => CLK, Q => n_1359, 
                           QN => n250);
   REGS_reg_86_25_inst : DFF_X1 port map( D => n11582, CK => CLK, Q => n_1360, 
                           QN => n251);
   REGS_reg_86_24_inst : DFF_X1 port map( D => n11581, CK => CLK, Q => n_1361, 
                           QN => n252);
   REGS_reg_85_31_inst : DFF_X1 port map( D => n11620, CK => CLK, Q => n_1362, 
                           QN => n253);
   REGS_reg_85_30_inst : DFF_X1 port map( D => n11619, CK => CLK, Q => n_1363, 
                           QN => n254);
   REGS_reg_85_29_inst : DFF_X1 port map( D => n11618, CK => CLK, Q => n_1364, 
                           QN => n255);
   REGS_reg_85_28_inst : DFF_X1 port map( D => n11617, CK => CLK, Q => n_1365, 
                           QN => n256);
   REGS_reg_85_27_inst : DFF_X1 port map( D => n11616, CK => CLK, Q => n_1366, 
                           QN => n257);
   REGS_reg_85_26_inst : DFF_X1 port map( D => n11615, CK => CLK, Q => n_1367, 
                           QN => n258);
   REGS_reg_85_25_inst : DFF_X1 port map( D => n11614, CK => CLK, Q => n_1368, 
                           QN => n259);
   REGS_reg_85_24_inst : DFF_X1 port map( D => n11613, CK => CLK, Q => n_1369, 
                           QN => n260);
   REGS_reg_84_31_inst : DFF_X1 port map( D => n11652, CK => CLK, Q => n52656, 
                           QN => n261);
   REGS_reg_84_30_inst : DFF_X1 port map( D => n11651, CK => CLK, Q => n52657, 
                           QN => n262);
   REGS_reg_84_29_inst : DFF_X1 port map( D => n11650, CK => CLK, Q => n52658, 
                           QN => n263);
   REGS_reg_84_28_inst : DFF_X1 port map( D => n11649, CK => CLK, Q => n52659, 
                           QN => n264);
   REGS_reg_84_27_inst : DFF_X1 port map( D => n11648, CK => CLK, Q => n52660, 
                           QN => n265);
   REGS_reg_84_26_inst : DFF_X1 port map( D => n11647, CK => CLK, Q => n52661, 
                           QN => n266);
   REGS_reg_84_25_inst : DFF_X1 port map( D => n11646, CK => CLK, Q => n52662, 
                           QN => n267);
   REGS_reg_84_24_inst : DFF_X1 port map( D => n11645, CK => CLK, Q => n52663, 
                           QN => n268);
   REGS_reg_81_31_inst : DFF_X1 port map( D => n11748, CK => CLK, Q => n_1370, 
                           QN => n269);
   REGS_reg_81_30_inst : DFF_X1 port map( D => n11747, CK => CLK, Q => n_1371, 
                           QN => n270);
   REGS_reg_81_29_inst : DFF_X1 port map( D => n11746, CK => CLK, Q => n_1372, 
                           QN => n271);
   REGS_reg_81_28_inst : DFF_X1 port map( D => n11745, CK => CLK, Q => n_1373, 
                           QN => n272);
   REGS_reg_81_27_inst : DFF_X1 port map( D => n11744, CK => CLK, Q => n_1374, 
                           QN => n273);
   REGS_reg_81_26_inst : DFF_X1 port map( D => n11743, CK => CLK, Q => n_1375, 
                           QN => n274);
   REGS_reg_81_25_inst : DFF_X1 port map( D => n11742, CK => CLK, Q => n_1376, 
                           QN => n275);
   REGS_reg_81_24_inst : DFF_X1 port map( D => n11741, CK => CLK, Q => n_1377, 
                           QN => n276);
   REGS_reg_80_31_inst : DFF_X1 port map( D => n11780, CK => CLK, Q => n1639, 
                           QN => n277);
   REGS_reg_80_30_inst : DFF_X1 port map( D => n11779, CK => CLK, Q => n1640, 
                           QN => n278);
   REGS_reg_80_29_inst : DFF_X1 port map( D => n11778, CK => CLK, Q => n1641, 
                           QN => n279);
   REGS_reg_80_28_inst : DFF_X1 port map( D => n11777, CK => CLK, Q => n1642, 
                           QN => n280);
   REGS_reg_80_27_inst : DFF_X1 port map( D => n11776, CK => CLK, Q => n1643, 
                           QN => n281);
   REGS_reg_80_26_inst : DFF_X1 port map( D => n11775, CK => CLK, Q => n1644, 
                           QN => n282);
   REGS_reg_80_25_inst : DFF_X1 port map( D => n11774, CK => CLK, Q => n1645, 
                           QN => n283);
   REGS_reg_80_24_inst : DFF_X1 port map( D => n11773, CK => CLK, Q => n1646, 
                           QN => n284);
   REGS_reg_79_31_inst : DFF_X1 port map( D => n11812, CK => CLK, Q => n51728, 
                           QN => n285);
   REGS_reg_79_30_inst : DFF_X1 port map( D => n11811, CK => CLK, Q => n51729, 
                           QN => n286);
   REGS_reg_79_29_inst : DFF_X1 port map( D => n11810, CK => CLK, Q => n51730, 
                           QN => n287);
   REGS_reg_79_28_inst : DFF_X1 port map( D => n11809, CK => CLK, Q => n51731, 
                           QN => n288);
   REGS_reg_79_27_inst : DFF_X1 port map( D => n11808, CK => CLK, Q => n51732, 
                           QN => n289);
   REGS_reg_79_26_inst : DFF_X1 port map( D => n11807, CK => CLK, Q => n51733, 
                           QN => n290);
   REGS_reg_79_25_inst : DFF_X1 port map( D => n11806, CK => CLK, Q => n51734, 
                           QN => n291);
   REGS_reg_79_24_inst : DFF_X1 port map( D => n11805, CK => CLK, Q => n51735, 
                           QN => n292);
   REGS_reg_78_31_inst : DFF_X1 port map( D => n11844, CK => CLK, Q => n51736, 
                           QN => n293);
   REGS_reg_78_30_inst : DFF_X1 port map( D => n11843, CK => CLK, Q => n51737, 
                           QN => n294);
   REGS_reg_78_29_inst : DFF_X1 port map( D => n11842, CK => CLK, Q => n51738, 
                           QN => n295);
   REGS_reg_78_28_inst : DFF_X1 port map( D => n11841, CK => CLK, Q => n51739, 
                           QN => n296);
   REGS_reg_78_27_inst : DFF_X1 port map( D => n11840, CK => CLK, Q => n51740, 
                           QN => n297);
   REGS_reg_78_26_inst : DFF_X1 port map( D => n11839, CK => CLK, Q => n51741, 
                           QN => n298);
   REGS_reg_78_25_inst : DFF_X1 port map( D => n11838, CK => CLK, Q => n51742, 
                           QN => n299);
   REGS_reg_78_24_inst : DFF_X1 port map( D => n11837, CK => CLK, Q => n51743, 
                           QN => n300);
   REGS_reg_77_31_inst : DFF_X1 port map( D => n11876, CK => CLK, Q => n_1378, 
                           QN => n4044);
   REGS_reg_77_30_inst : DFF_X1 port map( D => n11875, CK => CLK, Q => n_1379, 
                           QN => n4045);
   REGS_reg_77_29_inst : DFF_X1 port map( D => n11874, CK => CLK, Q => n_1380, 
                           QN => n4046);
   REGS_reg_77_28_inst : DFF_X1 port map( D => n11873, CK => CLK, Q => n_1381, 
                           QN => n4047);
   REGS_reg_77_27_inst : DFF_X1 port map( D => n11872, CK => CLK, Q => n_1382, 
                           QN => n4048);
   REGS_reg_77_26_inst : DFF_X1 port map( D => n11871, CK => CLK, Q => n_1383, 
                           QN => n4049);
   REGS_reg_77_25_inst : DFF_X1 port map( D => n11870, CK => CLK, Q => n_1384, 
                           QN => n4050);
   REGS_reg_77_24_inst : DFF_X1 port map( D => n11869, CK => CLK, Q => n_1385, 
                           QN => n4051);
   REGS_reg_76_31_inst : DFF_X1 port map( D => n11908, CK => CLK, Q => n_1386, 
                           QN => n4052);
   REGS_reg_76_30_inst : DFF_X1 port map( D => n11907, CK => CLK, Q => n_1387, 
                           QN => n4053);
   REGS_reg_76_29_inst : DFF_X1 port map( D => n11906, CK => CLK, Q => n_1388, 
                           QN => n4054);
   REGS_reg_76_28_inst : DFF_X1 port map( D => n11905, CK => CLK, Q => n_1389, 
                           QN => n4055);
   REGS_reg_76_27_inst : DFF_X1 port map( D => n11904, CK => CLK, Q => n_1390, 
                           QN => n4056);
   REGS_reg_76_26_inst : DFF_X1 port map( D => n11903, CK => CLK, Q => n_1391, 
                           QN => n4057);
   REGS_reg_76_25_inst : DFF_X1 port map( D => n11902, CK => CLK, Q => n_1392, 
                           QN => n4058);
   REGS_reg_76_24_inst : DFF_X1 port map( D => n11901, CK => CLK, Q => n_1393, 
                           QN => n4059);
   REGS_reg_75_31_inst : DFF_X1 port map( D => n11940, CK => CLK, Q => n436, QN
                           => n301);
   REGS_reg_75_30_inst : DFF_X1 port map( D => n11939, CK => CLK, Q => n437, QN
                           => n302);
   REGS_reg_75_29_inst : DFF_X1 port map( D => n11938, CK => CLK, Q => n438, QN
                           => n303);
   REGS_reg_75_28_inst : DFF_X1 port map( D => n11937, CK => CLK, Q => n439, QN
                           => n304);
   REGS_reg_75_27_inst : DFF_X1 port map( D => n11936, CK => CLK, Q => n440, QN
                           => n305);
   REGS_reg_75_26_inst : DFF_X1 port map( D => n11935, CK => CLK, Q => n441, QN
                           => n306);
   REGS_reg_75_25_inst : DFF_X1 port map( D => n11934, CK => CLK, Q => n442, QN
                           => n307);
   REGS_reg_75_24_inst : DFF_X1 port map( D => n11933, CK => CLK, Q => n443, QN
                           => n308);
   REGS_reg_74_31_inst : DFF_X1 port map( D => n11972, CK => CLK, Q => n444, QN
                           => n309);
   REGS_reg_74_30_inst : DFF_X1 port map( D => n11971, CK => CLK, Q => n445, QN
                           => n310);
   REGS_reg_74_29_inst : DFF_X1 port map( D => n11970, CK => CLK, Q => n446, QN
                           => n311);
   REGS_reg_74_28_inst : DFF_X1 port map( D => n11969, CK => CLK, Q => n447, QN
                           => n312);
   REGS_reg_74_27_inst : DFF_X1 port map( D => n11968, CK => CLK, Q => n448, QN
                           => n313);
   REGS_reg_74_26_inst : DFF_X1 port map( D => n11967, CK => CLK, Q => n449, QN
                           => n314);
   REGS_reg_74_25_inst : DFF_X1 port map( D => n11966, CK => CLK, Q => n450, QN
                           => n315);
   REGS_reg_74_24_inst : DFF_X1 port map( D => n11965, CK => CLK, Q => n451, QN
                           => n316);
   REGS_reg_73_31_inst : DFF_X1 port map( D => n12004, CK => CLK, Q => n_1394, 
                           QN => n317);
   REGS_reg_73_30_inst : DFF_X1 port map( D => n12003, CK => CLK, Q => n_1395, 
                           QN => n318);
   REGS_reg_73_29_inst : DFF_X1 port map( D => n12002, CK => CLK, Q => n_1396, 
                           QN => n319);
   REGS_reg_73_28_inst : DFF_X1 port map( D => n12001, CK => CLK, Q => n_1397, 
                           QN => n320);
   REGS_reg_73_27_inst : DFF_X1 port map( D => n12000, CK => CLK, Q => n_1398, 
                           QN => n321);
   REGS_reg_73_26_inst : DFF_X1 port map( D => n11999, CK => CLK, Q => n_1399, 
                           QN => n322);
   REGS_reg_73_25_inst : DFF_X1 port map( D => n11998, CK => CLK, Q => n_1400, 
                           QN => n323);
   REGS_reg_73_24_inst : DFF_X1 port map( D => n11997, CK => CLK, Q => n_1401, 
                           QN => n324);
   REGS_reg_72_31_inst : DFF_X1 port map( D => n12036, CK => CLK, Q => n_1402, 
                           QN => n325);
   REGS_reg_72_30_inst : DFF_X1 port map( D => n12035, CK => CLK, Q => n_1403, 
                           QN => n326);
   REGS_reg_72_29_inst : DFF_X1 port map( D => n12034, CK => CLK, Q => n_1404, 
                           QN => n327);
   REGS_reg_72_28_inst : DFF_X1 port map( D => n12033, CK => CLK, Q => n_1405, 
                           QN => n328);
   REGS_reg_72_27_inst : DFF_X1 port map( D => n12032, CK => CLK, Q => n_1406, 
                           QN => n329);
   REGS_reg_72_26_inst : DFF_X1 port map( D => n12031, CK => CLK, Q => n_1407, 
                           QN => n330);
   REGS_reg_72_25_inst : DFF_X1 port map( D => n12030, CK => CLK, Q => n_1408, 
                           QN => n331);
   REGS_reg_72_24_inst : DFF_X1 port map( D => n12029, CK => CLK, Q => n_1409, 
                           QN => n332);
   REGS_reg_71_31_inst : DFF_X1 port map( D => n12068, CK => CLK, Q => n51760, 
                           QN => n333);
   REGS_reg_71_30_inst : DFF_X1 port map( D => n12067, CK => CLK, Q => n51761, 
                           QN => n334);
   REGS_reg_71_29_inst : DFF_X1 port map( D => n12066, CK => CLK, Q => n51762, 
                           QN => n335);
   REGS_reg_71_28_inst : DFF_X1 port map( D => n12065, CK => CLK, Q => n51763, 
                           QN => n336);
   REGS_reg_71_27_inst : DFF_X1 port map( D => n12064, CK => CLK, Q => n51764, 
                           QN => n337);
   REGS_reg_71_26_inst : DFF_X1 port map( D => n12063, CK => CLK, Q => n51765, 
                           QN => n338);
   REGS_reg_71_25_inst : DFF_X1 port map( D => n12062, CK => CLK, Q => n51766, 
                           QN => n339);
   REGS_reg_71_24_inst : DFF_X1 port map( D => n12061, CK => CLK, Q => n51767, 
                           QN => n356);
   REGS_reg_70_31_inst : DFF_X1 port map( D => n12100, CK => CLK, Q => n51768, 
                           QN => n357);
   REGS_reg_70_30_inst : DFF_X1 port map( D => n12099, CK => CLK, Q => n51769, 
                           QN => n358);
   REGS_reg_70_29_inst : DFF_X1 port map( D => n12098, CK => CLK, Q => n51770, 
                           QN => n359);
   REGS_reg_70_28_inst : DFF_X1 port map( D => n12097, CK => CLK, Q => n51771, 
                           QN => n360);
   REGS_reg_70_27_inst : DFF_X1 port map( D => n12096, CK => CLK, Q => n51772, 
                           QN => n361);
   REGS_reg_70_26_inst : DFF_X1 port map( D => n12095, CK => CLK, Q => n51773, 
                           QN => n362);
   REGS_reg_70_25_inst : DFF_X1 port map( D => n12094, CK => CLK, Q => n51774, 
                           QN => n363);
   REGS_reg_70_24_inst : DFF_X1 port map( D => n12093, CK => CLK, Q => n51775, 
                           QN => n364);
   REGS_reg_69_31_inst : DFF_X1 port map( D => n12132, CK => CLK, Q => n16356, 
                           QN => n4060);
   REGS_reg_69_30_inst : DFF_X1 port map( D => n12131, CK => CLK, Q => n16355, 
                           QN => n4061);
   REGS_reg_69_29_inst : DFF_X1 port map( D => n12130, CK => CLK, Q => n16354, 
                           QN => n4062);
   REGS_reg_69_28_inst : DFF_X1 port map( D => n12129, CK => CLK, Q => n16353, 
                           QN => n4063);
   REGS_reg_69_27_inst : DFF_X1 port map( D => n12128, CK => CLK, Q => n16352, 
                           QN => n4064);
   REGS_reg_69_26_inst : DFF_X1 port map( D => n12127, CK => CLK, Q => n16351, 
                           QN => n4065);
   REGS_reg_69_25_inst : DFF_X1 port map( D => n12126, CK => CLK, Q => n16350, 
                           QN => n4066);
   REGS_reg_69_24_inst : DFF_X1 port map( D => n12125, CK => CLK, Q => n16349, 
                           QN => n4067);
   REGS_reg_68_31_inst : DFF_X1 port map( D => n12164, CK => CLK, Q => n16348, 
                           QN => n4068);
   REGS_reg_68_30_inst : DFF_X1 port map( D => n12163, CK => CLK, Q => n16347, 
                           QN => n4069);
   REGS_reg_68_29_inst : DFF_X1 port map( D => n12162, CK => CLK, Q => n16346, 
                           QN => n4070);
   REGS_reg_68_28_inst : DFF_X1 port map( D => n12161, CK => CLK, Q => n16345, 
                           QN => n4071);
   REGS_reg_68_27_inst : DFF_X1 port map( D => n12160, CK => CLK, Q => n16344, 
                           QN => n4072);
   REGS_reg_68_26_inst : DFF_X1 port map( D => n12159, CK => CLK, Q => n16343, 
                           QN => n4073);
   REGS_reg_68_25_inst : DFF_X1 port map( D => n12158, CK => CLK, Q => n16342, 
                           QN => n4074);
   REGS_reg_68_24_inst : DFF_X1 port map( D => n12157, CK => CLK, Q => n16341, 
                           QN => n4075);
   REGS_reg_64_31_inst : DFF_X1 port map( D => n12292, CK => CLK, Q => n_1410, 
                           QN => n365);
   REGS_reg_64_30_inst : DFF_X1 port map( D => n12291, CK => CLK, Q => n_1411, 
                           QN => n366);
   REGS_reg_64_29_inst : DFF_X1 port map( D => n12290, CK => CLK, Q => n_1412, 
                           QN => n367);
   REGS_reg_64_28_inst : DFF_X1 port map( D => n12289, CK => CLK, Q => n_1413, 
                           QN => n368);
   REGS_reg_64_27_inst : DFF_X1 port map( D => n12288, CK => CLK, Q => n_1414, 
                           QN => n369);
   REGS_reg_64_26_inst : DFF_X1 port map( D => n12287, CK => CLK, Q => n_1415, 
                           QN => n370);
   REGS_reg_64_25_inst : DFF_X1 port map( D => n12286, CK => CLK, Q => n_1416, 
                           QN => n371);
   REGS_reg_64_24_inst : DFF_X1 port map( D => n12285, CK => CLK, Q => n_1417, 
                           QN => n388);
   REGS_reg_134_31_inst : DFF_X1 port map( D => n10052, CK => CLK, Q => n51776,
                           QN => n1259);
   REGS_reg_134_30_inst : DFF_X1 port map( D => n10051, CK => CLK, Q => n51777,
                           QN => n1260);
   REGS_reg_134_29_inst : DFF_X1 port map( D => n10050, CK => CLK, Q => n51778,
                           QN => n1261);
   REGS_reg_134_28_inst : DFF_X1 port map( D => n10049, CK => CLK, Q => n51779,
                           QN => n1262);
   REGS_reg_134_27_inst : DFF_X1 port map( D => n10048, CK => CLK, Q => n51780,
                           QN => n1263);
   REGS_reg_134_26_inst : DFF_X1 port map( D => n10047, CK => CLK, Q => n51781,
                           QN => n1264);
   REGS_reg_134_25_inst : DFF_X1 port map( D => n10046, CK => CLK, Q => n51782,
                           QN => n1265);
   REGS_reg_134_24_inst : DFF_X1 port map( D => n10045, CK => CLK, Q => n51783,
                           QN => n1266);
   REGS_reg_135_31_inst : DFF_X1 port map( D => n10020, CK => CLK, Q => n52760,
                           QN => n1267);
   REGS_reg_135_30_inst : DFF_X1 port map( D => n10019, CK => CLK, Q => n52761,
                           QN => n1268);
   REGS_reg_135_29_inst : DFF_X1 port map( D => n10018, CK => CLK, Q => n52762,
                           QN => n1269);
   REGS_reg_135_28_inst : DFF_X1 port map( D => n10017, CK => CLK, Q => n52763,
                           QN => n1270);
   REGS_reg_135_27_inst : DFF_X1 port map( D => n10016, CK => CLK, Q => n52764,
                           QN => n1271);
   REGS_reg_135_26_inst : DFF_X1 port map( D => n10015, CK => CLK, Q => n52765,
                           QN => n1272);
   REGS_reg_135_25_inst : DFF_X1 port map( D => n10014, CK => CLK, Q => n52766,
                           QN => n1273);
   REGS_reg_135_24_inst : DFF_X1 port map( D => n10013, CK => CLK, Q => n52767,
                           QN => n1274);
   REGS_reg_135_23_inst : DFF_X1 port map( D => n10012, CK => CLK, Q => n52768,
                           QN => n1275);
   REGS_reg_135_22_inst : DFF_X1 port map( D => n10011, CK => CLK, Q => n52769,
                           QN => n1276);
   REGS_reg_135_21_inst : DFF_X1 port map( D => n10010, CK => CLK, Q => n52770,
                           QN => n1277);
   REGS_reg_135_20_inst : DFF_X1 port map( D => n10009, CK => CLK, Q => n52771,
                           QN => n1278);
   REGS_reg_135_19_inst : DFF_X1 port map( D => n10008, CK => CLK, Q => n52772,
                           QN => n1279);
   REGS_reg_135_10_inst : DFF_X1 port map( D => n9999, CK => CLK, Q => n52773, 
                           QN => n1280);
   REGS_reg_135_9_inst : DFF_X1 port map( D => n9998, CK => CLK, Q => n52774, 
                           QN => n1281);
   REGS_reg_135_8_inst : DFF_X1 port map( D => n9997, CK => CLK, Q => n52775, 
                           QN => n1282);
   REGS_reg_135_7_inst : DFF_X1 port map( D => n9996, CK => CLK, Q => n52776, 
                           QN => n1283);
   REGS_reg_135_6_inst : DFF_X1 port map( D => n9995, CK => CLK, Q => n52777, 
                           QN => n1284);
   REGS_reg_135_5_inst : DFF_X1 port map( D => n9994, CK => CLK, Q => n52778, 
                           QN => n1285);
   REGS_reg_135_4_inst : DFF_X1 port map( D => n9993, CK => CLK, Q => n52779, 
                           QN => n1286);
   REGS_reg_135_3_inst : DFF_X1 port map( D => n9992, CK => CLK, Q => n52780, 
                           QN => n1287);
   REGS_reg_135_2_inst : DFF_X1 port map( D => n9991, CK => CLK, Q => n52781, 
                           QN => n1288);
   REGS_reg_135_1_inst : DFF_X1 port map( D => n9990, CK => CLK, Q => n52782, 
                           QN => n1289);
   REGS_reg_135_0_inst : DFF_X1 port map( D => n9989, CK => CLK, Q => n52783, 
                           QN => n1290);
   REGS_reg_133_23_inst : DFF_X1 port map( D => n10076, CK => CLK, Q => n52784,
                           QN => n1291);
   REGS_reg_133_22_inst : DFF_X1 port map( D => n10075, CK => CLK, Q => n52785,
                           QN => n1292);
   REGS_reg_133_21_inst : DFF_X1 port map( D => n10074, CK => CLK, Q => n52786,
                           QN => n1293);
   REGS_reg_133_20_inst : DFF_X1 port map( D => n10073, CK => CLK, Q => n52787,
                           QN => n1294);
   REGS_reg_133_19_inst : DFF_X1 port map( D => n10072, CK => CLK, Q => n52788,
                           QN => n1295);
   REGS_reg_133_18_inst : DFF_X1 port map( D => n10071, CK => CLK, Q => n52789,
                           QN => n1296);
   REGS_reg_133_17_inst : DFF_X1 port map( D => n10070, CK => CLK, Q => n52790,
                           QN => n1297);
   REGS_reg_133_16_inst : DFF_X1 port map( D => n10069, CK => CLK, Q => n52791,
                           QN => n1298);
   REGS_reg_133_15_inst : DFF_X1 port map( D => n10068, CK => CLK, Q => n52792,
                           QN => n1299);
   REGS_reg_133_14_inst : DFF_X1 port map( D => n10067, CK => CLK, Q => n52793,
                           QN => n1300);
   REGS_reg_133_13_inst : DFF_X1 port map( D => n10066, CK => CLK, Q => n52794,
                           QN => n1301);
   REGS_reg_133_12_inst : DFF_X1 port map( D => n10065, CK => CLK, Q => n52795,
                           QN => n1302);
   REGS_reg_133_11_inst : DFF_X1 port map( D => n10064, CK => CLK, Q => n52796,
                           QN => n1303);
   REGS_reg_133_10_inst : DFF_X1 port map( D => n10063, CK => CLK, Q => n52797,
                           QN => n1304);
   REGS_reg_133_9_inst : DFF_X1 port map( D => n10062, CK => CLK, Q => n52798, 
                           QN => n1305);
   REGS_reg_133_8_inst : DFF_X1 port map( D => n10061, CK => CLK, Q => n52799, 
                           QN => n1306);
   REGS_reg_133_7_inst : DFF_X1 port map( D => n10060, CK => CLK, Q => n52800, 
                           QN => n1307);
   REGS_reg_133_6_inst : DFF_X1 port map( D => n10059, CK => CLK, Q => n52801, 
                           QN => n1308);
   REGS_reg_133_5_inst : DFF_X1 port map( D => n10058, CK => CLK, Q => n52802, 
                           QN => n1309);
   REGS_reg_133_4_inst : DFF_X1 port map( D => n10057, CK => CLK, Q => n52803, 
                           QN => n1310);
   REGS_reg_133_3_inst : DFF_X1 port map( D => n10056, CK => CLK, Q => n52804, 
                           QN => n1311);
   REGS_reg_133_2_inst : DFF_X1 port map( D => n10055, CK => CLK, Q => n52805, 
                           QN => n1312);
   REGS_reg_133_1_inst : DFF_X1 port map( D => n10054, CK => CLK, Q => n52806, 
                           QN => n1313);
   REGS_reg_133_0_inst : DFF_X1 port map( D => n10053, CK => CLK, Q => n52807, 
                           QN => n1314);
   REGS_reg_132_23_inst : DFF_X1 port map( D => n10108, CK => CLK, Q => n_1418,
                           QN => n1315);
   REGS_reg_132_22_inst : DFF_X1 port map( D => n10107, CK => CLK, Q => n_1419,
                           QN => n1316);
   REGS_reg_132_21_inst : DFF_X1 port map( D => n10106, CK => CLK, Q => n_1420,
                           QN => n1317);
   REGS_reg_132_20_inst : DFF_X1 port map( D => n10105, CK => CLK, Q => n_1421,
                           QN => n1318);
   REGS_reg_132_19_inst : DFF_X1 port map( D => n10104, CK => CLK, Q => n_1422,
                           QN => n1319);
   REGS_reg_132_18_inst : DFF_X1 port map( D => n10103, CK => CLK, Q => n_1423,
                           QN => n1320);
   REGS_reg_132_17_inst : DFF_X1 port map( D => n10102, CK => CLK, Q => n_1424,
                           QN => n1321);
   REGS_reg_132_16_inst : DFF_X1 port map( D => n10101, CK => CLK, Q => n_1425,
                           QN => n1322);
   REGS_reg_132_15_inst : DFF_X1 port map( D => n10100, CK => CLK, Q => n_1426,
                           QN => n1323);
   REGS_reg_132_14_inst : DFF_X1 port map( D => n10099, CK => CLK, Q => n_1427,
                           QN => n1324);
   REGS_reg_132_13_inst : DFF_X1 port map( D => n10098, CK => CLK, Q => n_1428,
                           QN => n1325);
   REGS_reg_132_12_inst : DFF_X1 port map( D => n10097, CK => CLK, Q => n_1429,
                           QN => n1326);
   REGS_reg_132_11_inst : DFF_X1 port map( D => n10096, CK => CLK, Q => n_1430,
                           QN => n1327);
   REGS_reg_131_10_inst : DFF_X1 port map( D => n10127, CK => CLK, Q => n_1431,
                           QN => n1328);
   REGS_reg_131_9_inst : DFF_X1 port map( D => n10126, CK => CLK, Q => n_1432, 
                           QN => n1329);
   REGS_reg_131_8_inst : DFF_X1 port map( D => n10125, CK => CLK, Q => n_1433, 
                           QN => n1330);
   REGS_reg_131_7_inst : DFF_X1 port map( D => n10124, CK => CLK, Q => n_1434, 
                           QN => n1331);
   REGS_reg_131_6_inst : DFF_X1 port map( D => n10123, CK => CLK, Q => n_1435, 
                           QN => n1332);
   REGS_reg_131_5_inst : DFF_X1 port map( D => n10122, CK => CLK, Q => n_1436, 
                           QN => n1333);
   REGS_reg_131_4_inst : DFF_X1 port map( D => n10121, CK => CLK, Q => n_1437, 
                           QN => n1334);
   REGS_reg_131_3_inst : DFF_X1 port map( D => n10120, CK => CLK, Q => n_1438, 
                           QN => n1335);
   REGS_reg_131_2_inst : DFF_X1 port map( D => n10119, CK => CLK, Q => n_1439, 
                           QN => n1336);
   REGS_reg_131_1_inst : DFF_X1 port map( D => n10118, CK => CLK, Q => n_1440, 
                           QN => n1337);
   REGS_reg_131_0_inst : DFF_X1 port map( D => n10117, CK => CLK, Q => n_1441, 
                           QN => n1338);
   REGS_reg_132_10_inst : DFF_X1 port map( D => n10095, CK => CLK, Q => n_1442,
                           QN => n1339);
   REGS_reg_132_9_inst : DFF_X1 port map( D => n10094, CK => CLK, Q => n_1443, 
                           QN => n1340);
   REGS_reg_132_8_inst : DFF_X1 port map( D => n10093, CK => CLK, Q => n_1444, 
                           QN => n1341);
   REGS_reg_132_7_inst : DFF_X1 port map( D => n10092, CK => CLK, Q => n_1445, 
                           QN => n1342);
   REGS_reg_132_6_inst : DFF_X1 port map( D => n10091, CK => CLK, Q => n_1446, 
                           QN => n1343);
   REGS_reg_132_5_inst : DFF_X1 port map( D => n10090, CK => CLK, Q => n_1447, 
                           QN => n1344);
   REGS_reg_132_4_inst : DFF_X1 port map( D => n10089, CK => CLK, Q => n_1448, 
                           QN => n1345);
   REGS_reg_132_3_inst : DFF_X1 port map( D => n10088, CK => CLK, Q => n_1449, 
                           QN => n1346);
   REGS_reg_132_2_inst : DFF_X1 port map( D => n10087, CK => CLK, Q => n_1450, 
                           QN => n1347);
   REGS_reg_132_1_inst : DFF_X1 port map( D => n10086, CK => CLK, Q => n_1451, 
                           QN => n1348);
   REGS_reg_132_0_inst : DFF_X1 port map( D => n10085, CK => CLK, Q => n_1452, 
                           QN => n1349);
   REGS_reg_131_23_inst : DFF_X1 port map( D => n10140, CK => CLK, Q => n_1453,
                           QN => n1350);
   REGS_reg_131_22_inst : DFF_X1 port map( D => n10139, CK => CLK, Q => n_1454,
                           QN => n1351);
   REGS_reg_131_21_inst : DFF_X1 port map( D => n10138, CK => CLK, Q => n_1455,
                           QN => n1352);
   REGS_reg_131_20_inst : DFF_X1 port map( D => n10137, CK => CLK, Q => n_1456,
                           QN => n1353);
   REGS_reg_131_19_inst : DFF_X1 port map( D => n10136, CK => CLK, Q => n_1457,
                           QN => n1354);
   REGS_reg_131_18_inst : DFF_X1 port map( D => n10135, CK => CLK, Q => n_1458,
                           QN => n1355);
   REGS_reg_131_17_inst : DFF_X1 port map( D => n10134, CK => CLK, Q => n_1459,
                           QN => n1356);
   REGS_reg_131_16_inst : DFF_X1 port map( D => n10133, CK => CLK, Q => n_1460,
                           QN => n1357);
   REGS_reg_131_15_inst : DFF_X1 port map( D => n10132, CK => CLK, Q => n_1461,
                           QN => n1358);
   REGS_reg_131_14_inst : DFF_X1 port map( D => n10131, CK => CLK, Q => n_1462,
                           QN => n1359);
   REGS_reg_131_13_inst : DFF_X1 port map( D => n10130, CK => CLK, Q => n_1463,
                           QN => n1360);
   REGS_reg_131_12_inst : DFF_X1 port map( D => n10129, CK => CLK, Q => n_1464,
                           QN => n1361);
   REGS_reg_131_11_inst : DFF_X1 port map( D => n10128, CK => CLK, Q => n_1465,
                           QN => n1362);
   REGS_reg_130_23_inst : DFF_X1 port map( D => n10172, CK => CLK, Q => n_1466,
                           QN => n1363);
   REGS_reg_130_22_inst : DFF_X1 port map( D => n10171, CK => CLK, Q => n_1467,
                           QN => n1364);
   REGS_reg_130_21_inst : DFF_X1 port map( D => n10170, CK => CLK, Q => n_1468,
                           QN => n1365);
   REGS_reg_130_20_inst : DFF_X1 port map( D => n10169, CK => CLK, Q => n_1469,
                           QN => n1366);
   REGS_reg_130_19_inst : DFF_X1 port map( D => n10168, CK => CLK, Q => n_1470,
                           QN => n1367);
   REGS_reg_130_18_inst : DFF_X1 port map( D => n10167, CK => CLK, Q => n_1471,
                           QN => n1368);
   REGS_reg_130_17_inst : DFF_X1 port map( D => n10166, CK => CLK, Q => n_1472,
                           QN => n1369);
   REGS_reg_130_16_inst : DFF_X1 port map( D => n10165, CK => CLK, Q => n_1473,
                           QN => n1370);
   REGS_reg_130_15_inst : DFF_X1 port map( D => n10164, CK => CLK, Q => n_1474,
                           QN => n1371);
   REGS_reg_130_14_inst : DFF_X1 port map( D => n10163, CK => CLK, Q => n_1475,
                           QN => n1372);
   REGS_reg_130_13_inst : DFF_X1 port map( D => n10162, CK => CLK, Q => n_1476,
                           QN => n1373);
   REGS_reg_130_12_inst : DFF_X1 port map( D => n10161, CK => CLK, Q => n_1477,
                           QN => n1374);
   REGS_reg_130_11_inst : DFF_X1 port map( D => n10160, CK => CLK, Q => n_1478,
                           QN => n1375);
   REGS_reg_130_10_inst : DFF_X1 port map( D => n10159, CK => CLK, Q => n_1479,
                           QN => n1376);
   REGS_reg_130_9_inst : DFF_X1 port map( D => n10158, CK => CLK, Q => n_1480, 
                           QN => n1377);
   REGS_reg_130_8_inst : DFF_X1 port map( D => n10157, CK => CLK, Q => n_1481, 
                           QN => n1378);
   REGS_reg_130_7_inst : DFF_X1 port map( D => n10156, CK => CLK, Q => n_1482, 
                           QN => n1379);
   REGS_reg_130_6_inst : DFF_X1 port map( D => n10155, CK => CLK, Q => n_1483, 
                           QN => n1380);
   REGS_reg_130_5_inst : DFF_X1 port map( D => n10154, CK => CLK, Q => n_1484, 
                           QN => n1381);
   REGS_reg_130_4_inst : DFF_X1 port map( D => n10153, CK => CLK, Q => n_1485, 
                           QN => n1382);
   REGS_reg_130_3_inst : DFF_X1 port map( D => n10152, CK => CLK, Q => n_1486, 
                           QN => n1383);
   REGS_reg_130_2_inst : DFF_X1 port map( D => n10151, CK => CLK, Q => n_1487, 
                           QN => n1384);
   REGS_reg_130_1_inst : DFF_X1 port map( D => n10150, CK => CLK, Q => n_1488, 
                           QN => n1385);
   REGS_reg_130_0_inst : DFF_X1 port map( D => n10149, CK => CLK, Q => n_1489, 
                           QN => n1386);
   REGS_reg_129_23_inst : DFF_X1 port map( D => n10204, CK => CLK, Q => n_1490,
                           QN => n1387);
   REGS_reg_129_22_inst : DFF_X1 port map( D => n10203, CK => CLK, Q => n_1491,
                           QN => n1388);
   REGS_reg_129_21_inst : DFF_X1 port map( D => n10202, CK => CLK, Q => n_1492,
                           QN => n1389);
   REGS_reg_129_20_inst : DFF_X1 port map( D => n10201, CK => CLK, Q => n_1493,
                           QN => n1390);
   REGS_reg_129_19_inst : DFF_X1 port map( D => n10200, CK => CLK, Q => n_1494,
                           QN => n1391);
   REGS_reg_129_18_inst : DFF_X1 port map( D => n10199, CK => CLK, Q => n_1495,
                           QN => n1392);
   REGS_reg_129_17_inst : DFF_X1 port map( D => n10198, CK => CLK, Q => n_1496,
                           QN => n1393);
   REGS_reg_129_16_inst : DFF_X1 port map( D => n10197, CK => CLK, Q => n_1497,
                           QN => n1394);
   REGS_reg_129_15_inst : DFF_X1 port map( D => n10196, CK => CLK, Q => n_1498,
                           QN => n1395);
   REGS_reg_129_14_inst : DFF_X1 port map( D => n10195, CK => CLK, Q => n_1499,
                           QN => n1396);
   REGS_reg_129_13_inst : DFF_X1 port map( D => n10194, CK => CLK, Q => n_1500,
                           QN => n1397);
   REGS_reg_129_12_inst : DFF_X1 port map( D => n10193, CK => CLK, Q => n_1501,
                           QN => n1398);
   REGS_reg_129_11_inst : DFF_X1 port map( D => n10192, CK => CLK, Q => n_1502,
                           QN => n1399);
   REGS_reg_129_10_inst : DFF_X1 port map( D => n10191, CK => CLK, Q => n_1503,
                           QN => n1400);
   REGS_reg_129_9_inst : DFF_X1 port map( D => n10190, CK => CLK, Q => n_1504, 
                           QN => n1401);
   REGS_reg_129_8_inst : DFF_X1 port map( D => n10189, CK => CLK, Q => n_1505, 
                           QN => n1402);
   REGS_reg_129_7_inst : DFF_X1 port map( D => n10188, CK => CLK, Q => n_1506, 
                           QN => n1403);
   REGS_reg_129_6_inst : DFF_X1 port map( D => n10187, CK => CLK, Q => n_1507, 
                           QN => n1404);
   REGS_reg_129_5_inst : DFF_X1 port map( D => n10186, CK => CLK, Q => n_1508, 
                           QN => n1405);
   REGS_reg_129_4_inst : DFF_X1 port map( D => n10185, CK => CLK, Q => n_1509, 
                           QN => n1406);
   REGS_reg_129_3_inst : DFF_X1 port map( D => n10184, CK => CLK, Q => n_1510, 
                           QN => n1407);
   REGS_reg_129_2_inst : DFF_X1 port map( D => n10183, CK => CLK, Q => n_1511, 
                           QN => n1408);
   REGS_reg_129_1_inst : DFF_X1 port map( D => n10182, CK => CLK, Q => n_1512, 
                           QN => n1409);
   REGS_reg_129_0_inst : DFF_X1 port map( D => n10181, CK => CLK, Q => n_1513, 
                           QN => n1410);
   REGS_reg_128_23_inst : DFF_X1 port map( D => n10236, CK => CLK, Q => n15519,
                           QN => n1411);
   REGS_reg_128_22_inst : DFF_X1 port map( D => n10235, CK => CLK, Q => n15518,
                           QN => n1412);
   REGS_reg_128_21_inst : DFF_X1 port map( D => n10234, CK => CLK, Q => n15517,
                           QN => n1413);
   REGS_reg_128_20_inst : DFF_X1 port map( D => n10233, CK => CLK, Q => n15516,
                           QN => n1414);
   REGS_reg_128_19_inst : DFF_X1 port map( D => n10232, CK => CLK, Q => n15515,
                           QN => n1415);
   REGS_reg_128_18_inst : DFF_X1 port map( D => n10231, CK => CLK, Q => n15514,
                           QN => n1416);
   REGS_reg_128_17_inst : DFF_X1 port map( D => n10230, CK => CLK, Q => n15513,
                           QN => n1417);
   REGS_reg_128_16_inst : DFF_X1 port map( D => n10229, CK => CLK, Q => n15512,
                           QN => n1418);
   REGS_reg_128_15_inst : DFF_X1 port map( D => n10228, CK => CLK, Q => n15511,
                           QN => n1419);
   REGS_reg_128_14_inst : DFF_X1 port map( D => n10227, CK => CLK, Q => n15510,
                           QN => n1420);
   REGS_reg_128_13_inst : DFF_X1 port map( D => n10226, CK => CLK, Q => n15509,
                           QN => n1421);
   REGS_reg_128_12_inst : DFF_X1 port map( D => n10225, CK => CLK, Q => n15508,
                           QN => n1422);
   REGS_reg_128_11_inst : DFF_X1 port map( D => n10224, CK => CLK, Q => n15507,
                           QN => n1423);
   REGS_reg_128_10_inst : DFF_X1 port map( D => n10223, CK => CLK, Q => n15506,
                           QN => n1424);
   REGS_reg_128_9_inst : DFF_X1 port map( D => n10222, CK => CLK, Q => n15505, 
                           QN => n1425);
   REGS_reg_128_8_inst : DFF_X1 port map( D => n10221, CK => CLK, Q => n15504, 
                           QN => n1426);
   REGS_reg_128_7_inst : DFF_X1 port map( D => n10220, CK => CLK, Q => n15503, 
                           QN => n1427);
   REGS_reg_128_6_inst : DFF_X1 port map( D => n10219, CK => CLK, Q => n15502, 
                           QN => n1428);
   REGS_reg_128_5_inst : DFF_X1 port map( D => n10218, CK => CLK, Q => n15501, 
                           QN => n1429);
   REGS_reg_128_4_inst : DFF_X1 port map( D => n10217, CK => CLK, Q => n15500, 
                           QN => n1430);
   REGS_reg_128_3_inst : DFF_X1 port map( D => n10216, CK => CLK, Q => n15499, 
                           QN => n1431);
   REGS_reg_128_2_inst : DFF_X1 port map( D => n10215, CK => CLK, Q => n15466, 
                           QN => n1432);
   REGS_reg_128_1_inst : DFF_X1 port map( D => n10214, CK => CLK, Q => n15465, 
                           QN => n1433);
   REGS_reg_128_0_inst : DFF_X1 port map( D => n10213, CK => CLK, Q => n15464, 
                           QN => n1434);
   REGS_reg_31_23_inst : DFF_X1 port map( D => n13340, CK => CLK, Q => n52856, 
                           QN => n1435);
   REGS_reg_31_22_inst : DFF_X1 port map( D => n13339, CK => CLK, Q => n52857, 
                           QN => n1436);
   REGS_reg_31_21_inst : DFF_X1 port map( D => n13338, CK => CLK, Q => n52858, 
                           QN => n1437);
   REGS_reg_31_20_inst : DFF_X1 port map( D => n13337, CK => CLK, Q => n52859, 
                           QN => n1438);
   REGS_reg_31_19_inst : DFF_X1 port map( D => n13336, CK => CLK, Q => n52860, 
                           QN => n1439);
   REGS_reg_31_18_inst : DFF_X1 port map( D => n13335, CK => CLK, Q => n52861, 
                           QN => n1440);
   REGS_reg_31_17_inst : DFF_X1 port map( D => n13334, CK => CLK, Q => n52862, 
                           QN => n1441);
   REGS_reg_31_16_inst : DFF_X1 port map( D => n13333, CK => CLK, Q => n52863, 
                           QN => n1442);
   REGS_reg_31_15_inst : DFF_X1 port map( D => n13332, CK => CLK, Q => n52864, 
                           QN => n1443);
   REGS_reg_31_14_inst : DFF_X1 port map( D => n13331, CK => CLK, Q => n52865, 
                           QN => n1444);
   REGS_reg_31_13_inst : DFF_X1 port map( D => n13330, CK => CLK, Q => n52866, 
                           QN => n1445);
   REGS_reg_31_12_inst : DFF_X1 port map( D => n13329, CK => CLK, Q => n52867, 
                           QN => n1446);
   REGS_reg_31_11_inst : DFF_X1 port map( D => n13328, CK => CLK, Q => n52868, 
                           QN => n1447);
   REGS_reg_31_10_inst : DFF_X1 port map( D => n13327, CK => CLK, Q => n52869, 
                           QN => n1448);
   REGS_reg_31_9_inst : DFF_X1 port map( D => n13326, CK => CLK, Q => n52870, 
                           QN => n1449);
   REGS_reg_31_8_inst : DFF_X1 port map( D => n13325, CK => CLK, Q => n52871, 
                           QN => n1450);
   REGS_reg_31_7_inst : DFF_X1 port map( D => n13324, CK => CLK, Q => n52872, 
                           QN => n1451);
   REGS_reg_31_6_inst : DFF_X1 port map( D => n13323, CK => CLK, Q => n52873, 
                           QN => n1452);
   REGS_reg_31_5_inst : DFF_X1 port map( D => n13322, CK => CLK, Q => n52874, 
                           QN => n1453);
   REGS_reg_31_4_inst : DFF_X1 port map( D => n13321, CK => CLK, Q => n52875, 
                           QN => n1454);
   REGS_reg_31_3_inst : DFF_X1 port map( D => n13320, CK => CLK, Q => n52876, 
                           QN => n1455);
   REGS_reg_31_2_inst : DFF_X1 port map( D => n13319, CK => CLK, Q => n52877, 
                           QN => n1456);
   REGS_reg_31_1_inst : DFF_X1 port map( D => n13318, CK => CLK, Q => n52878, 
                           QN => n1457);
   REGS_reg_31_0_inst : DFF_X1 port map( D => n13317, CK => CLK, Q => n52879, 
                           QN => n1458);
   REGS_reg_30_23_inst : DFF_X1 port map( D => n13372, CK => CLK, Q => n15850, 
                           QN => n1459);
   REGS_reg_30_22_inst : DFF_X1 port map( D => n13371, CK => CLK, Q => n15849, 
                           QN => n1460);
   REGS_reg_30_21_inst : DFF_X1 port map( D => n13370, CK => CLK, Q => n15848, 
                           QN => n1461);
   REGS_reg_30_20_inst : DFF_X1 port map( D => n13369, CK => CLK, Q => n15847, 
                           QN => n1462);
   REGS_reg_30_19_inst : DFF_X1 port map( D => n13368, CK => CLK, Q => n15846, 
                           QN => n1463);
   REGS_reg_30_18_inst : DFF_X1 port map( D => n13367, CK => CLK, Q => n15845, 
                           QN => n1464);
   REGS_reg_30_17_inst : DFF_X1 port map( D => n13366, CK => CLK, Q => n15844, 
                           QN => n1465);
   REGS_reg_30_16_inst : DFF_X1 port map( D => n13365, CK => CLK, Q => n15843, 
                           QN => n1466);
   REGS_reg_30_15_inst : DFF_X1 port map( D => n13364, CK => CLK, Q => n15842, 
                           QN => n1467);
   REGS_reg_30_14_inst : DFF_X1 port map( D => n13363, CK => CLK, Q => n15841, 
                           QN => n1468);
   REGS_reg_30_13_inst : DFF_X1 port map( D => n13362, CK => CLK, Q => n15840, 
                           QN => n1469);
   REGS_reg_30_12_inst : DFF_X1 port map( D => n13361, CK => CLK, Q => n15839, 
                           QN => n1470);
   REGS_reg_30_11_inst : DFF_X1 port map( D => n13360, CK => CLK, Q => n15838, 
                           QN => n1471);
   REGS_reg_30_10_inst : DFF_X1 port map( D => n13359, CK => CLK, Q => n15837, 
                           QN => n1472);
   REGS_reg_30_9_inst : DFF_X1 port map( D => n13358, CK => CLK, Q => n15836, 
                           QN => n1473);
   REGS_reg_30_8_inst : DFF_X1 port map( D => n13357, CK => CLK, Q => n15835, 
                           QN => n1474);
   REGS_reg_30_7_inst : DFF_X1 port map( D => n13356, CK => CLK, Q => n15834, 
                           QN => n1475);
   REGS_reg_30_6_inst : DFF_X1 port map( D => n13355, CK => CLK, Q => n15833, 
                           QN => n1476);
   REGS_reg_30_5_inst : DFF_X1 port map( D => n13354, CK => CLK, Q => n15832, 
                           QN => n1477);
   REGS_reg_30_4_inst : DFF_X1 port map( D => n13353, CK => CLK, Q => n15831, 
                           QN => n1478);
   REGS_reg_30_3_inst : DFF_X1 port map( D => n13352, CK => CLK, Q => n15830, 
                           QN => n1479);
   REGS_reg_30_2_inst : DFF_X1 port map( D => n13351, CK => CLK, Q => n15829, 
                           QN => n1480);
   REGS_reg_30_1_inst : DFF_X1 port map( D => n13350, CK => CLK, Q => n15828, 
                           QN => n1481);
   REGS_reg_30_0_inst : DFF_X1 port map( D => n13349, CK => CLK, Q => n15827, 
                           QN => n1482);
   REGS_reg_29_23_inst : DFF_X1 port map( D => n13404, CK => CLK, Q => n15826, 
                           QN => n1483);
   REGS_reg_29_22_inst : DFF_X1 port map( D => n13403, CK => CLK, Q => n15825, 
                           QN => n1484);
   REGS_reg_29_21_inst : DFF_X1 port map( D => n13402, CK => CLK, Q => n15824, 
                           QN => n1485);
   REGS_reg_29_20_inst : DFF_X1 port map( D => n13401, CK => CLK, Q => n15823, 
                           QN => n1486);
   REGS_reg_29_19_inst : DFF_X1 port map( D => n13400, CK => CLK, Q => n15822, 
                           QN => n1487);
   REGS_reg_29_18_inst : DFF_X1 port map( D => n13399, CK => CLK, Q => n15821, 
                           QN => n1488);
   REGS_reg_29_17_inst : DFF_X1 port map( D => n13398, CK => CLK, Q => n15820, 
                           QN => n1489);
   REGS_reg_29_16_inst : DFF_X1 port map( D => n13397, CK => CLK, Q => n15819, 
                           QN => n1490);
   REGS_reg_29_15_inst : DFF_X1 port map( D => n13396, CK => CLK, Q => n15818, 
                           QN => n1491);
   REGS_reg_29_14_inst : DFF_X1 port map( D => n13395, CK => CLK, Q => n15817, 
                           QN => n1492);
   REGS_reg_29_13_inst : DFF_X1 port map( D => n13394, CK => CLK, Q => n15816, 
                           QN => n1493);
   REGS_reg_29_12_inst : DFF_X1 port map( D => n13393, CK => CLK, Q => n15815, 
                           QN => n1494);
   REGS_reg_29_11_inst : DFF_X1 port map( D => n13392, CK => CLK, Q => n15814, 
                           QN => n1495);
   REGS_reg_29_10_inst : DFF_X1 port map( D => n13391, CK => CLK, Q => n15813, 
                           QN => n1496);
   REGS_reg_29_9_inst : DFF_X1 port map( D => n13390, CK => CLK, Q => n15812, 
                           QN => n1497);
   REGS_reg_29_8_inst : DFF_X1 port map( D => n13389, CK => CLK, Q => n15811, 
                           QN => n1498);
   REGS_reg_29_7_inst : DFF_X1 port map( D => n13388, CK => CLK, Q => n15810, 
                           QN => n1499);
   REGS_reg_29_6_inst : DFF_X1 port map( D => n13387, CK => CLK, Q => n15809, 
                           QN => n1500);
   REGS_reg_29_5_inst : DFF_X1 port map( D => n13386, CK => CLK, Q => n15808, 
                           QN => n1501);
   REGS_reg_29_4_inst : DFF_X1 port map( D => n13385, CK => CLK, Q => n15807, 
                           QN => n1502);
   REGS_reg_29_3_inst : DFF_X1 port map( D => n13384, CK => CLK, Q => n15806, 
                           QN => n1503);
   REGS_reg_29_2_inst : DFF_X1 port map( D => n13383, CK => CLK, Q => n15805, 
                           QN => n1504);
   REGS_reg_29_1_inst : DFF_X1 port map( D => n13382, CK => CLK, Q => n15804, 
                           QN => n1505);
   REGS_reg_29_0_inst : DFF_X1 port map( D => n13381, CK => CLK, Q => n15803, 
                           QN => n1506);
   REGS_reg_27_4_inst : DFF_X1 port map( D => n13449, CK => CLK, Q => n519, QN 
                           => n1507);
   REGS_reg_26_23_inst : DFF_X1 port map( D => n13500, CK => CLK, Q => n16208, 
                           QN => n1508);
   REGS_reg_26_22_inst : DFF_X1 port map( D => n13499, CK => CLK, Q => n16202, 
                           QN => n1509);
   REGS_reg_26_21_inst : DFF_X1 port map( D => n13498, CK => CLK, Q => n16196, 
                           QN => n1510);
   REGS_reg_26_20_inst : DFF_X1 port map( D => n13497, CK => CLK, Q => n16190, 
                           QN => n1511);
   REGS_reg_26_19_inst : DFF_X1 port map( D => n13496, CK => CLK, Q => n16256, 
                           QN => n1512);
   REGS_reg_26_18_inst : DFF_X1 port map( D => n13495, CK => CLK, Q => n16250, 
                           QN => n1513);
   REGS_reg_26_17_inst : DFF_X1 port map( D => n13494, CK => CLK, Q => n16244, 
                           QN => n1514);
   REGS_reg_26_16_inst : DFF_X1 port map( D => n13493, CK => CLK, Q => n16238, 
                           QN => n1515);
   REGS_reg_26_15_inst : DFF_X1 port map( D => n13492, CK => CLK, Q => n16232, 
                           QN => n1516);
   REGS_reg_26_14_inst : DFF_X1 port map( D => n13491, CK => CLK, Q => n16280, 
                           QN => n1517);
   REGS_reg_26_13_inst : DFF_X1 port map( D => n13490, CK => CLK, Q => n_1514, 
                           QN => n1520);
   REGS_reg_26_12_inst : DFF_X1 port map( D => n13489, CK => CLK, Q => n_1515, 
                           QN => n1522);
   REGS_reg_26_11_inst : DFF_X1 port map( D => n13488, CK => CLK, Q => n_1516, 
                           QN => n1524);
   REGS_reg_26_10_inst : DFF_X1 port map( D => n13487, CK => CLK, Q => n_1517, 
                           QN => n1526);
   REGS_reg_26_9_inst : DFF_X1 port map( D => n13486, CK => CLK, Q => n_1518, 
                           QN => n1528);
   REGS_reg_26_8_inst : DFF_X1 port map( D => n13485, CK => CLK, Q => n_1519, 
                           QN => n1530);
   REGS_reg_26_7_inst : DFF_X1 port map( D => n13484, CK => CLK, Q => n_1520, 
                           QN => n1532);
   REGS_reg_26_6_inst : DFF_X1 port map( D => n13483, CK => CLK, Q => n_1521, 
                           QN => n1534);
   REGS_reg_26_5_inst : DFF_X1 port map( D => n13482, CK => CLK, Q => n_1522, 
                           QN => n1536);
   REGS_reg_26_4_inst : DFF_X1 port map( D => n13481, CK => CLK, Q => n_1523, 
                           QN => n1538);
   REGS_reg_26_3_inst : DFF_X1 port map( D => n13480, CK => CLK, Q => n_1524, 
                           QN => n1540);
   REGS_reg_26_2_inst : DFF_X1 port map( D => n13479, CK => CLK, Q => n_1525, 
                           QN => n1542);
   REGS_reg_26_1_inst : DFF_X1 port map( D => n13478, CK => CLK, Q => n_1526, 
                           QN => n1544);
   REGS_reg_26_0_inst : DFF_X1 port map( D => n13477, CK => CLK, Q => n_1527, 
                           QN => n1546);
   REGS_reg_25_23_inst : DFF_X1 port map( D => n13532, CK => CLK, Q => n16207, 
                           QN => n1547);
   REGS_reg_25_22_inst : DFF_X1 port map( D => n13531, CK => CLK, Q => n16201, 
                           QN => n1548);
   REGS_reg_25_21_inst : DFF_X1 port map( D => n13530, CK => CLK, Q => n16195, 
                           QN => n1549);
   REGS_reg_25_20_inst : DFF_X1 port map( D => n13529, CK => CLK, Q => n16189, 
                           QN => n1550);
   REGS_reg_25_19_inst : DFF_X1 port map( D => n13528, CK => CLK, Q => n16255, 
                           QN => n1551);
   REGS_reg_25_18_inst : DFF_X1 port map( D => n13527, CK => CLK, Q => n16249, 
                           QN => n1552);
   REGS_reg_25_17_inst : DFF_X1 port map( D => n13526, CK => CLK, Q => n16243, 
                           QN => n1553);
   REGS_reg_25_16_inst : DFF_X1 port map( D => n13525, CK => CLK, Q => n16237, 
                           QN => n1554);
   REGS_reg_25_15_inst : DFF_X1 port map( D => n13524, CK => CLK, Q => n16231, 
                           QN => n1555);
   REGS_reg_25_14_inst : DFF_X1 port map( D => n13523, CK => CLK, Q => n16279, 
                           QN => n1556);
   REGS_reg_25_13_inst : DFF_X1 port map( D => n13522, CK => CLK, Q => n_1528, 
                           QN => n1557);
   REGS_reg_25_12_inst : DFF_X1 port map( D => n13521, CK => CLK, Q => n_1529, 
                           QN => n1558);
   REGS_reg_25_11_inst : DFF_X1 port map( D => n13520, CK => CLK, Q => n_1530, 
                           QN => n1589);
   REGS_reg_25_10_inst : DFF_X1 port map( D => n13519, CK => CLK, Q => n_1531, 
                           QN => n1590);
   REGS_reg_25_9_inst : DFF_X1 port map( D => n13518, CK => CLK, Q => n_1532, 
                           QN => n1607);
   REGS_reg_25_8_inst : DFF_X1 port map( D => n13517, CK => CLK, Q => n_1533, 
                           QN => n1608);
   REGS_reg_25_7_inst : DFF_X1 port map( D => n13516, CK => CLK, Q => n_1534, 
                           QN => n1609);
   REGS_reg_25_6_inst : DFF_X1 port map( D => n13515, CK => CLK, Q => n_1535, 
                           QN => n1610);
   REGS_reg_25_5_inst : DFF_X1 port map( D => n13514, CK => CLK, Q => n_1536, 
                           QN => n1611);
   REGS_reg_25_4_inst : DFF_X1 port map( D => n13513, CK => CLK, Q => n_1537, 
                           QN => n1612);
   REGS_reg_25_3_inst : DFF_X1 port map( D => n13512, CK => CLK, Q => n_1538, 
                           QN => n1613);
   REGS_reg_25_2_inst : DFF_X1 port map( D => n13511, CK => CLK, Q => n_1539, 
                           QN => n1614);
   REGS_reg_25_1_inst : DFF_X1 port map( D => n13510, CK => CLK, Q => n_1540, 
                           QN => n1615);
   REGS_reg_25_0_inst : DFF_X1 port map( D => n13509, CK => CLK, Q => n_1541, 
                           QN => n1616);
   REGS_reg_24_23_inst : DFF_X1 port map( D => n13564, CK => CLK, Q => n15874, 
                           QN => n1617);
   REGS_reg_24_22_inst : DFF_X1 port map( D => n13563, CK => CLK, Q => n15869, 
                           QN => n1618);
   REGS_reg_24_21_inst : DFF_X1 port map( D => n13562, CK => CLK, Q => n15864, 
                           QN => n1619);
   REGS_reg_24_20_inst : DFF_X1 port map( D => n13561, CK => CLK, Q => n15859, 
                           QN => n1620);
   REGS_reg_24_19_inst : DFF_X1 port map( D => n13560, CK => CLK, Q => n15854, 
                           QN => n1621);
   REGS_reg_24_18_inst : DFF_X1 port map( D => n13559, CK => CLK, Q => n15801, 
                           QN => n1622);
   REGS_reg_24_17_inst : DFF_X1 port map( D => n13558, CK => CLK, Q => n15796, 
                           QN => n1623);
   REGS_reg_24_16_inst : DFF_X1 port map( D => n13557, CK => CLK, Q => n15791, 
                           QN => n1624);
   REGS_reg_24_15_inst : DFF_X1 port map( D => n13556, CK => CLK, Q => n15786, 
                           QN => n1625);
   REGS_reg_24_14_inst : DFF_X1 port map( D => n13555, CK => CLK, Q => n15781, 
                           QN => n1626);
   REGS_reg_24_13_inst : DFF_X1 port map( D => n13554, CK => CLK, Q => n15776, 
                           QN => n1627);
   REGS_reg_24_12_inst : DFF_X1 port map( D => n13553, CK => CLK, Q => n15771, 
                           QN => n1628);
   REGS_reg_24_11_inst : DFF_X1 port map( D => n13552, CK => CLK, Q => n15766, 
                           QN => n1629);
   REGS_reg_24_10_inst : DFF_X1 port map( D => n13551, CK => CLK, Q => n15761, 
                           QN => n1630);
   REGS_reg_24_9_inst : DFF_X1 port map( D => n13550, CK => CLK, Q => n15756, 
                           QN => n1647);
   REGS_reg_24_8_inst : DFF_X1 port map( D => n13549, CK => CLK, Q => n15751, 
                           QN => n1648);
   REGS_reg_24_7_inst : DFF_X1 port map( D => n13548, CK => CLK, Q => n15912, 
                           QN => n1649);
   REGS_reg_24_6_inst : DFF_X1 port map( D => n13547, CK => CLK, Q => n15907, 
                           QN => n1650);
   REGS_reg_24_5_inst : DFF_X1 port map( D => n13546, CK => CLK, Q => n15902, 
                           QN => n1651);
   REGS_reg_24_4_inst : DFF_X1 port map( D => n13545, CK => CLK, Q => n15897, 
                           QN => n1652);
   REGS_reg_24_3_inst : DFF_X1 port map( D => n13544, CK => CLK, Q => n15892, 
                           QN => n1653);
   REGS_reg_24_2_inst : DFF_X1 port map( D => n13543, CK => CLK, Q => n15914, 
                           QN => n1654);
   REGS_reg_24_1_inst : DFF_X1 port map( D => n13542, CK => CLK, Q => n15884, 
                           QN => n1655);
   REGS_reg_24_0_inst : DFF_X1 port map( D => n13541, CK => CLK, Q => n15879, 
                           QN => n1656);
   REGS_reg_23_23_inst : DFF_X1 port map( D => n13596, CK => CLK, Q => n15875, 
                           QN => n1657);
   REGS_reg_23_22_inst : DFF_X1 port map( D => n13595, CK => CLK, Q => n15870, 
                           QN => n1658);
   REGS_reg_23_21_inst : DFF_X1 port map( D => n13594, CK => CLK, Q => n15865, 
                           QN => n1659);
   REGS_reg_23_20_inst : DFF_X1 port map( D => n13593, CK => CLK, Q => n15860, 
                           QN => n1660);
   REGS_reg_23_19_inst : DFF_X1 port map( D => n13592, CK => CLK, Q => n15855, 
                           QN => n1661);
   REGS_reg_23_18_inst : DFF_X1 port map( D => n13591, CK => CLK, Q => n15802, 
                           QN => n1662);
   REGS_reg_23_17_inst : DFF_X1 port map( D => n13590, CK => CLK, Q => n15797, 
                           QN => n1663);
   REGS_reg_23_16_inst : DFF_X1 port map( D => n13589, CK => CLK, Q => n15792, 
                           QN => n1664);
   REGS_reg_23_15_inst : DFF_X1 port map( D => n13588, CK => CLK, Q => n15787, 
                           QN => n1665);
   REGS_reg_23_14_inst : DFF_X1 port map( D => n13587, CK => CLK, Q => n15782, 
                           QN => n1666);
   REGS_reg_23_13_inst : DFF_X1 port map( D => n13586, CK => CLK, Q => n15777, 
                           QN => n1667);
   REGS_reg_23_12_inst : DFF_X1 port map( D => n13585, CK => CLK, Q => n15772, 
                           QN => n1668);
   REGS_reg_23_11_inst : DFF_X1 port map( D => n13584, CK => CLK, Q => n15767, 
                           QN => n1693);
   REGS_reg_23_10_inst : DFF_X1 port map( D => n13583, CK => CLK, Q => n15762, 
                           QN => n1694);
   REGS_reg_23_9_inst : DFF_X1 port map( D => n13582, CK => CLK, Q => n15757, 
                           QN => n1695);
   REGS_reg_23_8_inst : DFF_X1 port map( D => n13581, CK => CLK, Q => n15752, 
                           QN => n1696);
   REGS_reg_23_7_inst : DFF_X1 port map( D => n13580, CK => CLK, Q => n15913, 
                           QN => n1697);
   REGS_reg_23_6_inst : DFF_X1 port map( D => n13579, CK => CLK, Q => n15908, 
                           QN => n1698);
   REGS_reg_23_5_inst : DFF_X1 port map( D => n13578, CK => CLK, Q => n15903, 
                           QN => n1699);
   REGS_reg_23_4_inst : DFF_X1 port map( D => n13577, CK => CLK, Q => n15898, 
                           QN => n1700);
   REGS_reg_23_3_inst : DFF_X1 port map( D => n13576, CK => CLK, Q => n15893, 
                           QN => n1701);
   REGS_reg_23_2_inst : DFF_X1 port map( D => n13575, CK => CLK, Q => n15915, 
                           QN => n1702);
   REGS_reg_23_1_inst : DFF_X1 port map( D => n13574, CK => CLK, Q => n15885, 
                           QN => n1703);
   REGS_reg_23_0_inst : DFF_X1 port map( D => n13573, CK => CLK, Q => n15880, 
                           QN => n1704);
   REGS_reg_22_23_inst : DFF_X1 port map( D => n13628, CK => CLK, Q => n_1542, 
                           QN => n1705);
   REGS_reg_22_22_inst : DFF_X1 port map( D => n13627, CK => CLK, Q => n_1543, 
                           QN => n1706);
   REGS_reg_22_21_inst : DFF_X1 port map( D => n13626, CK => CLK, Q => n_1544, 
                           QN => n1707);
   REGS_reg_22_20_inst : DFF_X1 port map( D => n13625, CK => CLK, Q => n_1545, 
                           QN => n1708);
   REGS_reg_22_19_inst : DFF_X1 port map( D => n13624, CK => CLK, Q => n_1546, 
                           QN => n1709);
   REGS_reg_22_18_inst : DFF_X1 port map( D => n13623, CK => CLK, Q => n_1547, 
                           QN => n1710);
   REGS_reg_22_17_inst : DFF_X1 port map( D => n13622, CK => CLK, Q => n_1548, 
                           QN => n1711);
   REGS_reg_22_16_inst : DFF_X1 port map( D => n13621, CK => CLK, Q => n_1549, 
                           QN => n1712);
   REGS_reg_22_15_inst : DFF_X1 port map( D => n13620, CK => CLK, Q => n_1550, 
                           QN => n1713);
   REGS_reg_22_14_inst : DFF_X1 port map( D => n13619, CK => CLK, Q => n_1551, 
                           QN => n1714);
   REGS_reg_22_13_inst : DFF_X1 port map( D => n13618, CK => CLK, Q => n_1552, 
                           QN => n1715);
   REGS_reg_22_12_inst : DFF_X1 port map( D => n13617, CK => CLK, Q => n_1553, 
                           QN => n1716);
   REGS_reg_22_11_inst : DFF_X1 port map( D => n13616, CK => CLK, Q => n_1554, 
                           QN => n1717);
   REGS_reg_22_10_inst : DFF_X1 port map( D => n13615, CK => CLK, Q => n_1555, 
                           QN => n1718);
   REGS_reg_22_9_inst : DFF_X1 port map( D => n13614, CK => CLK, Q => n_1556, 
                           QN => n1719);
   REGS_reg_22_8_inst : DFF_X1 port map( D => n13613, CK => CLK, Q => n_1557, 
                           QN => n1720);
   REGS_reg_22_7_inst : DFF_X1 port map( D => n13612, CK => CLK, Q => n_1558, 
                           QN => n1721);
   REGS_reg_22_6_inst : DFF_X1 port map( D => n13611, CK => CLK, Q => n_1559, 
                           QN => n1722);
   REGS_reg_22_5_inst : DFF_X1 port map( D => n13610, CK => CLK, Q => n_1560, 
                           QN => n1723);
   REGS_reg_22_4_inst : DFF_X1 port map( D => n13609, CK => CLK, Q => n_1561, 
                           QN => n1724);
   REGS_reg_22_3_inst : DFF_X1 port map( D => n13608, CK => CLK, Q => n_1562, 
                           QN => n1725);
   REGS_reg_22_2_inst : DFF_X1 port map( D => n13607, CK => CLK, Q => n_1563, 
                           QN => n1726);
   REGS_reg_22_1_inst : DFF_X1 port map( D => n13606, CK => CLK, Q => n_1564, 
                           QN => n1727);
   REGS_reg_22_0_inst : DFF_X1 port map( D => n13605, CK => CLK, Q => n_1565, 
                           QN => n1728);
   REGS_reg_21_23_inst : DFF_X1 port map( D => n13660, CK => CLK, Q => n15610, 
                           QN => n1729);
   REGS_reg_21_22_inst : DFF_X1 port map( D => n13659, CK => CLK, Q => n15609, 
                           QN => n1730);
   REGS_reg_21_21_inst : DFF_X1 port map( D => n13658, CK => CLK, Q => n15608, 
                           QN => n1731);
   REGS_reg_21_20_inst : DFF_X1 port map( D => n13657, CK => CLK, Q => n15607, 
                           QN => n1732);
   REGS_reg_21_19_inst : DFF_X1 port map( D => n13656, CK => CLK, Q => n15606, 
                           QN => n1733);
   REGS_reg_21_18_inst : DFF_X1 port map( D => n13655, CK => CLK, Q => n15605, 
                           QN => n1734);
   REGS_reg_21_17_inst : DFF_X1 port map( D => n13654, CK => CLK, Q => n15604, 
                           QN => n1735);
   REGS_reg_21_16_inst : DFF_X1 port map( D => n13653, CK => CLK, Q => n15603, 
                           QN => n1736);
   REGS_reg_21_15_inst : DFF_X1 port map( D => n13652, CK => CLK, Q => n15602, 
                           QN => n1737);
   REGS_reg_21_14_inst : DFF_X1 port map( D => n13651, CK => CLK, Q => n15601, 
                           QN => n1738);
   REGS_reg_62_23_inst : DFF_X1 port map( D => n12348, CK => CLK, Q => n592, QN
                           => n2779);
   REGS_reg_62_22_inst : DFF_X1 port map( D => n12347, CK => CLK, Q => n593, QN
                           => n2780);
   REGS_reg_62_21_inst : DFF_X1 port map( D => n12346, CK => CLK, Q => n594, QN
                           => n2781);
   REGS_reg_62_20_inst : DFF_X1 port map( D => n12345, CK => CLK, Q => n595, QN
                           => n2782);
   REGS_reg_62_19_inst : DFF_X1 port map( D => n12344, CK => CLK, Q => n596, QN
                           => n2783);
   REGS_reg_62_18_inst : DFF_X1 port map( D => n12343, CK => CLK, Q => n597, QN
                           => n2784);
   REGS_reg_62_17_inst : DFF_X1 port map( D => n12342, CK => CLK, Q => n598, QN
                           => n2785);
   REGS_reg_62_16_inst : DFF_X1 port map( D => n12341, CK => CLK, Q => n599, QN
                           => n2786);
   REGS_reg_62_15_inst : DFF_X1 port map( D => n12340, CK => CLK, Q => n600, QN
                           => n2787);
   REGS_reg_62_14_inst : DFF_X1 port map( D => n12339, CK => CLK, Q => n601, QN
                           => n2788);
   REGS_reg_62_13_inst : DFF_X1 port map( D => n12338, CK => CLK, Q => n602, QN
                           => n2789);
   REGS_reg_62_12_inst : DFF_X1 port map( D => n12337, CK => CLK, Q => n603, QN
                           => n2790);
   REGS_reg_62_11_inst : DFF_X1 port map( D => n12336, CK => CLK, Q => n604, QN
                           => n2839);
   REGS_reg_62_10_inst : DFF_X1 port map( D => n12335, CK => CLK, Q => n605, QN
                           => n2840);
   REGS_reg_62_9_inst : DFF_X1 port map( D => n12334, CK => CLK, Q => n606, QN 
                           => n2841);
   REGS_reg_62_8_inst : DFF_X1 port map( D => n12333, CK => CLK, Q => n607, QN 
                           => n2842);
   REGS_reg_62_7_inst : DFF_X1 port map( D => n12332, CK => CLK, Q => n608, QN 
                           => n2843);
   REGS_reg_62_6_inst : DFF_X1 port map( D => n12331, CK => CLK, Q => n609, QN 
                           => n2844);
   REGS_reg_62_5_inst : DFF_X1 port map( D => n12330, CK => CLK, Q => n610, QN 
                           => n2845);
   REGS_reg_62_4_inst : DFF_X1 port map( D => n12329, CK => CLK, Q => n611, QN 
                           => n2846);
   REGS_reg_62_3_inst : DFF_X1 port map( D => n12328, CK => CLK, Q => n612, QN 
                           => n2847);
   REGS_reg_62_2_inst : DFF_X1 port map( D => n12327, CK => CLK, Q => n613, QN 
                           => n2848);
   REGS_reg_62_1_inst : DFF_X1 port map( D => n12326, CK => CLK, Q => n614, QN 
                           => n2849);
   REGS_reg_62_0_inst : DFF_X1 port map( D => n12325, CK => CLK, Q => n615, QN 
                           => n2850);
   REGS_reg_61_23_inst : DFF_X1 port map( D => n12380, CK => CLK, Q => n616, QN
                           => n2851);
   REGS_reg_61_22_inst : DFF_X1 port map( D => n12379, CK => CLK, Q => n617, QN
                           => n2852);
   REGS_reg_61_21_inst : DFF_X1 port map( D => n12378, CK => CLK, Q => n618, QN
                           => n2853);
   REGS_reg_61_20_inst : DFF_X1 port map( D => n12377, CK => CLK, Q => n619, QN
                           => n2854);
   REGS_reg_61_19_inst : DFF_X1 port map( D => n12376, CK => CLK, Q => n620, QN
                           => n2855);
   REGS_reg_61_18_inst : DFF_X1 port map( D => n12375, CK => CLK, Q => n621, QN
                           => n2856);
   REGS_reg_61_17_inst : DFF_X1 port map( D => n12374, CK => CLK, Q => n622, QN
                           => n2857);
   REGS_reg_61_16_inst : DFF_X1 port map( D => n12373, CK => CLK, Q => n623, QN
                           => n2858);
   REGS_reg_61_15_inst : DFF_X1 port map( D => n12372, CK => CLK, Q => n624, QN
                           => n2859);
   REGS_reg_61_14_inst : DFF_X1 port map( D => n12371, CK => CLK, Q => n625, QN
                           => n2860);
   REGS_reg_61_13_inst : DFF_X1 port map( D => n12370, CK => CLK, Q => n626, QN
                           => n2861);
   REGS_reg_61_12_inst : DFF_X1 port map( D => n12369, CK => CLK, Q => n627, QN
                           => n2862);
   REGS_reg_61_11_inst : DFF_X1 port map( D => n12368, CK => CLK, Q => n628, QN
                           => n2863);
   REGS_reg_61_10_inst : DFF_X1 port map( D => n12367, CK => CLK, Q => n629, QN
                           => n2864);
   REGS_reg_61_9_inst : DFF_X1 port map( D => n12366, CK => CLK, Q => n630, QN 
                           => n2865);
   REGS_reg_61_8_inst : DFF_X1 port map( D => n12365, CK => CLK, Q => n631, QN 
                           => n2866);
   REGS_reg_61_7_inst : DFF_X1 port map( D => n12364, CK => CLK, Q => n632, QN 
                           => n2867);
   REGS_reg_61_6_inst : DFF_X1 port map( D => n12363, CK => CLK, Q => n633, QN 
                           => n2868);
   REGS_reg_61_5_inst : DFF_X1 port map( D => n12362, CK => CLK, Q => n634, QN 
                           => n2869);
   REGS_reg_61_4_inst : DFF_X1 port map( D => n12361, CK => CLK, Q => n635, QN 
                           => n2870);
   REGS_reg_61_3_inst : DFF_X1 port map( D => n12360, CK => CLK, Q => n636, QN 
                           => n2871);
   REGS_reg_61_2_inst : DFF_X1 port map( D => n12359, CK => CLK, Q => n637, QN 
                           => n2872);
   REGS_reg_61_1_inst : DFF_X1 port map( D => n12358, CK => CLK, Q => n638, QN 
                           => n2873);
   REGS_reg_61_0_inst : DFF_X1 port map( D => n12357, CK => CLK, Q => n639, QN 
                           => n2874);
   REGS_reg_59_23_inst : DFF_X1 port map( D => n12444, CK => CLK, Q => n16789, 
                           QN => n4714);
   REGS_reg_59_22_inst : DFF_X1 port map( D => n12443, CK => CLK, Q => n16788, 
                           QN => n4715);
   REGS_reg_59_21_inst : DFF_X1 port map( D => n12442, CK => CLK, Q => n16787, 
                           QN => n4716);
   REGS_reg_59_20_inst : DFF_X1 port map( D => n12441, CK => CLK, Q => n16786, 
                           QN => n4717);
   REGS_reg_59_19_inst : DFF_X1 port map( D => n12440, CK => CLK, Q => n16785, 
                           QN => n4718);
   REGS_reg_59_18_inst : DFF_X1 port map( D => n12439, CK => CLK, Q => n16784, 
                           QN => n4719);
   REGS_reg_59_17_inst : DFF_X1 port map( D => n12438, CK => CLK, Q => n16783, 
                           QN => n4720);
   REGS_reg_59_16_inst : DFF_X1 port map( D => n12437, CK => CLK, Q => n16782, 
                           QN => n4721);
   REGS_reg_59_15_inst : DFF_X1 port map( D => n12436, CK => CLK, Q => n16781, 
                           QN => n4722);
   REGS_reg_59_14_inst : DFF_X1 port map( D => n12435, CK => CLK, Q => n16780, 
                           QN => n4723);
   REGS_reg_59_13_inst : DFF_X1 port map( D => n12434, CK => CLK, Q => n16779, 
                           QN => n4724);
   REGS_reg_59_12_inst : DFF_X1 port map( D => n12433, CK => CLK, Q => n16778, 
                           QN => n4725);
   REGS_reg_59_11_inst : DFF_X1 port map( D => n12432, CK => CLK, Q => n16777, 
                           QN => n4726);
   REGS_reg_59_10_inst : DFF_X1 port map( D => n12431, CK => CLK, Q => n16776, 
                           QN => n4727);
   REGS_reg_59_9_inst : DFF_X1 port map( D => n12430, CK => CLK, Q => n16775, 
                           QN => n4728);
   REGS_reg_59_8_inst : DFF_X1 port map( D => n12429, CK => CLK, Q => n16774, 
                           QN => n4729);
   REGS_reg_59_7_inst : DFF_X1 port map( D => n12428, CK => CLK, Q => n16773, 
                           QN => n4730);
   REGS_reg_59_6_inst : DFF_X1 port map( D => n12427, CK => CLK, Q => n16772, 
                           QN => n4731);
   REGS_reg_59_5_inst : DFF_X1 port map( D => n12426, CK => CLK, Q => n16771, 
                           QN => n4732);
   REGS_reg_59_4_inst : DFF_X1 port map( D => n12425, CK => CLK, Q => n16770, 
                           QN => n4733);
   REGS_reg_59_3_inst : DFF_X1 port map( D => n12424, CK => CLK, Q => n16769, 
                           QN => n4734);
   REGS_reg_59_2_inst : DFF_X1 port map( D => n12423, CK => CLK, Q => n16768, 
                           QN => n4735);
   REGS_reg_59_1_inst : DFF_X1 port map( D => n12422, CK => CLK, Q => n16767, 
                           QN => n4736);
   REGS_reg_59_0_inst : DFF_X1 port map( D => n12421, CK => CLK, Q => n16766, 
                           QN => n4737);
   REGS_reg_58_23_inst : DFF_X1 port map( D => n12476, CK => CLK, Q => n_1566, 
                           QN => n2875);
   REGS_reg_58_22_inst : DFF_X1 port map( D => n12475, CK => CLK, Q => n_1567, 
                           QN => n2876);
   REGS_reg_58_21_inst : DFF_X1 port map( D => n12474, CK => CLK, Q => n_1568, 
                           QN => n2877);
   REGS_reg_58_20_inst : DFF_X1 port map( D => n12473, CK => CLK, Q => n_1569, 
                           QN => n2878);
   REGS_reg_58_19_inst : DFF_X1 port map( D => n12472, CK => CLK, Q => n_1570, 
                           QN => n2879);
   REGS_reg_58_18_inst : DFF_X1 port map( D => n12471, CK => CLK, Q => n_1571, 
                           QN => n2880);
   REGS_reg_58_17_inst : DFF_X1 port map( D => n12470, CK => CLK, Q => n_1572, 
                           QN => n2881);
   REGS_reg_58_16_inst : DFF_X1 port map( D => n12469, CK => CLK, Q => n_1573, 
                           QN => n2882);
   REGS_reg_58_15_inst : DFF_X1 port map( D => n12468, CK => CLK, Q => n_1574, 
                           QN => n2883);
   REGS_reg_58_14_inst : DFF_X1 port map( D => n12467, CK => CLK, Q => n_1575, 
                           QN => n2884);
   REGS_reg_58_13_inst : DFF_X1 port map( D => n12466, CK => CLK, Q => n_1576, 
                           QN => n2885);
   REGS_reg_58_12_inst : DFF_X1 port map( D => n12465, CK => CLK, Q => n_1577, 
                           QN => n2886);
   REGS_reg_58_11_inst : DFF_X1 port map( D => n12464, CK => CLK, Q => n_1578, 
                           QN => n2907);
   REGS_reg_58_10_inst : DFF_X1 port map( D => n12463, CK => CLK, Q => n_1579, 
                           QN => n2908);
   REGS_reg_58_9_inst : DFF_X1 port map( D => n12462, CK => CLK, Q => n_1580, 
                           QN => n2925);
   REGS_reg_58_8_inst : DFF_X1 port map( D => n12461, CK => CLK, Q => n_1581, 
                           QN => n2926);
   REGS_reg_58_7_inst : DFF_X1 port map( D => n12460, CK => CLK, Q => n_1582, 
                           QN => n2927);
   REGS_reg_58_6_inst : DFF_X1 port map( D => n12459, CK => CLK, Q => n_1583, 
                           QN => n2928);
   REGS_reg_58_5_inst : DFF_X1 port map( D => n12458, CK => CLK, Q => n_1584, 
                           QN => n2929);
   REGS_reg_58_4_inst : DFF_X1 port map( D => n12457, CK => CLK, Q => n_1585, 
                           QN => n2930);
   REGS_reg_58_3_inst : DFF_X1 port map( D => n12456, CK => CLK, Q => n_1586, 
                           QN => n2931);
   REGS_reg_58_2_inst : DFF_X1 port map( D => n12455, CK => CLK, Q => n_1587, 
                           QN => n2932);
   REGS_reg_58_1_inst : DFF_X1 port map( D => n12454, CK => CLK, Q => n_1588, 
                           QN => n2933);
   REGS_reg_58_0_inst : DFF_X1 port map( D => n12453, CK => CLK, Q => n_1589, 
                           QN => n2934);
   REGS_reg_57_23_inst : DFF_X1 port map( D => n12508, CK => CLK, Q => n_1590, 
                           QN => n2935);
   REGS_reg_57_22_inst : DFF_X1 port map( D => n12507, CK => CLK, Q => n_1591, 
                           QN => n2936);
   REGS_reg_57_21_inst : DFF_X1 port map( D => n12506, CK => CLK, Q => n_1592, 
                           QN => n2937);
   REGS_reg_57_20_inst : DFF_X1 port map( D => n12505, CK => CLK, Q => n_1593, 
                           QN => n2938);
   REGS_reg_57_19_inst : DFF_X1 port map( D => n12504, CK => CLK, Q => n_1594, 
                           QN => n2939);
   REGS_reg_57_18_inst : DFF_X1 port map( D => n12503, CK => CLK, Q => n_1595, 
                           QN => n2940);
   REGS_reg_57_17_inst : DFF_X1 port map( D => n12502, CK => CLK, Q => n_1596, 
                           QN => n2941);
   REGS_reg_57_16_inst : DFF_X1 port map( D => n12501, CK => CLK, Q => n_1597, 
                           QN => n2942);
   REGS_reg_57_15_inst : DFF_X1 port map( D => n12500, CK => CLK, Q => n_1598, 
                           QN => n2943);
   REGS_reg_57_14_inst : DFF_X1 port map( D => n12499, CK => CLK, Q => n_1599, 
                           QN => n2944);
   REGS_reg_57_13_inst : DFF_X1 port map( D => n12498, CK => CLK, Q => n_1600, 
                           QN => n2945);
   REGS_reg_57_12_inst : DFF_X1 port map( D => n12497, CK => CLK, Q => n_1601, 
                           QN => n2946);
   REGS_reg_57_11_inst : DFF_X1 port map( D => n12496, CK => CLK, Q => n_1602, 
                           QN => n2947);
   REGS_reg_57_10_inst : DFF_X1 port map( D => n12495, CK => CLK, Q => n_1603, 
                           QN => n2948);
   REGS_reg_57_9_inst : DFF_X1 port map( D => n12494, CK => CLK, Q => n_1604, 
                           QN => n2949);
   REGS_reg_57_8_inst : DFF_X1 port map( D => n12493, CK => CLK, Q => n_1605, 
                           QN => n2950);
   REGS_reg_57_7_inst : DFF_X1 port map( D => n12492, CK => CLK, Q => n_1606, 
                           QN => n2951);
   REGS_reg_57_6_inst : DFF_X1 port map( D => n12491, CK => CLK, Q => n_1607, 
                           QN => n2952);
   REGS_reg_57_5_inst : DFF_X1 port map( D => n12490, CK => CLK, Q => n_1608, 
                           QN => n2953);
   REGS_reg_57_4_inst : DFF_X1 port map( D => n12489, CK => CLK, Q => n_1609, 
                           QN => n2954);
   REGS_reg_57_3_inst : DFF_X1 port map( D => n12488, CK => CLK, Q => n_1610, 
                           QN => n2955);
   REGS_reg_57_2_inst : DFF_X1 port map( D => n12487, CK => CLK, Q => n_1611, 
                           QN => n2956);
   REGS_reg_57_1_inst : DFF_X1 port map( D => n12486, CK => CLK, Q => n_1612, 
                           QN => n2957);
   REGS_reg_57_0_inst : DFF_X1 port map( D => n12485, CK => CLK, Q => n_1613, 
                           QN => n2958);
   REGS_reg_56_23_inst : DFF_X1 port map( D => n12540, CK => CLK, Q => n640, QN
                           => n2959);
   REGS_reg_56_22_inst : DFF_X1 port map( D => n12539, CK => CLK, Q => n641, QN
                           => n2960);
   REGS_reg_56_21_inst : DFF_X1 port map( D => n12538, CK => CLK, Q => n642, QN
                           => n2961);
   REGS_reg_56_20_inst : DFF_X1 port map( D => n12537, CK => CLK, Q => n643, QN
                           => n2962);
   REGS_reg_56_19_inst : DFF_X1 port map( D => n12536, CK => CLK, Q => n644, QN
                           => n2963);
   REGS_reg_56_18_inst : DFF_X1 port map( D => n12535, CK => CLK, Q => n645, QN
                           => n2964);
   REGS_reg_56_17_inst : DFF_X1 port map( D => n12534, CK => CLK, Q => n646, QN
                           => n2965);
   REGS_reg_56_16_inst : DFF_X1 port map( D => n12533, CK => CLK, Q => n647, QN
                           => n2966);
   REGS_reg_56_15_inst : DFF_X1 port map( D => n12532, CK => CLK, Q => n648, QN
                           => n2967);
   REGS_reg_56_14_inst : DFF_X1 port map( D => n12531, CK => CLK, Q => n649, QN
                           => n2968);
   REGS_reg_56_13_inst : DFF_X1 port map( D => n12530, CK => CLK, Q => n650, QN
                           => n2969);
   REGS_reg_56_12_inst : DFF_X1 port map( D => n12529, CK => CLK, Q => n651, QN
                           => n2970);
   REGS_reg_56_11_inst : DFF_X1 port map( D => n12528, CK => CLK, Q => n652, QN
                           => n2971);
   REGS_reg_56_10_inst : DFF_X1 port map( D => n12527, CK => CLK, Q => n653, QN
                           => n2972);
   REGS_reg_56_9_inst : DFF_X1 port map( D => n12526, CK => CLK, Q => n654, QN 
                           => n2973);
   REGS_reg_56_8_inst : DFF_X1 port map( D => n12525, CK => CLK, Q => n655, QN 
                           => n2974);
   REGS_reg_56_7_inst : DFF_X1 port map( D => n12524, CK => CLK, Q => n656, QN 
                           => n2975);
   REGS_reg_56_6_inst : DFF_X1 port map( D => n12523, CK => CLK, Q => n657, QN 
                           => n2976);
   REGS_reg_56_5_inst : DFF_X1 port map( D => n12522, CK => CLK, Q => n658, QN 
                           => n2977);
   REGS_reg_56_4_inst : DFF_X1 port map( D => n12521, CK => CLK, Q => n659, QN 
                           => n2978);
   REGS_reg_56_3_inst : DFF_X1 port map( D => n12520, CK => CLK, Q => n660, QN 
                           => n3027);
   REGS_reg_56_2_inst : DFF_X1 port map( D => n12519, CK => CLK, Q => n661, QN 
                           => n3028);
   REGS_reg_56_1_inst : DFF_X1 port map( D => n12518, CK => CLK, Q => n662, QN 
                           => n3029);
   REGS_reg_56_0_inst : DFF_X1 port map( D => n12517, CK => CLK, Q => n663, QN 
                           => n3030);
   REGS_reg_55_23_inst : DFF_X1 port map( D => n12572, CK => CLK, Q => n664, QN
                           => n3031);
   REGS_reg_55_22_inst : DFF_X1 port map( D => n12571, CK => CLK, Q => n665, QN
                           => n3032);
   REGS_reg_55_21_inst : DFF_X1 port map( D => n12570, CK => CLK, Q => n666, QN
                           => n3033);
   REGS_reg_55_20_inst : DFF_X1 port map( D => n12569, CK => CLK, Q => n667, QN
                           => n3034);
   REGS_reg_55_19_inst : DFF_X1 port map( D => n12568, CK => CLK, Q => n668, QN
                           => n3035);
   REGS_reg_55_18_inst : DFF_X1 port map( D => n12567, CK => CLK, Q => n669, QN
                           => n3036);
   REGS_reg_55_17_inst : DFF_X1 port map( D => n12566, CK => CLK, Q => n670, QN
                           => n3037);
   REGS_reg_55_16_inst : DFF_X1 port map( D => n12565, CK => CLK, Q => n671, QN
                           => n3038);
   REGS_reg_55_15_inst : DFF_X1 port map( D => n12564, CK => CLK, Q => n672, QN
                           => n3039);
   REGS_reg_55_14_inst : DFF_X1 port map( D => n12563, CK => CLK, Q => n673, QN
                           => n3040);
   REGS_reg_55_13_inst : DFF_X1 port map( D => n12562, CK => CLK, Q => n674, QN
                           => n3041);
   REGS_reg_55_12_inst : DFF_X1 port map( D => n12561, CK => CLK, Q => n675, QN
                           => n3042);
   REGS_reg_55_11_inst : DFF_X1 port map( D => n12560, CK => CLK, Q => n676, QN
                           => n3043);
   REGS_reg_55_10_inst : DFF_X1 port map( D => n12559, CK => CLK, Q => n677, QN
                           => n3044);
   REGS_reg_55_9_inst : DFF_X1 port map( D => n12558, CK => CLK, Q => n678, QN 
                           => n3045);
   REGS_reg_55_8_inst : DFF_X1 port map( D => n12557, CK => CLK, Q => n679, QN 
                           => n3046);
   REGS_reg_55_7_inst : DFF_X1 port map( D => n12556, CK => CLK, Q => n680, QN 
                           => n3047);
   REGS_reg_55_6_inst : DFF_X1 port map( D => n12555, CK => CLK, Q => n681, QN 
                           => n3048);
   REGS_reg_55_5_inst : DFF_X1 port map( D => n12554, CK => CLK, Q => n682, QN 
                           => n3049);
   REGS_reg_55_4_inst : DFF_X1 port map( D => n12553, CK => CLK, Q => n683, QN 
                           => n3050);
   REGS_reg_55_3_inst : DFF_X1 port map( D => n12552, CK => CLK, Q => n684, QN 
                           => n3051);
   REGS_reg_55_2_inst : DFF_X1 port map( D => n12551, CK => CLK, Q => n685, QN 
                           => n3052);
   REGS_reg_55_1_inst : DFF_X1 port map( D => n12550, CK => CLK, Q => n686, QN 
                           => n3053);
   REGS_reg_55_0_inst : DFF_X1 port map( D => n12549, CK => CLK, Q => n687, QN 
                           => n3054);
   REGS_reg_54_23_inst : DFF_X1 port map( D => n12604, CK => CLK, Q => n688, QN
                           => n3055);
   REGS_reg_54_22_inst : DFF_X1 port map( D => n12603, CK => CLK, Q => n689, QN
                           => n3056);
   REGS_reg_54_21_inst : DFF_X1 port map( D => n12602, CK => CLK, Q => n690, QN
                           => n3057);
   REGS_reg_54_20_inst : DFF_X1 port map( D => n12601, CK => CLK, Q => n691, QN
                           => n3058);
   REGS_reg_54_19_inst : DFF_X1 port map( D => n12600, CK => CLK, Q => n692, QN
                           => n3059);
   REGS_reg_54_18_inst : DFF_X1 port map( D => n12599, CK => CLK, Q => n693, QN
                           => n3060);
   REGS_reg_54_17_inst : DFF_X1 port map( D => n12598, CK => CLK, Q => n694, QN
                           => n3061);
   REGS_reg_54_16_inst : DFF_X1 port map( D => n12597, CK => CLK, Q => n695, QN
                           => n3062);
   REGS_reg_54_15_inst : DFF_X1 port map( D => n12596, CK => CLK, Q => n696, QN
                           => n3063);
   REGS_reg_54_14_inst : DFF_X1 port map( D => n12595, CK => CLK, Q => n697, QN
                           => n3064);
   REGS_reg_54_13_inst : DFF_X1 port map( D => n12594, CK => CLK, Q => n698, QN
                           => n3065);
   REGS_reg_54_12_inst : DFF_X1 port map( D => n12593, CK => CLK, Q => n699, QN
                           => n3066);
   REGS_reg_54_11_inst : DFF_X1 port map( D => n12592, CK => CLK, Q => n700, QN
                           => n3067);
   REGS_reg_54_10_inst : DFF_X1 port map( D => n12591, CK => CLK, Q => n701, QN
                           => n3068);
   REGS_reg_54_9_inst : DFF_X1 port map( D => n12590, CK => CLK, Q => n702, QN 
                           => n3069);
   REGS_reg_54_8_inst : DFF_X1 port map( D => n12589, CK => CLK, Q => n703, QN 
                           => n3070);
   REGS_reg_54_7_inst : DFF_X1 port map( D => n12588, CK => CLK, Q => n704, QN 
                           => n3071);
   REGS_reg_54_6_inst : DFF_X1 port map( D => n12587, CK => CLK, Q => n705, QN 
                           => n3072);
   REGS_reg_54_5_inst : DFF_X1 port map( D => n12586, CK => CLK, Q => n706, QN 
                           => n3073);
   REGS_reg_54_4_inst : DFF_X1 port map( D => n12585, CK => CLK, Q => n707, QN 
                           => n3074);
   REGS_reg_54_3_inst : DFF_X1 port map( D => n12584, CK => CLK, Q => n708, QN 
                           => n3075);
   REGS_reg_54_2_inst : DFF_X1 port map( D => n12583, CK => CLK, Q => n709, QN 
                           => n3076);
   REGS_reg_54_1_inst : DFF_X1 port map( D => n12582, CK => CLK, Q => n710, QN 
                           => n3077);
   REGS_reg_54_0_inst : DFF_X1 port map( D => n12581, CK => CLK, Q => n711, QN 
                           => n3078);
   REGS_reg_53_23_inst : DFF_X1 port map( D => n12636, CK => CLK, Q => n712, QN
                           => n3079);
   REGS_reg_53_22_inst : DFF_X1 port map( D => n12635, CK => CLK, Q => n713, QN
                           => n3080);
   REGS_reg_53_21_inst : DFF_X1 port map( D => n12634, CK => CLK, Q => n714, QN
                           => n3081);
   REGS_reg_53_20_inst : DFF_X1 port map( D => n12633, CK => CLK, Q => n715, QN
                           => n3082);
   REGS_reg_53_19_inst : DFF_X1 port map( D => n12632, CK => CLK, Q => n716, QN
                           => n3083);
   REGS_reg_53_18_inst : DFF_X1 port map( D => n12631, CK => CLK, Q => n717, QN
                           => n3084);
   REGS_reg_53_17_inst : DFF_X1 port map( D => n12630, CK => CLK, Q => n718, QN
                           => n3085);
   REGS_reg_53_16_inst : DFF_X1 port map( D => n12629, CK => CLK, Q => n719, QN
                           => n3086);
   REGS_reg_53_15_inst : DFF_X1 port map( D => n12628, CK => CLK, Q => n720, QN
                           => n3087);
   REGS_reg_53_14_inst : DFF_X1 port map( D => n12627, CK => CLK, Q => n721, QN
                           => n3088);
   REGS_reg_53_13_inst : DFF_X1 port map( D => n12626, CK => CLK, Q => n722, QN
                           => n3089);
   REGS_reg_53_12_inst : DFF_X1 port map( D => n12625, CK => CLK, Q => n723, QN
                           => n3090);
   REGS_reg_53_11_inst : DFF_X1 port map( D => n12624, CK => CLK, Q => n724, QN
                           => n3091);
   REGS_reg_53_10_inst : DFF_X1 port map( D => n12623, CK => CLK, Q => n725, QN
                           => n3092);
   REGS_reg_53_9_inst : DFF_X1 port map( D => n12622, CK => CLK, Q => n726, QN 
                           => n3093);
   REGS_reg_53_8_inst : DFF_X1 port map( D => n12621, CK => CLK, Q => n727, QN 
                           => n3094);
   REGS_reg_53_7_inst : DFF_X1 port map( D => n12620, CK => CLK, Q => n728, QN 
                           => n3095);
   REGS_reg_53_6_inst : DFF_X1 port map( D => n12619, CK => CLK, Q => n729, QN 
                           => n3096);
   REGS_reg_53_5_inst : DFF_X1 port map( D => n12618, CK => CLK, Q => n730, QN 
                           => n3097);
   REGS_reg_53_4_inst : DFF_X1 port map( D => n12617, CK => CLK, Q => n731, QN 
                           => n3098);
   REGS_reg_53_3_inst : DFF_X1 port map( D => n12616, CK => CLK, Q => n732, QN 
                           => n3123);
   REGS_reg_53_2_inst : DFF_X1 port map( D => n12615, CK => CLK, Q => n733, QN 
                           => n3124);
   REGS_reg_53_1_inst : DFF_X1 port map( D => n12614, CK => CLK, Q => n734, QN 
                           => n3125);
   REGS_reg_53_0_inst : DFF_X1 port map( D => n12613, CK => CLK, Q => n735, QN 
                           => n3126);
   REGS_reg_52_23_inst : DFF_X1 port map( D => n12668, CK => CLK, Q => n16765, 
                           QN => n4738);
   REGS_reg_52_22_inst : DFF_X1 port map( D => n12667, CK => CLK, Q => n16764, 
                           QN => n4739);
   REGS_reg_52_21_inst : DFF_X1 port map( D => n12666, CK => CLK, Q => n16763, 
                           QN => n4740);
   REGS_reg_52_20_inst : DFF_X1 port map( D => n12665, CK => CLK, Q => n16762, 
                           QN => n4741);
   REGS_reg_52_19_inst : DFF_X1 port map( D => n12664, CK => CLK, Q => n16761, 
                           QN => n4742);
   REGS_reg_52_18_inst : DFF_X1 port map( D => n12663, CK => CLK, Q => n16760, 
                           QN => n4743);
   REGS_reg_52_17_inst : DFF_X1 port map( D => n12662, CK => CLK, Q => n16759, 
                           QN => n4744);
   REGS_reg_52_16_inst : DFF_X1 port map( D => n12661, CK => CLK, Q => n16758, 
                           QN => n4745);
   REGS_reg_52_15_inst : DFF_X1 port map( D => n12660, CK => CLK, Q => n16757, 
                           QN => n4746);
   REGS_reg_52_14_inst : DFF_X1 port map( D => n12659, CK => CLK, Q => n16756, 
                           QN => n4747);
   REGS_reg_52_13_inst : DFF_X1 port map( D => n12658, CK => CLK, Q => n16755, 
                           QN => n4748);
   REGS_reg_52_12_inst : DFF_X1 port map( D => n12657, CK => CLK, Q => n16754, 
                           QN => n4749);
   REGS_reg_52_11_inst : DFF_X1 port map( D => n12656, CK => CLK, Q => n16753, 
                           QN => n4750);
   REGS_reg_52_10_inst : DFF_X1 port map( D => n12655, CK => CLK, Q => n16752, 
                           QN => n4751);
   REGS_reg_52_9_inst : DFF_X1 port map( D => n12654, CK => CLK, Q => n16751, 
                           QN => n4752);
   REGS_reg_52_8_inst : DFF_X1 port map( D => n12653, CK => CLK, Q => n16750, 
                           QN => n4753);
   REGS_reg_52_7_inst : DFF_X1 port map( D => n12652, CK => CLK, Q => n16749, 
                           QN => n4754);
   REGS_reg_52_6_inst : DFF_X1 port map( D => n12651, CK => CLK, Q => n16748, 
                           QN => n4755);
   REGS_reg_52_5_inst : DFF_X1 port map( D => n12650, CK => CLK, Q => n16747, 
                           QN => n4756);
   REGS_reg_52_4_inst : DFF_X1 port map( D => n12649, CK => CLK, Q => n16746, 
                           QN => n4757);
   REGS_reg_52_3_inst : DFF_X1 port map( D => n12648, CK => CLK, Q => n16745, 
                           QN => n4758);
   REGS_reg_52_2_inst : DFF_X1 port map( D => n12647, CK => CLK, Q => n16744, 
                           QN => n4759);
   REGS_reg_52_1_inst : DFF_X1 port map( D => n12646, CK => CLK, Q => n16743, 
                           QN => n4760);
   REGS_reg_52_0_inst : DFF_X1 port map( D => n12645, CK => CLK, Q => n16742, 
                           QN => n4761);
   REGS_reg_51_23_inst : DFF_X1 port map( D => n12700, CK => CLK, Q => n16741, 
                           QN => n4762);
   REGS_reg_51_22_inst : DFF_X1 port map( D => n12699, CK => CLK, Q => n16740, 
                           QN => n4763);
   REGS_reg_51_21_inst : DFF_X1 port map( D => n12698, CK => CLK, Q => n16739, 
                           QN => n4764);
   REGS_reg_51_20_inst : DFF_X1 port map( D => n12697, CK => CLK, Q => n16738, 
                           QN => n4765);
   REGS_reg_51_19_inst : DFF_X1 port map( D => n12696, CK => CLK, Q => n16737, 
                           QN => n4766);
   REGS_reg_51_18_inst : DFF_X1 port map( D => n12695, CK => CLK, Q => n16736, 
                           QN => n4767);
   REGS_reg_51_17_inst : DFF_X1 port map( D => n12694, CK => CLK, Q => n16735, 
                           QN => n4768);
   REGS_reg_51_16_inst : DFF_X1 port map( D => n12693, CK => CLK, Q => n16734, 
                           QN => n4769);
   REGS_reg_51_15_inst : DFF_X1 port map( D => n12692, CK => CLK, Q => n16733, 
                           QN => n4770);
   REGS_reg_51_14_inst : DFF_X1 port map( D => n12691, CK => CLK, Q => n16732, 
                           QN => n4771);
   REGS_reg_51_13_inst : DFF_X1 port map( D => n12690, CK => CLK, Q => n16731, 
                           QN => n4772);
   REGS_reg_51_12_inst : DFF_X1 port map( D => n12689, CK => CLK, Q => n16730, 
                           QN => n4773);
   REGS_reg_51_11_inst : DFF_X1 port map( D => n12688, CK => CLK, Q => n16729, 
                           QN => n4774);
   REGS_reg_51_10_inst : DFF_X1 port map( D => n12687, CK => CLK, Q => n16728, 
                           QN => n4775);
   REGS_reg_51_9_inst : DFF_X1 port map( D => n12686, CK => CLK, Q => n16727, 
                           QN => n4776);
   REGS_reg_51_8_inst : DFF_X1 port map( D => n12685, CK => CLK, Q => n16726, 
                           QN => n4777);
   REGS_reg_51_7_inst : DFF_X1 port map( D => n12684, CK => CLK, Q => n16725, 
                           QN => n4778);
   REGS_reg_51_6_inst : DFF_X1 port map( D => n12683, CK => CLK, Q => n16724, 
                           QN => n4779);
   REGS_reg_51_5_inst : DFF_X1 port map( D => n12682, CK => CLK, Q => n16723, 
                           QN => n4780);
   REGS_reg_51_4_inst : DFF_X1 port map( D => n12681, CK => CLK, Q => n16722, 
                           QN => n4781);
   REGS_reg_51_3_inst : DFF_X1 port map( D => n12680, CK => CLK, Q => n16721, 
                           QN => n4782);
   REGS_reg_51_2_inst : DFF_X1 port map( D => n12679, CK => CLK, Q => n16720, 
                           QN => n4783);
   REGS_reg_51_1_inst : DFF_X1 port map( D => n12678, CK => CLK, Q => n16719, 
                           QN => n4784);
   REGS_reg_51_0_inst : DFF_X1 port map( D => n12677, CK => CLK, Q => n16718, 
                           QN => n4785);
   REGS_reg_50_23_inst : DFF_X1 port map( D => n12732, CK => CLK, Q => n53124, 
                           QN => n3127);
   REGS_reg_50_22_inst : DFF_X1 port map( D => n12731, CK => CLK, Q => n53125, 
                           QN => n3128);
   REGS_reg_50_21_inst : DFF_X1 port map( D => n12730, CK => CLK, Q => n53126, 
                           QN => n3129);
   REGS_reg_50_20_inst : DFF_X1 port map( D => n12729, CK => CLK, Q => n53127, 
                           QN => n3130);
   REGS_reg_50_19_inst : DFF_X1 port map( D => n12728, CK => CLK, Q => n53128, 
                           QN => n3131);
   REGS_reg_50_18_inst : DFF_X1 port map( D => n12727, CK => CLK, Q => n53129, 
                           QN => n3132);
   REGS_reg_50_17_inst : DFF_X1 port map( D => n12726, CK => CLK, Q => n53130, 
                           QN => n3133);
   REGS_reg_50_16_inst : DFF_X1 port map( D => n12725, CK => CLK, Q => n53131, 
                           QN => n3134);
   REGS_reg_50_15_inst : DFF_X1 port map( D => n12724, CK => CLK, Q => n53132, 
                           QN => n3135);
   REGS_reg_50_14_inst : DFF_X1 port map( D => n12723, CK => CLK, Q => n53133, 
                           QN => n3136);
   REGS_reg_50_13_inst : DFF_X1 port map( D => n12722, CK => CLK, Q => n53134, 
                           QN => n3137);
   REGS_reg_50_12_inst : DFF_X1 port map( D => n12721, CK => CLK, Q => n53135, 
                           QN => n3138);
   REGS_reg_50_11_inst : DFF_X1 port map( D => n12720, CK => CLK, Q => n53136, 
                           QN => n3139);
   REGS_reg_50_10_inst : DFF_X1 port map( D => n12719, CK => CLK, Q => n53137, 
                           QN => n3140);
   REGS_reg_50_9_inst : DFF_X1 port map( D => n12718, CK => CLK, Q => n53138, 
                           QN => n3141);
   REGS_reg_50_8_inst : DFF_X1 port map( D => n12717, CK => CLK, Q => n53139, 
                           QN => n3142);
   REGS_reg_50_7_inst : DFF_X1 port map( D => n12716, CK => CLK, Q => n53140, 
                           QN => n3143);
   REGS_reg_50_6_inst : DFF_X1 port map( D => n12715, CK => CLK, Q => n53141, 
                           QN => n3144);
   REGS_reg_50_5_inst : DFF_X1 port map( D => n12714, CK => CLK, Q => n53142, 
                           QN => n3145);
   REGS_reg_50_4_inst : DFF_X1 port map( D => n12713, CK => CLK, Q => n53143, 
                           QN => n3146);
   REGS_reg_50_3_inst : DFF_X1 port map( D => n12712, CK => CLK, Q => n53144, 
                           QN => n3147);
   REGS_reg_50_2_inst : DFF_X1 port map( D => n12711, CK => CLK, Q => n53145, 
                           QN => n3148);
   REGS_reg_50_1_inst : DFF_X1 port map( D => n12710, CK => CLK, Q => n53146, 
                           QN => n3149);
   REGS_reg_50_0_inst : DFF_X1 port map( D => n12709, CK => CLK, Q => n53147, 
                           QN => n3150);
   REGS_reg_48_9_inst : DFF_X1 port map( D => n12782, CK => CLK, Q => n53186, 
                           QN => n3151);
   REGS_reg_48_8_inst : DFF_X1 port map( D => n12781, CK => CLK, Q => n53187, 
                           QN => n3152);
   REGS_reg_48_7_inst : DFF_X1 port map( D => n12780, CK => CLK, Q => n53188, 
                           QN => n3153);
   REGS_reg_48_6_inst : DFF_X1 port map( D => n12779, CK => CLK, Q => n53189, 
                           QN => n3154);
   REGS_reg_48_5_inst : DFF_X1 port map( D => n12778, CK => CLK, Q => n53190, 
                           QN => n3155);
   REGS_reg_48_4_inst : DFF_X1 port map( D => n12777, CK => CLK, Q => n53191, 
                           QN => n3156);
   REGS_reg_48_3_inst : DFF_X1 port map( D => n12776, CK => CLK, Q => n53192, 
                           QN => n3157);
   REGS_reg_48_2_inst : DFF_X1 port map( D => n12775, CK => CLK, Q => n53193, 
                           QN => n3158);
   REGS_reg_48_1_inst : DFF_X1 port map( D => n12774, CK => CLK, Q => n53194, 
                           QN => n3159);
   REGS_reg_48_0_inst : DFF_X1 port map( D => n12773, CK => CLK, Q => n53195, 
                           QN => n3160);
   REGS_reg_47_23_inst : DFF_X1 port map( D => n12828, CK => CLK, Q => n16717, 
                           QN => n4824);
   REGS_reg_47_22_inst : DFF_X1 port map( D => n12827, CK => CLK, Q => n16716, 
                           QN => n4825);
   REGS_reg_47_21_inst : DFF_X1 port map( D => n12826, CK => CLK, Q => n16715, 
                           QN => n4826);
   REGS_reg_47_20_inst : DFF_X1 port map( D => n12825, CK => CLK, Q => n16714, 
                           QN => n4827);
   REGS_reg_47_19_inst : DFF_X1 port map( D => n12824, CK => CLK, Q => n16713, 
                           QN => n4828);
   REGS_reg_47_18_inst : DFF_X1 port map( D => n12823, CK => CLK, Q => n16712, 
                           QN => n4829);
   REGS_reg_47_17_inst : DFF_X1 port map( D => n12822, CK => CLK, Q => n16711, 
                           QN => n4830);
   REGS_reg_47_16_inst : DFF_X1 port map( D => n12821, CK => CLK, Q => n16710, 
                           QN => n4831);
   REGS_reg_47_15_inst : DFF_X1 port map( D => n12820, CK => CLK, Q => n16709, 
                           QN => n4832);
   REGS_reg_47_14_inst : DFF_X1 port map( D => n12819, CK => CLK, Q => n16708, 
                           QN => n4833);
   REGS_reg_47_13_inst : DFF_X1 port map( D => n12818, CK => CLK, Q => n16308, 
                           QN => n3161);
   REGS_reg_47_12_inst : DFF_X1 port map( D => n12817, CK => CLK, Q => n16306, 
                           QN => n3162);
   REGS_reg_47_11_inst : DFF_X1 port map( D => n12816, CK => CLK, Q => n16304, 
                           QN => n3163);
   REGS_reg_47_10_inst : DFF_X1 port map( D => n12815, CK => CLK, Q => n16302, 
                           QN => n3164);
   REGS_reg_47_9_inst : DFF_X1 port map( D => n12814, CK => CLK, Q => n16300, 
                           QN => n3165);
   REGS_reg_47_8_inst : DFF_X1 port map( D => n12813, CK => CLK, Q => n16298, 
                           QN => n3166);
   REGS_reg_47_7_inst : DFF_X1 port map( D => n12812, CK => CLK, Q => n16334, 
                           QN => n3167);
   REGS_reg_47_6_inst : DFF_X1 port map( D => n12811, CK => CLK, Q => n16332, 
                           QN => n3168);
   REGS_reg_47_5_inst : DFF_X1 port map( D => n12810, CK => CLK, Q => n16330, 
                           QN => n3169);
   REGS_reg_47_4_inst : DFF_X1 port map( D => n12809, CK => CLK, Q => n16328, 
                           QN => n3170);
   REGS_reg_47_3_inst : DFF_X1 port map( D => n12808, CK => CLK, Q => n16326, 
                           QN => n3171);
   REGS_reg_47_2_inst : DFF_X1 port map( D => n12807, CK => CLK, Q => n16324, 
                           QN => n3172);
   REGS_reg_47_1_inst : DFF_X1 port map( D => n12806, CK => CLK, Q => n16322, 
                           QN => n3173);
   REGS_reg_47_0_inst : DFF_X1 port map( D => n12805, CK => CLK, Q => n16320, 
                           QN => n3174);
   REGS_reg_46_23_inst : DFF_X1 port map( D => n12860, CK => CLK, Q => n16707, 
                           QN => n4834);
   REGS_reg_46_22_inst : DFF_X1 port map( D => n12859, CK => CLK, Q => n16706, 
                           QN => n4835);
   REGS_reg_46_21_inst : DFF_X1 port map( D => n12858, CK => CLK, Q => n16705, 
                           QN => n4836);
   REGS_reg_46_20_inst : DFF_X1 port map( D => n12857, CK => CLK, Q => n16704, 
                           QN => n4837);
   REGS_reg_46_19_inst : DFF_X1 port map( D => n12856, CK => CLK, Q => n16703, 
                           QN => n4838);
   REGS_reg_46_18_inst : DFF_X1 port map( D => n12855, CK => CLK, Q => n16702, 
                           QN => n4839);
   REGS_reg_46_17_inst : DFF_X1 port map( D => n12854, CK => CLK, Q => n16701, 
                           QN => n4840);
   REGS_reg_46_16_inst : DFF_X1 port map( D => n12853, CK => CLK, Q => n16700, 
                           QN => n4841);
   REGS_reg_46_15_inst : DFF_X1 port map( D => n12852, CK => CLK, Q => n16699, 
                           QN => n4842);
   REGS_reg_46_14_inst : DFF_X1 port map( D => n12851, CK => CLK, Q => n16698, 
                           QN => n4843);
   REGS_reg_46_13_inst : DFF_X1 port map( D => n12850, CK => CLK, Q => n16697, 
                           QN => n4844);
   REGS_reg_46_12_inst : DFF_X1 port map( D => n12849, CK => CLK, Q => n16696, 
                           QN => n4845);
   REGS_reg_46_11_inst : DFF_X1 port map( D => n12848, CK => CLK, Q => n16695, 
                           QN => n4846);
   REGS_reg_46_10_inst : DFF_X1 port map( D => n12847, CK => CLK, Q => n16694, 
                           QN => n4847);
   REGS_reg_46_9_inst : DFF_X1 port map( D => n12846, CK => CLK, Q => n16693, 
                           QN => n4848);
   REGS_reg_46_8_inst : DFF_X1 port map( D => n12845, CK => CLK, Q => n16692, 
                           QN => n4849);
   REGS_reg_46_7_inst : DFF_X1 port map( D => n12844, CK => CLK, Q => n16691, 
                           QN => n4850);
   REGS_reg_46_6_inst : DFF_X1 port map( D => n12843, CK => CLK, Q => n16690, 
                           QN => n4851);
   REGS_reg_46_5_inst : DFF_X1 port map( D => n12842, CK => CLK, Q => n16689, 
                           QN => n4852);
   REGS_reg_46_4_inst : DFF_X1 port map( D => n12841, CK => CLK, Q => n16688, 
                           QN => n4853);
   REGS_reg_46_3_inst : DFF_X1 port map( D => n12840, CK => CLK, Q => n16687, 
                           QN => n4854);
   REGS_reg_46_2_inst : DFF_X1 port map( D => n12839, CK => CLK, Q => n16686, 
                           QN => n4855);
   REGS_reg_46_1_inst : DFF_X1 port map( D => n12838, CK => CLK, Q => n16685, 
                           QN => n4856);
   REGS_reg_46_0_inst : DFF_X1 port map( D => n12837, CK => CLK, Q => n16684, 
                           QN => n4857);
   REGS_reg_45_23_inst : DFF_X1 port map( D => n12892, CK => CLK, Q => n736, QN
                           => n3175);
   REGS_reg_45_22_inst : DFF_X1 port map( D => n12891, CK => CLK, Q => n737, QN
                           => n3176);
   REGS_reg_45_21_inst : DFF_X1 port map( D => n12890, CK => CLK, Q => n738, QN
                           => n3177);
   REGS_reg_45_20_inst : DFF_X1 port map( D => n12889, CK => CLK, Q => n739, QN
                           => n3178);
   REGS_reg_45_19_inst : DFF_X1 port map( D => n12888, CK => CLK, Q => n740, QN
                           => n3179);
   REGS_reg_45_18_inst : DFF_X1 port map( D => n12887, CK => CLK, Q => n741, QN
                           => n3180);
   REGS_reg_45_17_inst : DFF_X1 port map( D => n12886, CK => CLK, Q => n742, QN
                           => n3181);
   REGS_reg_45_16_inst : DFF_X1 port map( D => n12885, CK => CLK, Q => n743, QN
                           => n3182);
   REGS_reg_45_15_inst : DFF_X1 port map( D => n12884, CK => CLK, Q => n744, QN
                           => n3183);
   REGS_reg_45_14_inst : DFF_X1 port map( D => n12883, CK => CLK, Q => n745, QN
                           => n3184);
   REGS_reg_45_13_inst : DFF_X1 port map( D => n12882, CK => CLK, Q => n746, QN
                           => n3185);
   REGS_reg_45_12_inst : DFF_X1 port map( D => n12881, CK => CLK, Q => n747, QN
                           => n3186);
   REGS_reg_45_11_inst : DFF_X1 port map( D => n12880, CK => CLK, Q => n748, QN
                           => n3187);
   REGS_reg_45_10_inst : DFF_X1 port map( D => n12879, CK => CLK, Q => n749, QN
                           => n3188);
   REGS_reg_45_9_inst : DFF_X1 port map( D => n12878, CK => CLK, Q => n750, QN 
                           => n3189);
   REGS_reg_45_8_inst : DFF_X1 port map( D => n12877, CK => CLK, Q => n751, QN 
                           => n3190);
   REGS_reg_45_7_inst : DFF_X1 port map( D => n12876, CK => CLK, Q => n752, QN 
                           => n3191);
   REGS_reg_45_6_inst : DFF_X1 port map( D => n12875, CK => CLK, Q => n753, QN 
                           => n3192);
   REGS_reg_45_5_inst : DFF_X1 port map( D => n12874, CK => CLK, Q => n754, QN 
                           => n3193);
   REGS_reg_45_4_inst : DFF_X1 port map( D => n12873, CK => CLK, Q => n755, QN 
                           => n3194);
   REGS_reg_45_3_inst : DFF_X1 port map( D => n12872, CK => CLK, Q => n756, QN 
                           => n3195);
   REGS_reg_45_2_inst : DFF_X1 port map( D => n12871, CK => CLK, Q => n757, QN 
                           => n3196);
   REGS_reg_45_1_inst : DFF_X1 port map( D => n12870, CK => CLK, Q => n758, QN 
                           => n3197);
   REGS_reg_45_0_inst : DFF_X1 port map( D => n12869, CK => CLK, Q => n759, QN 
                           => n3198);
   REGS_reg_44_9_inst : DFF_X1 port map( D => n12910, CK => CLK, Q => n_1614, 
                           QN => n3199);
   REGS_reg_44_8_inst : DFF_X1 port map( D => n12909, CK => CLK, Q => n_1615, 
                           QN => n3200);
   REGS_reg_44_7_inst : DFF_X1 port map( D => n12908, CK => CLK, Q => n_1616, 
                           QN => n3201);
   REGS_reg_44_6_inst : DFF_X1 port map( D => n12907, CK => CLK, Q => n_1617, 
                           QN => n3202);
   REGS_reg_44_5_inst : DFF_X1 port map( D => n12906, CK => CLK, Q => n_1618, 
                           QN => n3203);
   REGS_reg_44_4_inst : DFF_X1 port map( D => n12905, CK => CLK, Q => n_1619, 
                           QN => n3204);
   REGS_reg_44_3_inst : DFF_X1 port map( D => n12904, CK => CLK, Q => n_1620, 
                           QN => n3205);
   REGS_reg_44_2_inst : DFF_X1 port map( D => n12903, CK => CLK, Q => n_1621, 
                           QN => n3206);
   REGS_reg_44_1_inst : DFF_X1 port map( D => n12902, CK => CLK, Q => n_1622, 
                           QN => n3207);
   REGS_reg_44_0_inst : DFF_X1 port map( D => n12901, CK => CLK, Q => n_1623, 
                           QN => n3208);
   REGS_reg_43_23_inst : DFF_X1 port map( D => n12956, CK => CLK, Q => n16529, 
                           QN => n4858);
   REGS_reg_43_22_inst : DFF_X1 port map( D => n12955, CK => CLK, Q => n16528, 
                           QN => n4859);
   REGS_reg_43_21_inst : DFF_X1 port map( D => n12954, CK => CLK, Q => n16527, 
                           QN => n4860);
   REGS_reg_43_20_inst : DFF_X1 port map( D => n12953, CK => CLK, Q => n16526, 
                           QN => n4861);
   REGS_reg_43_19_inst : DFF_X1 port map( D => n12952, CK => CLK, Q => n16525, 
                           QN => n4862);
   REGS_reg_43_18_inst : DFF_X1 port map( D => n12951, CK => CLK, Q => n16524, 
                           QN => n4863);
   REGS_reg_43_17_inst : DFF_X1 port map( D => n12950, CK => CLK, Q => n16523, 
                           QN => n4864);
   REGS_reg_43_16_inst : DFF_X1 port map( D => n12949, CK => CLK, Q => n16522, 
                           QN => n4865);
   REGS_reg_43_15_inst : DFF_X1 port map( D => n12948, CK => CLK, Q => n16521, 
                           QN => n4866);
   REGS_reg_43_14_inst : DFF_X1 port map( D => n12947, CK => CLK, Q => n16520, 
                           QN => n4867);
   REGS_reg_43_13_inst : DFF_X1 port map( D => n12946, CK => CLK, Q => n16519, 
                           QN => n4868);
   REGS_reg_43_12_inst : DFF_X1 port map( D => n12945, CK => CLK, Q => n16518, 
                           QN => n4869);
   REGS_reg_43_11_inst : DFF_X1 port map( D => n12944, CK => CLK, Q => n16517, 
                           QN => n4870);
   REGS_reg_43_10_inst : DFF_X1 port map( D => n12943, CK => CLK, Q => n16516, 
                           QN => n4871);
   REGS_reg_43_9_inst : DFF_X1 port map( D => n12942, CK => CLK, Q => n16515, 
                           QN => n4872);
   REGS_reg_43_8_inst : DFF_X1 port map( D => n12941, CK => CLK, Q => n16514, 
                           QN => n4873);
   REGS_reg_43_7_inst : DFF_X1 port map( D => n12940, CK => CLK, Q => n16513, 
                           QN => n4874);
   REGS_reg_43_6_inst : DFF_X1 port map( D => n12939, CK => CLK, Q => n16512, 
                           QN => n4875);
   REGS_reg_43_5_inst : DFF_X1 port map( D => n12938, CK => CLK, Q => n16511, 
                           QN => n4876);
   REGS_reg_43_4_inst : DFF_X1 port map( D => n12937, CK => CLK, Q => n16510, 
                           QN => n4877);
   REGS_reg_43_3_inst : DFF_X1 port map( D => n12936, CK => CLK, Q => n16509, 
                           QN => n4878);
   REGS_reg_43_2_inst : DFF_X1 port map( D => n12935, CK => CLK, Q => n16508, 
                           QN => n4879);
   REGS_reg_43_1_inst : DFF_X1 port map( D => n12934, CK => CLK, Q => n16507, 
                           QN => n4880);
   REGS_reg_43_0_inst : DFF_X1 port map( D => n12933, CK => CLK, Q => n16506, 
                           QN => n4881);
   REGS_reg_42_23_inst : DFF_X1 port map( D => n12988, CK => CLK, Q => n16683, 
                           QN => n4882);
   REGS_reg_42_22_inst : DFF_X1 port map( D => n12987, CK => CLK, Q => n16682, 
                           QN => n4883);
   REGS_reg_42_21_inst : DFF_X1 port map( D => n12986, CK => CLK, Q => n16681, 
                           QN => n4884);
   REGS_reg_42_20_inst : DFF_X1 port map( D => n12985, CK => CLK, Q => n16680, 
                           QN => n4885);
   REGS_reg_42_19_inst : DFF_X1 port map( D => n12984, CK => CLK, Q => n16679, 
                           QN => n4886);
   REGS_reg_42_18_inst : DFF_X1 port map( D => n12983, CK => CLK, Q => n16678, 
                           QN => n4887);
   REGS_reg_42_17_inst : DFF_X1 port map( D => n12982, CK => CLK, Q => n16677, 
                           QN => n4888);
   REGS_reg_42_16_inst : DFF_X1 port map( D => n12981, CK => CLK, Q => n16676, 
                           QN => n4889);
   REGS_reg_42_15_inst : DFF_X1 port map( D => n12980, CK => CLK, Q => n16675, 
                           QN => n4890);
   REGS_reg_42_14_inst : DFF_X1 port map( D => n12979, CK => CLK, Q => n16674, 
                           QN => n4891);
   REGS_reg_42_13_inst : DFF_X1 port map( D => n12978, CK => CLK, Q => n16673, 
                           QN => n4892);
   REGS_reg_42_12_inst : DFF_X1 port map( D => n12977, CK => CLK, Q => n16672, 
                           QN => n4893);
   REGS_reg_42_11_inst : DFF_X1 port map( D => n12976, CK => CLK, Q => n16671, 
                           QN => n4894);
   REGS_reg_42_10_inst : DFF_X1 port map( D => n12975, CK => CLK, Q => n16670, 
                           QN => n4895);
   REGS_reg_42_9_inst : DFF_X1 port map( D => n12974, CK => CLK, Q => n16669, 
                           QN => n4896);
   REGS_reg_42_8_inst : DFF_X1 port map( D => n12973, CK => CLK, Q => n16668, 
                           QN => n4897);
   REGS_reg_42_7_inst : DFF_X1 port map( D => n12972, CK => CLK, Q => n16667, 
                           QN => n4898);
   REGS_reg_42_6_inst : DFF_X1 port map( D => n12971, CK => CLK, Q => n16666, 
                           QN => n4899);
   REGS_reg_42_5_inst : DFF_X1 port map( D => n12970, CK => CLK, Q => n16665, 
                           QN => n4900);
   REGS_reg_42_4_inst : DFF_X1 port map( D => n12969, CK => CLK, Q => n16664, 
                           QN => n4901);
   REGS_reg_42_3_inst : DFF_X1 port map( D => n12968, CK => CLK, Q => n16663, 
                           QN => n4902);
   REGS_reg_42_2_inst : DFF_X1 port map( D => n12967, CK => CLK, Q => n16662, 
                           QN => n4903);
   REGS_reg_42_1_inst : DFF_X1 port map( D => n12966, CK => CLK, Q => n16661, 
                           QN => n4904);
   REGS_reg_42_0_inst : DFF_X1 port map( D => n12965, CK => CLK, Q => n16660, 
                           QN => n4905);
   REGS_reg_41_23_inst : DFF_X1 port map( D => n13020, CK => CLK, Q => n_1624, 
                           QN => n3209);
   REGS_reg_41_22_inst : DFF_X1 port map( D => n13019, CK => CLK, Q => n_1625, 
                           QN => n3210);
   REGS_reg_41_21_inst : DFF_X1 port map( D => n13018, CK => CLK, Q => n_1626, 
                           QN => n3211);
   REGS_reg_41_20_inst : DFF_X1 port map( D => n13017, CK => CLK, Q => n_1627, 
                           QN => n3212);
   REGS_reg_41_19_inst : DFF_X1 port map( D => n13016, CK => CLK, Q => n_1628, 
                           QN => n3213);
   REGS_reg_41_18_inst : DFF_X1 port map( D => n13015, CK => CLK, Q => n_1629, 
                           QN => n3214);
   REGS_reg_41_17_inst : DFF_X1 port map( D => n13014, CK => CLK, Q => n_1630, 
                           QN => n3215);
   REGS_reg_41_16_inst : DFF_X1 port map( D => n13013, CK => CLK, Q => n_1631, 
                           QN => n3216);
   REGS_reg_41_15_inst : DFF_X1 port map( D => n13012, CK => CLK, Q => n_1632, 
                           QN => n3217);
   REGS_reg_41_14_inst : DFF_X1 port map( D => n13011, CK => CLK, Q => n_1633, 
                           QN => n3218);
   REGS_reg_41_13_inst : DFF_X1 port map( D => n13010, CK => CLK, Q => n_1634, 
                           QN => n3219);
   REGS_reg_41_12_inst : DFF_X1 port map( D => n13009, CK => CLK, Q => n_1635, 
                           QN => n3220);
   REGS_reg_41_11_inst : DFF_X1 port map( D => n13008, CK => CLK, Q => n_1636, 
                           QN => n3221);
   REGS_reg_41_10_inst : DFF_X1 port map( D => n13007, CK => CLK, Q => n_1637, 
                           QN => n3222);
   REGS_reg_41_9_inst : DFF_X1 port map( D => n13006, CK => CLK, Q => n_1638, 
                           QN => n3223);
   REGS_reg_41_8_inst : DFF_X1 port map( D => n13005, CK => CLK, Q => n_1639, 
                           QN => n3224);
   REGS_reg_41_7_inst : DFF_X1 port map( D => n13004, CK => CLK, Q => n_1640, 
                           QN => n3225);
   REGS_reg_41_6_inst : DFF_X1 port map( D => n13003, CK => CLK, Q => n_1641, 
                           QN => n3226);
   REGS_reg_41_5_inst : DFF_X1 port map( D => n13002, CK => CLK, Q => n_1642, 
                           QN => n3227);
   REGS_reg_41_4_inst : DFF_X1 port map( D => n13001, CK => CLK, Q => n_1643, 
                           QN => n3228);
   REGS_reg_41_3_inst : DFF_X1 port map( D => n13000, CK => CLK, Q => n_1644, 
                           QN => n3229);
   REGS_reg_41_2_inst : DFF_X1 port map( D => n12999, CK => CLK, Q => n_1645, 
                           QN => n3230);
   REGS_reg_41_1_inst : DFF_X1 port map( D => n12998, CK => CLK, Q => n_1646, 
                           QN => n3231);
   REGS_reg_41_0_inst : DFF_X1 port map( D => n12997, CK => CLK, Q => n_1647, 
                           QN => n3232);
   REGS_reg_40_23_inst : DFF_X1 port map( D => n13052, CK => CLK, Q => n_1648, 
                           QN => n3233);
   REGS_reg_40_22_inst : DFF_X1 port map( D => n13051, CK => CLK, Q => n_1649, 
                           QN => n3234);
   REGS_reg_40_21_inst : DFF_X1 port map( D => n13050, CK => CLK, Q => n_1650, 
                           QN => n3235);
   REGS_reg_40_20_inst : DFF_X1 port map( D => n13049, CK => CLK, Q => n_1651, 
                           QN => n3236);
   REGS_reg_40_19_inst : DFF_X1 port map( D => n13048, CK => CLK, Q => n_1652, 
                           QN => n3237);
   REGS_reg_40_18_inst : DFF_X1 port map( D => n13047, CK => CLK, Q => n_1653, 
                           QN => n3238);
   REGS_reg_40_17_inst : DFF_X1 port map( D => n13046, CK => CLK, Q => n_1654, 
                           QN => n3239);
   REGS_reg_40_16_inst : DFF_X1 port map( D => n13045, CK => CLK, Q => n_1655, 
                           QN => n3240);
   REGS_reg_40_15_inst : DFF_X1 port map( D => n13044, CK => CLK, Q => n_1656, 
                           QN => n3241);
   REGS_reg_40_14_inst : DFF_X1 port map( D => n13043, CK => CLK, Q => n_1657, 
                           QN => n3242);
   REGS_reg_40_13_inst : DFF_X1 port map( D => n13042, CK => CLK, Q => n_1658, 
                           QN => n3243);
   REGS_reg_40_12_inst : DFF_X1 port map( D => n13041, CK => CLK, Q => n_1659, 
                           QN => n3244);
   REGS_reg_40_11_inst : DFF_X1 port map( D => n13040, CK => CLK, Q => n_1660, 
                           QN => n3245);
   REGS_reg_40_10_inst : DFF_X1 port map( D => n13039, CK => CLK, Q => n_1661, 
                           QN => n3246);
   REGS_reg_40_9_inst : DFF_X1 port map( D => n13038, CK => CLK, Q => n_1662, 
                           QN => n3247);
   REGS_reg_40_8_inst : DFF_X1 port map( D => n13037, CK => CLK, Q => n_1663, 
                           QN => n3248);
   REGS_reg_40_7_inst : DFF_X1 port map( D => n13036, CK => CLK, Q => n_1664, 
                           QN => n3249);
   REGS_reg_40_6_inst : DFF_X1 port map( D => n13035, CK => CLK, Q => n_1665, 
                           QN => n3250);
   REGS_reg_40_5_inst : DFF_X1 port map( D => n13034, CK => CLK, Q => n_1666, 
                           QN => n3251);
   REGS_reg_40_4_inst : DFF_X1 port map( D => n13033, CK => CLK, Q => n_1667, 
                           QN => n3252);
   REGS_reg_40_3_inst : DFF_X1 port map( D => n13032, CK => CLK, Q => n_1668, 
                           QN => n3253);
   REGS_reg_40_2_inst : DFF_X1 port map( D => n13031, CK => CLK, Q => n_1669, 
                           QN => n3254);
   REGS_reg_40_1_inst : DFF_X1 port map( D => n13030, CK => CLK, Q => n_1670, 
                           QN => n3255);
   REGS_reg_40_0_inst : DFF_X1 port map( D => n13029, CK => CLK, Q => n_1671, 
                           QN => n3256);
   REGS_reg_35_23_inst : DFF_X1 port map( D => n13212, CK => CLK, Q => n16505, 
                           QN => n4954);
   REGS_reg_35_22_inst : DFF_X1 port map( D => n13211, CK => CLK, Q => n16504, 
                           QN => n4955);
   REGS_reg_35_21_inst : DFF_X1 port map( D => n13210, CK => CLK, Q => n16503, 
                           QN => n4956);
   REGS_reg_35_20_inst : DFF_X1 port map( D => n13209, CK => CLK, Q => n16502, 
                           QN => n4957);
   REGS_reg_35_19_inst : DFF_X1 port map( D => n13208, CK => CLK, Q => n16501, 
                           QN => n4958);
   REGS_reg_35_18_inst : DFF_X1 port map( D => n13207, CK => CLK, Q => n16500, 
                           QN => n4959);
   REGS_reg_35_17_inst : DFF_X1 port map( D => n13206, CK => CLK, Q => n16499, 
                           QN => n4960);
   REGS_reg_35_16_inst : DFF_X1 port map( D => n13205, CK => CLK, Q => n16498, 
                           QN => n4961);
   REGS_reg_35_15_inst : DFF_X1 port map( D => n13204, CK => CLK, Q => n16497, 
                           QN => n4962);
   REGS_reg_35_14_inst : DFF_X1 port map( D => n13203, CK => CLK, Q => n16496, 
                           QN => n4963);
   REGS_reg_35_13_inst : DFF_X1 port map( D => n13202, CK => CLK, Q => n16495, 
                           QN => n4964);
   REGS_reg_35_12_inst : DFF_X1 port map( D => n13201, CK => CLK, Q => n16494, 
                           QN => n4965);
   REGS_reg_35_11_inst : DFF_X1 port map( D => n13200, CK => CLK, Q => n16493, 
                           QN => n4966);
   REGS_reg_35_10_inst : DFF_X1 port map( D => n13199, CK => CLK, Q => n16492, 
                           QN => n4967);
   REGS_reg_35_9_inst : DFF_X1 port map( D => n13198, CK => CLK, Q => n16491, 
                           QN => n4968);
   REGS_reg_35_8_inst : DFF_X1 port map( D => n13197, CK => CLK, Q => n16490, 
                           QN => n4969);
   REGS_reg_35_7_inst : DFF_X1 port map( D => n13196, CK => CLK, Q => n16489, 
                           QN => n4970);
   REGS_reg_35_6_inst : DFF_X1 port map( D => n13195, CK => CLK, Q => n16488, 
                           QN => n4971);
   REGS_reg_35_5_inst : DFF_X1 port map( D => n13194, CK => CLK, Q => n16487, 
                           QN => n4972);
   REGS_reg_35_4_inst : DFF_X1 port map( D => n13193, CK => CLK, Q => n16486, 
                           QN => n4973);
   REGS_reg_35_3_inst : DFF_X1 port map( D => n13192, CK => CLK, Q => n16485, 
                           QN => n4974);
   REGS_reg_35_2_inst : DFF_X1 port map( D => n13191, CK => CLK, Q => n16484, 
                           QN => n4975);
   REGS_reg_35_1_inst : DFF_X1 port map( D => n13190, CK => CLK, Q => n16483, 
                           QN => n4976);
   REGS_reg_35_0_inst : DFF_X1 port map( D => n13189, CK => CLK, Q => n16482, 
                           QN => n4977);
   REGS_reg_34_23_inst : DFF_X1 port map( D => n13244, CK => CLK, Q => n16659, 
                           QN => n4978);
   REGS_reg_34_22_inst : DFF_X1 port map( D => n13243, CK => CLK, Q => n16658, 
                           QN => n4979);
   REGS_reg_34_21_inst : DFF_X1 port map( D => n13242, CK => CLK, Q => n16657, 
                           QN => n4980);
   REGS_reg_34_20_inst : DFF_X1 port map( D => n13241, CK => CLK, Q => n16656, 
                           QN => n4981);
   REGS_reg_34_19_inst : DFF_X1 port map( D => n13240, CK => CLK, Q => n16655, 
                           QN => n4982);
   REGS_reg_34_18_inst : DFF_X1 port map( D => n13239, CK => CLK, Q => n16654, 
                           QN => n4983);
   REGS_reg_34_17_inst : DFF_X1 port map( D => n13238, CK => CLK, Q => n16653, 
                           QN => n4984);
   REGS_reg_34_16_inst : DFF_X1 port map( D => n13237, CK => CLK, Q => n16652, 
                           QN => n4985);
   REGS_reg_34_15_inst : DFF_X1 port map( D => n13236, CK => CLK, Q => n16651, 
                           QN => n4986);
   REGS_reg_34_14_inst : DFF_X1 port map( D => n13235, CK => CLK, Q => n16650, 
                           QN => n4987);
   REGS_reg_34_13_inst : DFF_X1 port map( D => n13234, CK => CLK, Q => n16649, 
                           QN => n4988);
   REGS_reg_34_12_inst : DFF_X1 port map( D => n13233, CK => CLK, Q => n16648, 
                           QN => n4989);
   REGS_reg_34_11_inst : DFF_X1 port map( D => n13232, CK => CLK, Q => n16647, 
                           QN => n4990);
   REGS_reg_34_10_inst : DFF_X1 port map( D => n13231, CK => CLK, Q => n16646, 
                           QN => n4991);
   REGS_reg_34_9_inst : DFF_X1 port map( D => n13230, CK => CLK, Q => n16645, 
                           QN => n4992);
   REGS_reg_34_8_inst : DFF_X1 port map( D => n13229, CK => CLK, Q => n16644, 
                           QN => n4993);
   REGS_reg_34_7_inst : DFF_X1 port map( D => n13228, CK => CLK, Q => n16643, 
                           QN => n4994);
   REGS_reg_34_6_inst : DFF_X1 port map( D => n13227, CK => CLK, Q => n16642, 
                           QN => n4995);
   REGS_reg_34_5_inst : DFF_X1 port map( D => n13226, CK => CLK, Q => n16641, 
                           QN => n4996);
   REGS_reg_34_4_inst : DFF_X1 port map( D => n13225, CK => CLK, Q => n16640, 
                           QN => n4997);
   REGS_reg_34_3_inst : DFF_X1 port map( D => n13224, CK => CLK, Q => n16639, 
                           QN => n4998);
   REGS_reg_34_2_inst : DFF_X1 port map( D => n13223, CK => CLK, Q => n16638, 
                           QN => n4999);
   REGS_reg_34_1_inst : DFF_X1 port map( D => n13222, CK => CLK, Q => n16637, 
                           QN => n5000);
   REGS_reg_34_0_inst : DFF_X1 port map( D => n13221, CK => CLK, Q => n16636, 
                           QN => n5001);
   REGS_reg_13_23_inst : DFF_X1 port map( D => n13916, CK => CLK, Q => n16635, 
                           QN => n4504);
   REGS_reg_13_22_inst : DFF_X1 port map( D => n13915, CK => CLK, Q => n16634, 
                           QN => n4505);
   REGS_reg_13_21_inst : DFF_X1 port map( D => n13914, CK => CLK, Q => n16633, 
                           QN => n4506);
   REGS_reg_13_20_inst : DFF_X1 port map( D => n13913, CK => CLK, Q => n16632, 
                           QN => n4507);
   REGS_reg_13_19_inst : DFF_X1 port map( D => n13912, CK => CLK, Q => n16631, 
                           QN => n4508);
   REGS_reg_13_18_inst : DFF_X1 port map( D => n13911, CK => CLK, Q => n16630, 
                           QN => n4509);
   REGS_reg_13_17_inst : DFF_X1 port map( D => n13910, CK => CLK, Q => n16629, 
                           QN => n4510);
   REGS_reg_13_16_inst : DFF_X1 port map( D => n13909, CK => CLK, Q => n16628, 
                           QN => n4511);
   REGS_reg_13_15_inst : DFF_X1 port map( D => n13908, CK => CLK, Q => n16627, 
                           QN => n4512);
   REGS_reg_13_14_inst : DFF_X1 port map( D => n13907, CK => CLK, Q => n16626, 
                           QN => n4513);
   REGS_reg_13_13_inst : DFF_X1 port map( D => n13906, CK => CLK, Q => n16625, 
                           QN => n4514);
   REGS_reg_13_12_inst : DFF_X1 port map( D => n13905, CK => CLK, Q => n16624, 
                           QN => n4515);
   REGS_reg_13_11_inst : DFF_X1 port map( D => n13904, CK => CLK, Q => n16623, 
                           QN => n4516);
   REGS_reg_13_10_inst : DFF_X1 port map( D => n13903, CK => CLK, Q => n16622, 
                           QN => n4517);
   REGS_reg_13_9_inst : DFF_X1 port map( D => n13902, CK => CLK, Q => n16621, 
                           QN => n4518);
   REGS_reg_13_8_inst : DFF_X1 port map( D => n13901, CK => CLK, Q => n16620, 
                           QN => n4519);
   REGS_reg_13_7_inst : DFF_X1 port map( D => n13900, CK => CLK, Q => n16619, 
                           QN => n4520);
   REGS_reg_13_6_inst : DFF_X1 port map( D => n13899, CK => CLK, Q => n16618, 
                           QN => n4521);
   REGS_reg_13_5_inst : DFF_X1 port map( D => n13898, CK => CLK, Q => n16617, 
                           QN => n4522);
   REGS_reg_13_4_inst : DFF_X1 port map( D => n13897, CK => CLK, Q => n16616, 
                           QN => n4523);
   REGS_reg_13_3_inst : DFF_X1 port map( D => n13896, CK => CLK, Q => n16615, 
                           QN => n4524);
   REGS_reg_13_2_inst : DFF_X1 port map( D => n13895, CK => CLK, Q => n16614, 
                           QN => n4525);
   REGS_reg_13_1_inst : DFF_X1 port map( D => n13894, CK => CLK, Q => n16613, 
                           QN => n4526);
   REGS_reg_13_0_inst : DFF_X1 port map( D => n13893, CK => CLK, Q => n16612, 
                           QN => n4527);
   REGS_reg_12_23_inst : DFF_X1 port map( D => n13948, CK => CLK, Q => n16611, 
                           QN => n4528);
   REGS_reg_12_22_inst : DFF_X1 port map( D => n13947, CK => CLK, Q => n16610, 
                           QN => n4529);
   REGS_reg_12_21_inst : DFF_X1 port map( D => n13946, CK => CLK, Q => n16609, 
                           QN => n4530);
   REGS_reg_12_20_inst : DFF_X1 port map( D => n13945, CK => CLK, Q => n16608, 
                           QN => n4531);
   REGS_reg_12_19_inst : DFF_X1 port map( D => n13944, CK => CLK, Q => n16607, 
                           QN => n4532);
   REGS_reg_12_18_inst : DFF_X1 port map( D => n13943, CK => CLK, Q => n16606, 
                           QN => n4533);
   REGS_reg_12_17_inst : DFF_X1 port map( D => n13942, CK => CLK, Q => n16605, 
                           QN => n4534);
   REGS_reg_12_16_inst : DFF_X1 port map( D => n13941, CK => CLK, Q => n16604, 
                           QN => n4535);
   REGS_reg_12_15_inst : DFF_X1 port map( D => n13940, CK => CLK, Q => n16603, 
                           QN => n4536);
   REGS_reg_12_14_inst : DFF_X1 port map( D => n13939, CK => CLK, Q => n16602, 
                           QN => n4537);
   REGS_reg_12_13_inst : DFF_X1 port map( D => n13938, CK => CLK, Q => n16601, 
                           QN => n4538);
   REGS_reg_12_12_inst : DFF_X1 port map( D => n13937, CK => CLK, Q => n16600, 
                           QN => n4539);
   REGS_reg_12_11_inst : DFF_X1 port map( D => n13936, CK => CLK, Q => n16599, 
                           QN => n4540);
   REGS_reg_12_10_inst : DFF_X1 port map( D => n13935, CK => CLK, Q => n16598, 
                           QN => n4541);
   REGS_reg_12_9_inst : DFF_X1 port map( D => n13934, CK => CLK, Q => n16597, 
                           QN => n4542);
   REGS_reg_12_8_inst : DFF_X1 port map( D => n13933, CK => CLK, Q => n16596, 
                           QN => n4543);
   REGS_reg_12_7_inst : DFF_X1 port map( D => n13932, CK => CLK, Q => n16595, 
                           QN => n4544);
   REGS_reg_12_6_inst : DFF_X1 port map( D => n13931, CK => CLK, Q => n16594, 
                           QN => n4545);
   REGS_reg_12_5_inst : DFF_X1 port map( D => n13930, CK => CLK, Q => n16593, 
                           QN => n4546);
   REGS_reg_12_4_inst : DFF_X1 port map( D => n13929, CK => CLK, Q => n16592, 
                           QN => n4547);
   REGS_reg_12_3_inst : DFF_X1 port map( D => n13928, CK => CLK, Q => n16591, 
                           QN => n4548);
   REGS_reg_12_2_inst : DFF_X1 port map( D => n13927, CK => CLK, Q => n16590, 
                           QN => n4549);
   REGS_reg_12_1_inst : DFF_X1 port map( D => n13926, CK => CLK, Q => n16589, 
                           QN => n4550);
   REGS_reg_12_0_inst : DFF_X1 port map( D => n13925, CK => CLK, Q => n16588, 
                           QN => n4551);
   REGS_reg_10_23_inst : DFF_X1 port map( D => n14012, CK => CLK, Q => n53476, 
                           QN => n2725);
   REGS_reg_10_22_inst : DFF_X1 port map( D => n14011, CK => CLK, Q => n53477, 
                           QN => n2726);
   REGS_reg_10_21_inst : DFF_X1 port map( D => n14010, CK => CLK, Q => n53478, 
                           QN => n2727);
   REGS_reg_10_20_inst : DFF_X1 port map( D => n14009, CK => CLK, Q => n53479, 
                           QN => n2728);
   REGS_reg_10_19_inst : DFF_X1 port map( D => n14008, CK => CLK, Q => n53480, 
                           QN => n2729);
   REGS_reg_10_18_inst : DFF_X1 port map( D => n14007, CK => CLK, Q => n53481, 
                           QN => n2730);
   REGS_reg_10_17_inst : DFF_X1 port map( D => n14006, CK => CLK, Q => n53482, 
                           QN => n2731);
   REGS_reg_10_16_inst : DFF_X1 port map( D => n14005, CK => CLK, Q => n53483, 
                           QN => n2732);
   REGS_reg_10_15_inst : DFF_X1 port map( D => n14004, CK => CLK, Q => n53484, 
                           QN => n2733);
   REGS_reg_10_14_inst : DFF_X1 port map( D => n14003, CK => CLK, Q => n53485, 
                           QN => n2734);
   REGS_reg_10_13_inst : DFF_X1 port map( D => n14002, CK => CLK, Q => n53486, 
                           QN => n2735);
   REGS_reg_10_12_inst : DFF_X1 port map( D => n14001, CK => CLK, Q => n53487, 
                           QN => n2736);
   REGS_reg_10_11_inst : DFF_X1 port map( D => n14000, CK => CLK, Q => n53488, 
                           QN => n2737);
   REGS_reg_10_10_inst : DFF_X1 port map( D => n13999, CK => CLK, Q => n53489, 
                           QN => n2738);
   REGS_reg_10_9_inst : DFF_X1 port map( D => n13998, CK => CLK, Q => n53490, 
                           QN => n2739);
   REGS_reg_10_8_inst : DFF_X1 port map( D => n13997, CK => CLK, Q => n53491, 
                           QN => n2740);
   REGS_reg_10_7_inst : DFF_X1 port map( D => n13996, CK => CLK, Q => n53492, 
                           QN => n2741);
   REGS_reg_10_6_inst : DFF_X1 port map( D => n13995, CK => CLK, Q => n53493, 
                           QN => n2742);
   REGS_reg_10_5_inst : DFF_X1 port map( D => n13994, CK => CLK, Q => n53494, 
                           QN => n2743);
   REGS_reg_10_4_inst : DFF_X1 port map( D => n13993, CK => CLK, Q => n53495, 
                           QN => n2744);
   REGS_reg_10_3_inst : DFF_X1 port map( D => n13992, CK => CLK, Q => n53496, 
                           QN => n2745);
   REGS_reg_10_2_inst : DFF_X1 port map( D => n13991, CK => CLK, Q => n53497, 
                           QN => n2746);
   REGS_reg_10_1_inst : DFF_X1 port map( D => n13990, CK => CLK, Q => n53498, 
                           QN => n2747);
   REGS_reg_10_0_inst : DFF_X1 port map( D => n13989, CK => CLK, Q => n53499, 
                           QN => n2748);
   REGS_reg_9_23_inst : DFF_X1 port map( D => n14044, CK => CLK, Q => n_1672, 
                           QN => n4576);
   REGS_reg_9_22_inst : DFF_X1 port map( D => n14043, CK => CLK, Q => n_1673, 
                           QN => n4577);
   REGS_reg_9_21_inst : DFF_X1 port map( D => n14042, CK => CLK, Q => n_1674, 
                           QN => n4578);
   REGS_reg_9_20_inst : DFF_X1 port map( D => n14041, CK => CLK, Q => n_1675, 
                           QN => n4579);
   REGS_reg_9_19_inst : DFF_X1 port map( D => n14040, CK => CLK, Q => n_1676, 
                           QN => n4580);
   REGS_reg_9_18_inst : DFF_X1 port map( D => n14039, CK => CLK, Q => n_1677, 
                           QN => n4581);
   REGS_reg_9_17_inst : DFF_X1 port map( D => n14038, CK => CLK, Q => n_1678, 
                           QN => n4582);
   REGS_reg_9_16_inst : DFF_X1 port map( D => n14037, CK => CLK, Q => n_1679, 
                           QN => n4583);
   REGS_reg_9_15_inst : DFF_X1 port map( D => n14036, CK => CLK, Q => n_1680, 
                           QN => n4584);
   REGS_reg_9_14_inst : DFF_X1 port map( D => n14035, CK => CLK, Q => n_1681, 
                           QN => n4585);
   REGS_reg_9_13_inst : DFF_X1 port map( D => n14034, CK => CLK, Q => n_1682, 
                           QN => n4586);
   REGS_reg_9_12_inst : DFF_X1 port map( D => n14033, CK => CLK, Q => n_1683, 
                           QN => n4587);
   REGS_reg_9_11_inst : DFF_X1 port map( D => n14032, CK => CLK, Q => n_1684, 
                           QN => n4588);
   REGS_reg_9_10_inst : DFF_X1 port map( D => n14031, CK => CLK, Q => n_1685, 
                           QN => n4589);
   REGS_reg_9_9_inst : DFF_X1 port map( D => n14030, CK => CLK, Q => n_1686, QN
                           => n4590);
   REGS_reg_9_8_inst : DFF_X1 port map( D => n14029, CK => CLK, Q => n_1687, QN
                           => n4591);
   REGS_reg_9_7_inst : DFF_X1 port map( D => n14028, CK => CLK, Q => n_1688, QN
                           => n4592);
   REGS_reg_9_6_inst : DFF_X1 port map( D => n14027, CK => CLK, Q => n_1689, QN
                           => n4593);
   REGS_reg_9_5_inst : DFF_X1 port map( D => n14026, CK => CLK, Q => n_1690, QN
                           => n4594);
   REGS_reg_9_4_inst : DFF_X1 port map( D => n14025, CK => CLK, Q => n_1691, QN
                           => n4595);
   REGS_reg_9_3_inst : DFF_X1 port map( D => n14024, CK => CLK, Q => n_1692, QN
                           => n4596);
   REGS_reg_9_2_inst : DFF_X1 port map( D => n14023, CK => CLK, Q => n_1693, QN
                           => n4597);
   REGS_reg_9_1_inst : DFF_X1 port map( D => n14022, CK => CLK, Q => n_1694, QN
                           => n4598);
   REGS_reg_9_0_inst : DFF_X1 port map( D => n14021, CK => CLK, Q => n_1695, QN
                           => n4599);
   REGS_reg_8_23_inst : DFF_X1 port map( D => n14076, CK => CLK, Q => n16798, 
                           QN => n4600);
   REGS_reg_8_22_inst : DFF_X1 port map( D => n14075, CK => CLK, Q => n16797, 
                           QN => n4601);
   REGS_reg_8_21_inst : DFF_X1 port map( D => n14074, CK => CLK, Q => n16796, 
                           QN => n4602);
   REGS_reg_8_20_inst : DFF_X1 port map( D => n14073, CK => CLK, Q => n16795, 
                           QN => n4603);
   REGS_reg_8_19_inst : DFF_X1 port map( D => n14072, CK => CLK, Q => n16806, 
                           QN => n4604);
   REGS_reg_8_18_inst : DFF_X1 port map( D => n14071, CK => CLK, Q => n16805, 
                           QN => n4605);
   REGS_reg_8_17_inst : DFF_X1 port map( D => n14070, CK => CLK, Q => n16804, 
                           QN => n4606);
   REGS_reg_8_16_inst : DFF_X1 port map( D => n14069, CK => CLK, Q => n16803, 
                           QN => n4607);
   REGS_reg_8_15_inst : DFF_X1 port map( D => n14068, CK => CLK, Q => n16802, 
                           QN => n4608);
   REGS_reg_8_14_inst : DFF_X1 port map( D => n14067, CK => CLK, Q => n16810, 
                           QN => n4609);
   REGS_reg_8_13_inst : DFF_X1 port map( D => n14066, CK => CLK, Q => n16809, 
                           QN => n4610);
   REGS_reg_8_12_inst : DFF_X1 port map( D => n14065, CK => CLK, Q => n16801, 
                           QN => n4611);
   REGS_reg_8_11_inst : DFF_X1 port map( D => n14064, CK => CLK, Q => n16808, 
                           QN => n4612);
   REGS_reg_8_10_inst : DFF_X1 port map( D => n14063, CK => CLK, Q => n16807, 
                           QN => n4613);
   REGS_reg_8_9_inst : DFF_X1 port map( D => n14062, CK => CLK, Q => n16800, QN
                           => n4614);
   REGS_reg_8_8_inst : DFF_X1 port map( D => n14061, CK => CLK, Q => n16794, QN
                           => n4615);
   REGS_reg_8_7_inst : DFF_X1 port map( D => n14060, CK => CLK, Q => n16799, QN
                           => n4616);
   REGS_reg_8_6_inst : DFF_X1 port map( D => n14059, CK => CLK, Q => n16793, QN
                           => n4617);
   REGS_reg_8_5_inst : DFF_X1 port map( D => n14058, CK => CLK, Q => n16792, QN
                           => n4618);
   REGS_reg_8_4_inst : DFF_X1 port map( D => n14057, CK => CLK, Q => n16791, QN
                           => n4619);
   REGS_reg_8_3_inst : DFF_X1 port map( D => n14056, CK => CLK, Q => n16790, QN
                           => n4620);
   REGS_reg_8_2_inst : DFF_X1 port map( D => n14055, CK => CLK, Q => n16813, QN
                           => n4621);
   REGS_reg_8_1_inst : DFF_X1 port map( D => n14054, CK => CLK, Q => n16812, QN
                           => n4622);
   REGS_reg_8_0_inst : DFF_X1 port map( D => n14053, CK => CLK, Q => n16811, QN
                           => n4623);
   REGS_reg_5_23_inst : DFF_X1 port map( D => n14172, CK => CLK, Q => n_1696, 
                           QN => n4648);
   REGS_reg_5_22_inst : DFF_X1 port map( D => n14171, CK => CLK, Q => n_1697, 
                           QN => n4649);
   REGS_reg_5_21_inst : DFF_X1 port map( D => n14170, CK => CLK, Q => n_1698, 
                           QN => n4650);
   REGS_reg_5_20_inst : DFF_X1 port map( D => n14169, CK => CLK, Q => n_1699, 
                           QN => n4651);
   REGS_reg_5_19_inst : DFF_X1 port map( D => n14168, CK => CLK, Q => n_1700, 
                           QN => n4652);
   REGS_reg_5_18_inst : DFF_X1 port map( D => n14167, CK => CLK, Q => n_1701, 
                           QN => n4653);
   REGS_reg_5_17_inst : DFF_X1 port map( D => n14166, CK => CLK, Q => n_1702, 
                           QN => n4654);
   REGS_reg_5_16_inst : DFF_X1 port map( D => n14165, CK => CLK, Q => n_1703, 
                           QN => n4655);
   REGS_reg_5_15_inst : DFF_X1 port map( D => n14164, CK => CLK, Q => n_1704, 
                           QN => n4656);
   REGS_reg_5_14_inst : DFF_X1 port map( D => n14163, CK => CLK, Q => n_1705, 
                           QN => n4657);
   REGS_reg_5_13_inst : DFF_X1 port map( D => n14162, CK => CLK, Q => n_1706, 
                           QN => n4658);
   REGS_reg_5_12_inst : DFF_X1 port map( D => n14161, CK => CLK, Q => n_1707, 
                           QN => n4659);
   REGS_reg_5_11_inst : DFF_X1 port map( D => n14160, CK => CLK, Q => n_1708, 
                           QN => n4660);
   REGS_reg_5_10_inst : DFF_X1 port map( D => n14159, CK => CLK, Q => n_1709, 
                           QN => n4661);
   REGS_reg_5_9_inst : DFF_X1 port map( D => n14158, CK => CLK, Q => n_1710, QN
                           => n4662);
   REGS_reg_5_8_inst : DFF_X1 port map( D => n14157, CK => CLK, Q => n_1711, QN
                           => n4663);
   REGS_reg_5_7_inst : DFF_X1 port map( D => n14156, CK => CLK, Q => n_1712, QN
                           => n4664);
   REGS_reg_5_6_inst : DFF_X1 port map( D => n14155, CK => CLK, Q => n_1713, QN
                           => n4665);
   REGS_reg_5_5_inst : DFF_X1 port map( D => n14154, CK => CLK, Q => n_1714, QN
                           => n4666);
   REGS_reg_5_4_inst : DFF_X1 port map( D => n14153, CK => CLK, Q => n_1715, QN
                           => n4667);
   REGS_reg_5_3_inst : DFF_X1 port map( D => n14152, CK => CLK, Q => n_1716, QN
                           => n4668);
   REGS_reg_5_2_inst : DFF_X1 port map( D => n14151, CK => CLK, Q => n_1717, QN
                           => n4669);
   REGS_reg_5_1_inst : DFF_X1 port map( D => n14150, CK => CLK, Q => n_1718, QN
                           => n4670);
   REGS_reg_5_0_inst : DFF_X1 port map( D => n14149, CK => CLK, Q => n_1719, QN
                           => n4671);
   REGS_reg_4_23_inst : DFF_X1 port map( D => n14204, CK => CLK, Q => n_1720, 
                           QN => n4672);
   REGS_reg_4_22_inst : DFF_X1 port map( D => n14203, CK => CLK, Q => n_1721, 
                           QN => n4673);
   REGS_reg_4_21_inst : DFF_X1 port map( D => n14202, CK => CLK, Q => n_1722, 
                           QN => n4674);
   REGS_reg_4_20_inst : DFF_X1 port map( D => n14201, CK => CLK, Q => n_1723, 
                           QN => n4675);
   REGS_reg_4_19_inst : DFF_X1 port map( D => n14200, CK => CLK, Q => n_1724, 
                           QN => n4676);
   REGS_reg_4_18_inst : DFF_X1 port map( D => n14199, CK => CLK, Q => n_1725, 
                           QN => n4677);
   REGS_reg_4_17_inst : DFF_X1 port map( D => n14198, CK => CLK, Q => n_1726, 
                           QN => n4678);
   REGS_reg_4_16_inst : DFF_X1 port map( D => n14197, CK => CLK, Q => n_1727, 
                           QN => n4679);
   REGS_reg_4_15_inst : DFF_X1 port map( D => n14196, CK => CLK, Q => n_1728, 
                           QN => n4680);
   REGS_reg_4_14_inst : DFF_X1 port map( D => n14195, CK => CLK, Q => n_1729, 
                           QN => n4681);
   REGS_reg_4_13_inst : DFF_X1 port map( D => n14194, CK => CLK, Q => n_1730, 
                           QN => n4682);
   REGS_reg_4_12_inst : DFF_X1 port map( D => n14193, CK => CLK, Q => n_1731, 
                           QN => n4683);
   REGS_reg_4_11_inst : DFF_X1 port map( D => n14192, CK => CLK, Q => n_1732, 
                           QN => n4684);
   REGS_reg_4_10_inst : DFF_X1 port map( D => n14191, CK => CLK, Q => n_1733, 
                           QN => n4685);
   REGS_reg_4_9_inst : DFF_X1 port map( D => n14190, CK => CLK, Q => n_1734, QN
                           => n4686);
   REGS_reg_4_8_inst : DFF_X1 port map( D => n14189, CK => CLK, Q => n_1735, QN
                           => n4687);
   REGS_reg_4_7_inst : DFF_X1 port map( D => n14188, CK => CLK, Q => n_1736, QN
                           => n4688);
   REGS_reg_4_6_inst : DFF_X1 port map( D => n14187, CK => CLK, Q => n_1737, QN
                           => n4689);
   REGS_reg_4_5_inst : DFF_X1 port map( D => n14186, CK => CLK, Q => n_1738, QN
                           => n4690);
   REGS_reg_4_4_inst : DFF_X1 port map( D => n14185, CK => CLK, Q => n_1739, QN
                           => n4691);
   REGS_reg_4_3_inst : DFF_X1 port map( D => n14184, CK => CLK, Q => n_1740, QN
                           => n4692);
   REGS_reg_4_2_inst : DFF_X1 port map( D => n14183, CK => CLK, Q => n_1741, QN
                           => n4693);
   REGS_reg_4_1_inst : DFF_X1 port map( D => n14182, CK => CLK, Q => n_1742, QN
                           => n4694);
   REGS_reg_4_0_inst : DFF_X1 port map( D => n14181, CK => CLK, Q => n_1743, QN
                           => n4695);
   REGS_reg_3_23_inst : DFF_X1 port map( D => n14236, CK => CLK, Q => n936, QN 
                           => n2749);
   REGS_reg_3_22_inst : DFF_X1 port map( D => n14235, CK => CLK, Q => n937, QN 
                           => n2750);
   REGS_reg_3_21_inst : DFF_X1 port map( D => n14234, CK => CLK, Q => n938, QN 
                           => n2751);
   REGS_reg_3_20_inst : DFF_X1 port map( D => n14233, CK => CLK, Q => n939, QN 
                           => n2752);
   REGS_reg_3_19_inst : DFF_X1 port map( D => n14232, CK => CLK, Q => n940, QN 
                           => n2753);
   REGS_reg_3_18_inst : DFF_X1 port map( D => n14231, CK => CLK, Q => n941, QN 
                           => n2754);
   REGS_reg_3_17_inst : DFF_X1 port map( D => n14230, CK => CLK, Q => n942, QN 
                           => n2755);
   REGS_reg_3_16_inst : DFF_X1 port map( D => n14229, CK => CLK, Q => n943, QN 
                           => n2756);
   REGS_reg_3_15_inst : DFF_X1 port map( D => n14228, CK => CLK, Q => n944, QN 
                           => n2757);
   REGS_reg_3_14_inst : DFF_X1 port map( D => n14227, CK => CLK, Q => n945, QN 
                           => n2758);
   REGS_reg_3_13_inst : DFF_X1 port map( D => n14226, CK => CLK, Q => n946, QN 
                           => n2759);
   REGS_reg_3_12_inst : DFF_X1 port map( D => n14225, CK => CLK, Q => n947, QN 
                           => n2760);
   REGS_reg_3_11_inst : DFF_X1 port map( D => n14224, CK => CLK, Q => n948, QN 
                           => n2761);
   REGS_reg_3_10_inst : DFF_X1 port map( D => n14223, CK => CLK, Q => n949, QN 
                           => n2762);
   REGS_reg_3_9_inst : DFF_X1 port map( D => n14222, CK => CLK, Q => n950, QN 
                           => n2763);
   REGS_reg_3_8_inst : DFF_X1 port map( D => n14221, CK => CLK, Q => n951, QN 
                           => n2764);
   REGS_reg_3_7_inst : DFF_X1 port map( D => n14220, CK => CLK, Q => n952, QN 
                           => n2765);
   REGS_reg_3_6_inst : DFF_X1 port map( D => n14219, CK => CLK, Q => n953, QN 
                           => n2766);
   REGS_reg_3_5_inst : DFF_X1 port map( D => n14218, CK => CLK, Q => n954, QN 
                           => n2767);
   REGS_reg_3_4_inst : DFF_X1 port map( D => n14217, CK => CLK, Q => n955, QN 
                           => n2768);
   REGS_reg_3_3_inst : DFF_X1 port map( D => n14216, CK => CLK, Q => n956, QN 
                           => n2769);
   REGS_reg_2_8_inst : DFF_X1 port map( D => n14253, CK => CLK, Q => n963, QN 
                           => n2770);
   REGS_reg_2_7_inst : DFF_X1 port map( D => n14252, CK => CLK, Q => n964, QN 
                           => n2771);
   REGS_reg_2_6_inst : DFF_X1 port map( D => n14251, CK => CLK, Q => n965, QN 
                           => n2772);
   REGS_reg_2_5_inst : DFF_X1 port map( D => n14250, CK => CLK, Q => n966, QN 
                           => n2773);
   REGS_reg_2_4_inst : DFF_X1 port map( D => n14249, CK => CLK, Q => n967, QN 
                           => n2774);
   REGS_reg_2_3_inst : DFF_X1 port map( D => n14248, CK => CLK, Q => n968, QN 
                           => n2775);
   REGS_reg_2_2_inst : DFF_X1 port map( D => n14247, CK => CLK, Q => n969, QN 
                           => n2776);
   REGS_reg_2_1_inst : DFF_X1 port map( D => n14246, CK => CLK, Q => n970, QN 
                           => n2777);
   REGS_reg_2_0_inst : DFF_X1 port map( D => n14245, CK => CLK, Q => n971, QN 
                           => n2778);
   REGS_reg_127_23_inst : DFF_X1 port map( D => n10268, CK => CLK, Q => n15463,
                           QN => n3257);
   REGS_reg_127_22_inst : DFF_X1 port map( D => n10267, CK => CLK, Q => n15462,
                           QN => n3258);
   REGS_reg_127_21_inst : DFF_X1 port map( D => n10266, CK => CLK, Q => n15461,
                           QN => n3259);
   REGS_reg_127_20_inst : DFF_X1 port map( D => n10265, CK => CLK, Q => n15460,
                           QN => n3260);
   REGS_reg_127_19_inst : DFF_X1 port map( D => n10264, CK => CLK, Q => n15459,
                           QN => n3261);
   REGS_reg_127_18_inst : DFF_X1 port map( D => n10263, CK => CLK, Q => n15458,
                           QN => n3262);
   REGS_reg_127_17_inst : DFF_X1 port map( D => n10262, CK => CLK, Q => n15457,
                           QN => n3263);
   REGS_reg_127_16_inst : DFF_X1 port map( D => n10261, CK => CLK, Q => n15456,
                           QN => n3264);
   REGS_reg_127_15_inst : DFF_X1 port map( D => n10260, CK => CLK, Q => n15455,
                           QN => n3265);
   REGS_reg_127_14_inst : DFF_X1 port map( D => n10259, CK => CLK, Q => n15454,
                           QN => n3266);
   REGS_reg_127_13_inst : DFF_X1 port map( D => n10258, CK => CLK, Q => n15453,
                           QN => n3267);
   REGS_reg_127_12_inst : DFF_X1 port map( D => n10257, CK => CLK, Q => n15452,
                           QN => n3268);
   REGS_reg_127_11_inst : DFF_X1 port map( D => n10256, CK => CLK, Q => n15451,
                           QN => n3269);
   REGS_reg_127_10_inst : DFF_X1 port map( D => n10255, CK => CLK, Q => n15450,
                           QN => n3270);
   REGS_reg_127_9_inst : DFF_X1 port map( D => n10254, CK => CLK, Q => n15449, 
                           QN => n3271);
   REGS_reg_127_8_inst : DFF_X1 port map( D => n10253, CK => CLK, Q => n15448, 
                           QN => n3272);
   REGS_reg_127_7_inst : DFF_X1 port map( D => n10252, CK => CLK, Q => n15447, 
                           QN => n3273);
   REGS_reg_127_6_inst : DFF_X1 port map( D => n10251, CK => CLK, Q => n15446, 
                           QN => n3274);
   REGS_reg_127_5_inst : DFF_X1 port map( D => n10250, CK => CLK, Q => n15445, 
                           QN => n3275);
   REGS_reg_127_4_inst : DFF_X1 port map( D => n10249, CK => CLK, Q => n15444, 
                           QN => n3276);
   REGS_reg_127_3_inst : DFF_X1 port map( D => n10248, CK => CLK, Q => n15443, 
                           QN => n3277);
   REGS_reg_127_2_inst : DFF_X1 port map( D => n10247, CK => CLK, Q => n15442, 
                           QN => n3278);
   REGS_reg_127_1_inst : DFF_X1 port map( D => n10246, CK => CLK, Q => n15441, 
                           QN => n3279);
   REGS_reg_127_0_inst : DFF_X1 port map( D => n10245, CK => CLK, Q => n15440, 
                           QN => n3280);
   REGS_reg_126_23_inst : DFF_X1 port map( D => n10300, CK => CLK, Q => n996, 
                           QN => n3281);
   REGS_reg_126_22_inst : DFF_X1 port map( D => n10299, CK => CLK, Q => n997, 
                           QN => n3282);
   REGS_reg_126_21_inst : DFF_X1 port map( D => n10298, CK => CLK, Q => n998, 
                           QN => n3283);
   REGS_reg_126_20_inst : DFF_X1 port map( D => n10297, CK => CLK, Q => n999, 
                           QN => n3284);
   REGS_reg_126_19_inst : DFF_X1 port map( D => n10296, CK => CLK, Q => n2299, 
                           QN => n5050);
   REGS_reg_126_18_inst : DFF_X1 port map( D => n10295, CK => CLK, Q => n2300, 
                           QN => n5051);
   REGS_reg_126_17_inst : DFF_X1 port map( D => n10294, CK => CLK, Q => n2301, 
                           QN => n5052);
   REGS_reg_126_16_inst : DFF_X1 port map( D => n10293, CK => CLK, Q => n2302, 
                           QN => n5053);
   REGS_reg_126_15_inst : DFF_X1 port map( D => n10292, CK => CLK, Q => n2303, 
                           QN => n5054);
   REGS_reg_126_14_inst : DFF_X1 port map( D => n10291, CK => CLK, Q => n2304, 
                           QN => n5055);
   REGS_reg_126_13_inst : DFF_X1 port map( D => n10290, CK => CLK, Q => n2305, 
                           QN => n5056);
   REGS_reg_126_12_inst : DFF_X1 port map( D => n10289, CK => CLK, Q => n2306, 
                           QN => n5057);
   REGS_reg_126_11_inst : DFF_X1 port map( D => n10288, CK => CLK, Q => n2307, 
                           QN => n5058);
   REGS_reg_126_10_inst : DFF_X1 port map( D => n10287, CK => CLK, Q => n2308, 
                           QN => n5059);
   REGS_reg_126_9_inst : DFF_X1 port map( D => n10286, CK => CLK, Q => n2309, 
                           QN => n5060);
   REGS_reg_126_8_inst : DFF_X1 port map( D => n10285, CK => CLK, Q => n2310, 
                           QN => n5061);
   REGS_reg_126_7_inst : DFF_X1 port map( D => n10284, CK => CLK, Q => n2311, 
                           QN => n5062);
   REGS_reg_126_6_inst : DFF_X1 port map( D => n10283, CK => CLK, Q => n2312, 
                           QN => n5063);
   REGS_reg_126_5_inst : DFF_X1 port map( D => n10282, CK => CLK, Q => n2313, 
                           QN => n5064);
   REGS_reg_126_4_inst : DFF_X1 port map( D => n10281, CK => CLK, Q => n2314, 
                           QN => n5065);
   REGS_reg_126_3_inst : DFF_X1 port map( D => n10280, CK => CLK, Q => n2315, 
                           QN => n5066);
   REGS_reg_126_2_inst : DFF_X1 port map( D => n10279, CK => CLK, Q => n2316, 
                           QN => n5067);
   REGS_reg_126_1_inst : DFF_X1 port map( D => n10278, CK => CLK, Q => n2317, 
                           QN => n5068);
   REGS_reg_126_0_inst : DFF_X1 port map( D => n10277, CK => CLK, Q => n2318, 
                           QN => n5069);
   REGS_reg_125_23_inst : DFF_X1 port map( D => n10332, CK => CLK, Q => n2319, 
                           QN => n5070);
   REGS_reg_125_22_inst : DFF_X1 port map( D => n10331, CK => CLK, Q => n2320, 
                           QN => n5071);
   REGS_reg_125_21_inst : DFF_X1 port map( D => n10330, CK => CLK, Q => n2321, 
                           QN => n5072);
   REGS_reg_125_20_inst : DFF_X1 port map( D => n10329, CK => CLK, Q => n2322, 
                           QN => n5073);
   REGS_reg_125_19_inst : DFF_X1 port map( D => n10328, CK => CLK, Q => n2323, 
                           QN => n5074);
   REGS_reg_125_18_inst : DFF_X1 port map( D => n10327, CK => CLK, Q => n2324, 
                           QN => n5075);
   REGS_reg_125_17_inst : DFF_X1 port map( D => n10326, CK => CLK, Q => n2325, 
                           QN => n5076);
   REGS_reg_125_16_inst : DFF_X1 port map( D => n10325, CK => CLK, Q => n2326, 
                           QN => n5077);
   REGS_reg_125_15_inst : DFF_X1 port map( D => n10324, CK => CLK, Q => n2327, 
                           QN => n5078);
   REGS_reg_125_14_inst : DFF_X1 port map( D => n10323, CK => CLK, Q => n2328, 
                           QN => n5079);
   REGS_reg_125_13_inst : DFF_X1 port map( D => n10322, CK => CLK, Q => n2329, 
                           QN => n5080);
   REGS_reg_125_12_inst : DFF_X1 port map( D => n10321, CK => CLK, Q => n2330, 
                           QN => n5081);
   REGS_reg_125_11_inst : DFF_X1 port map( D => n10320, CK => CLK, Q => n2331, 
                           QN => n5082);
   REGS_reg_125_10_inst : DFF_X1 port map( D => n10319, CK => CLK, Q => n2332, 
                           QN => n5083);
   REGS_reg_125_9_inst : DFF_X1 port map( D => n10318, CK => CLK, Q => n2333, 
                           QN => n5084);
   REGS_reg_125_8_inst : DFF_X1 port map( D => n10317, CK => CLK, Q => n2334, 
                           QN => n5085);
   REGS_reg_125_7_inst : DFF_X1 port map( D => n10316, CK => CLK, Q => n2335, 
                           QN => n5086);
   REGS_reg_125_6_inst : DFF_X1 port map( D => n10315, CK => CLK, Q => n2336, 
                           QN => n5087);
   REGS_reg_125_5_inst : DFF_X1 port map( D => n10314, CK => CLK, Q => n2337, 
                           QN => n5088);
   REGS_reg_125_4_inst : DFF_X1 port map( D => n10313, CK => CLK, Q => n2338, 
                           QN => n5089);
   REGS_reg_125_3_inst : DFF_X1 port map( D => n10312, CK => CLK, Q => n2339, 
                           QN => n5090);
   REGS_reg_125_2_inst : DFF_X1 port map( D => n10311, CK => CLK, Q => n2340, 
                           QN => n5091);
   REGS_reg_125_1_inst : DFF_X1 port map( D => n10310, CK => CLK, Q => n2341, 
                           QN => n5092);
   REGS_reg_125_0_inst : DFF_X1 port map( D => n10309, CK => CLK, Q => n2342, 
                           QN => n5093);
   REGS_reg_124_23_inst : DFF_X1 port map( D => n10364, CK => CLK, Q => n52160,
                           QN => n3285);
   REGS_reg_124_22_inst : DFF_X1 port map( D => n10363, CK => CLK, Q => n52161,
                           QN => n3286);
   REGS_reg_124_21_inst : DFF_X1 port map( D => n10362, CK => CLK, Q => n52162,
                           QN => n3287);
   REGS_reg_124_20_inst : DFF_X1 port map( D => n10361, CK => CLK, Q => n52163,
                           QN => n3288);
   REGS_reg_124_19_inst : DFF_X1 port map( D => n10360, CK => CLK, Q => n52164,
                           QN => n3289);
   REGS_reg_124_18_inst : DFF_X1 port map( D => n10359, CK => CLK, Q => n52165,
                           QN => n3290);
   REGS_reg_124_17_inst : DFF_X1 port map( D => n10358, CK => CLK, Q => n52166,
                           QN => n3291);
   REGS_reg_124_16_inst : DFF_X1 port map( D => n10357, CK => CLK, Q => n52167,
                           QN => n3292);
   REGS_reg_124_15_inst : DFF_X1 port map( D => n10356, CK => CLK, Q => n52168,
                           QN => n3293);
   REGS_reg_124_14_inst : DFF_X1 port map( D => n10355, CK => CLK, Q => n52169,
                           QN => n3294);
   REGS_reg_124_13_inst : DFF_X1 port map( D => n10354, CK => CLK, Q => n52170,
                           QN => n3295);
   REGS_reg_124_12_inst : DFF_X1 port map( D => n10353, CK => CLK, Q => n52171,
                           QN => n3296);
   REGS_reg_124_11_inst : DFF_X1 port map( D => n10352, CK => CLK, Q => n52172,
                           QN => n3297);
   REGS_reg_124_10_inst : DFF_X1 port map( D => n10351, CK => CLK, Q => n52173,
                           QN => n3298);
   REGS_reg_124_9_inst : DFF_X1 port map( D => n10350, CK => CLK, Q => n52174, 
                           QN => n3299);
   REGS_reg_124_8_inst : DFF_X1 port map( D => n10349, CK => CLK, Q => n52175, 
                           QN => n3300);
   REGS_reg_124_7_inst : DFF_X1 port map( D => n10348, CK => CLK, Q => n52176, 
                           QN => n3301);
   REGS_reg_124_6_inst : DFF_X1 port map( D => n10347, CK => CLK, Q => n52177, 
                           QN => n3302);
   REGS_reg_124_5_inst : DFF_X1 port map( D => n10346, CK => CLK, Q => n52178, 
                           QN => n3303);
   REGS_reg_124_4_inst : DFF_X1 port map( D => n10345, CK => CLK, Q => n52179, 
                           QN => n3304);
   REGS_reg_124_3_inst : DFF_X1 port map( D => n10344, CK => CLK, Q => n52180, 
                           QN => n3305);
   REGS_reg_124_2_inst : DFF_X1 port map( D => n10343, CK => CLK, Q => n52181, 
                           QN => n3306);
   REGS_reg_124_1_inst : DFF_X1 port map( D => n10342, CK => CLK, Q => n52182, 
                           QN => n3307);
   REGS_reg_124_0_inst : DFF_X1 port map( D => n10341, CK => CLK, Q => n52183, 
                           QN => n3308);
   REGS_reg_123_23_inst : DFF_X1 port map( D => n10396, CK => CLK, Q => n52184,
                           QN => n3309);
   REGS_reg_123_22_inst : DFF_X1 port map( D => n10395, CK => CLK, Q => n52185,
                           QN => n3310);
   REGS_reg_123_21_inst : DFF_X1 port map( D => n10394, CK => CLK, Q => n52186,
                           QN => n3311);
   REGS_reg_123_20_inst : DFF_X1 port map( D => n10393, CK => CLK, Q => n52187,
                           QN => n3312);
   REGS_reg_123_19_inst : DFF_X1 port map( D => n10392, CK => CLK, Q => n52188,
                           QN => n3313);
   REGS_reg_123_18_inst : DFF_X1 port map( D => n10391, CK => CLK, Q => n52189,
                           QN => n3314);
   REGS_reg_123_17_inst : DFF_X1 port map( D => n10390, CK => CLK, Q => n52190,
                           QN => n3315);
   REGS_reg_123_16_inst : DFF_X1 port map( D => n10389, CK => CLK, Q => n52191,
                           QN => n3316);
   REGS_reg_123_15_inst : DFF_X1 port map( D => n10388, CK => CLK, Q => n52192,
                           QN => n3317);
   REGS_reg_123_14_inst : DFF_X1 port map( D => n10387, CK => CLK, Q => n52193,
                           QN => n3318);
   REGS_reg_123_13_inst : DFF_X1 port map( D => n10386, CK => CLK, Q => n52194,
                           QN => n3319);
   REGS_reg_123_12_inst : DFF_X1 port map( D => n10385, CK => CLK, Q => n52195,
                           QN => n3320);
   REGS_reg_123_11_inst : DFF_X1 port map( D => n10384, CK => CLK, Q => n52196,
                           QN => n3321);
   REGS_reg_123_10_inst : DFF_X1 port map( D => n10383, CK => CLK, Q => n52197,
                           QN => n3322);
   REGS_reg_123_9_inst : DFF_X1 port map( D => n10382, CK => CLK, Q => n52198, 
                           QN => n3323);
   REGS_reg_123_8_inst : DFF_X1 port map( D => n10381, CK => CLK, Q => n52199, 
                           QN => n3324);
   REGS_reg_123_7_inst : DFF_X1 port map( D => n10380, CK => CLK, Q => n52200, 
                           QN => n3325);
   REGS_reg_123_6_inst : DFF_X1 port map( D => n10379, CK => CLK, Q => n52201, 
                           QN => n3326);
   REGS_reg_123_5_inst : DFF_X1 port map( D => n10378, CK => CLK, Q => n52202, 
                           QN => n3327);
   REGS_reg_123_4_inst : DFF_X1 port map( D => n10377, CK => CLK, Q => n52203, 
                           QN => n3328);
   REGS_reg_123_3_inst : DFF_X1 port map( D => n10376, CK => CLK, Q => n52204, 
                           QN => n3329);
   REGS_reg_123_2_inst : DFF_X1 port map( D => n10375, CK => CLK, Q => n52205, 
                           QN => n3330);
   REGS_reg_123_1_inst : DFF_X1 port map( D => n10374, CK => CLK, Q => n52206, 
                           QN => n3331);
   REGS_reg_123_0_inst : DFF_X1 port map( D => n10373, CK => CLK, Q => n52207, 
                           QN => n3332);
   REGS_reg_122_23_inst : DFF_X1 port map( D => n10428, CK => CLK, Q => n53632,
                           QN => n3333);
   REGS_reg_122_22_inst : DFF_X1 port map( D => n10427, CK => CLK, Q => n53633,
                           QN => n3334);
   REGS_reg_122_21_inst : DFF_X1 port map( D => n10426, CK => CLK, Q => n53634,
                           QN => n3335);
   REGS_reg_122_20_inst : DFF_X1 port map( D => n10425, CK => CLK, Q => n53635,
                           QN => n3336);
   REGS_reg_122_19_inst : DFF_X1 port map( D => n10424, CK => CLK, Q => n53636,
                           QN => n3337);
   REGS_reg_122_18_inst : DFF_X1 port map( D => n10423, CK => CLK, Q => n53637,
                           QN => n3338);
   REGS_reg_122_17_inst : DFF_X1 port map( D => n10422, CK => CLK, Q => n53638,
                           QN => n3339);
   REGS_reg_122_16_inst : DFF_X1 port map( D => n10421, CK => CLK, Q => n53639,
                           QN => n3340);
   REGS_reg_122_15_inst : DFF_X1 port map( D => n10420, CK => CLK, Q => n53640,
                           QN => n3341);
   REGS_reg_122_14_inst : DFF_X1 port map( D => n10419, CK => CLK, Q => n53641,
                           QN => n3342);
   REGS_reg_122_13_inst : DFF_X1 port map( D => n10418, CK => CLK, Q => n53642,
                           QN => n3343);
   REGS_reg_122_12_inst : DFF_X1 port map( D => n10417, CK => CLK, Q => n53643,
                           QN => n3344);
   REGS_reg_122_11_inst : DFF_X1 port map( D => n10416, CK => CLK, Q => n53644,
                           QN => n3345);
   REGS_reg_122_10_inst : DFF_X1 port map( D => n10415, CK => CLK, Q => n53645,
                           QN => n3346);
   REGS_reg_122_9_inst : DFF_X1 port map( D => n10414, CK => CLK, Q => n53646, 
                           QN => n3347);
   REGS_reg_122_8_inst : DFF_X1 port map( D => n10413, CK => CLK, Q => n53647, 
                           QN => n3348);
   REGS_reg_122_7_inst : DFF_X1 port map( D => n10412, CK => CLK, Q => n53648, 
                           QN => n3349);
   REGS_reg_122_6_inst : DFF_X1 port map( D => n10411, CK => CLK, Q => n53649, 
                           QN => n3350);
   REGS_reg_122_5_inst : DFF_X1 port map( D => n10410, CK => CLK, Q => n53650, 
                           QN => n3351);
   REGS_reg_122_4_inst : DFF_X1 port map( D => n10409, CK => CLK, Q => n53651, 
                           QN => n3352);
   REGS_reg_122_3_inst : DFF_X1 port map( D => n10408, CK => CLK, Q => n53652, 
                           QN => n3353);
   REGS_reg_122_2_inst : DFF_X1 port map( D => n10407, CK => CLK, Q => n53653, 
                           QN => n3354);
   REGS_reg_122_1_inst : DFF_X1 port map( D => n10406, CK => CLK, Q => n53654, 
                           QN => n3355);
   REGS_reg_122_0_inst : DFF_X1 port map( D => n10405, CK => CLK, Q => n53655, 
                           QN => n3356);
   REGS_reg_121_23_inst : DFF_X1 port map( D => n10460, CK => CLK, Q => n53656,
                           QN => n3357);
   REGS_reg_121_22_inst : DFF_X1 port map( D => n10459, CK => CLK, Q => n53657,
                           QN => n3358);
   REGS_reg_121_21_inst : DFF_X1 port map( D => n10458, CK => CLK, Q => n53658,
                           QN => n3359);
   REGS_reg_121_20_inst : DFF_X1 port map( D => n10457, CK => CLK, Q => n53659,
                           QN => n3360);
   REGS_reg_121_19_inst : DFF_X1 port map( D => n10456, CK => CLK, Q => n53660,
                           QN => n3361);
   REGS_reg_121_18_inst : DFF_X1 port map( D => n10455, CK => CLK, Q => n53661,
                           QN => n3362);
   REGS_reg_121_17_inst : DFF_X1 port map( D => n10454, CK => CLK, Q => n53662,
                           QN => n3363);
   REGS_reg_121_16_inst : DFF_X1 port map( D => n10453, CK => CLK, Q => n53663,
                           QN => n3364);
   REGS_reg_121_15_inst : DFF_X1 port map( D => n10452, CK => CLK, Q => n53664,
                           QN => n3365);
   REGS_reg_121_14_inst : DFF_X1 port map( D => n10451, CK => CLK, Q => n53665,
                           QN => n3366);
   REGS_reg_121_13_inst : DFF_X1 port map( D => n10450, CK => CLK, Q => n53666,
                           QN => n3367);
   REGS_reg_121_12_inst : DFF_X1 port map( D => n10449, CK => CLK, Q => n53667,
                           QN => n3368);
   REGS_reg_121_11_inst : DFF_X1 port map( D => n10448, CK => CLK, Q => n53668,
                           QN => n3369);
   REGS_reg_121_10_inst : DFF_X1 port map( D => n10447, CK => CLK, Q => n53669,
                           QN => n3370);
   REGS_reg_121_9_inst : DFF_X1 port map( D => n10446, CK => CLK, Q => n53670, 
                           QN => n3371);
   REGS_reg_121_8_inst : DFF_X1 port map( D => n10445, CK => CLK, Q => n53671, 
                           QN => n3372);
   REGS_reg_121_7_inst : DFF_X1 port map( D => n10444, CK => CLK, Q => n53672, 
                           QN => n3373);
   REGS_reg_121_6_inst : DFF_X1 port map( D => n10443, CK => CLK, Q => n53673, 
                           QN => n3374);
   REGS_reg_121_5_inst : DFF_X1 port map( D => n10442, CK => CLK, Q => n53674, 
                           QN => n3375);
   REGS_reg_121_4_inst : DFF_X1 port map( D => n10441, CK => CLK, Q => n53675, 
                           QN => n3376);
   REGS_reg_121_3_inst : DFF_X1 port map( D => n10440, CK => CLK, Q => n53676, 
                           QN => n3377);
   REGS_reg_121_2_inst : DFF_X1 port map( D => n10439, CK => CLK, Q => n53677, 
                           QN => n3378);
   REGS_reg_121_1_inst : DFF_X1 port map( D => n10438, CK => CLK, Q => n53678, 
                           QN => n3379);
   REGS_reg_121_0_inst : DFF_X1 port map( D => n10437, CK => CLK, Q => n53679, 
                           QN => n3380);
   REGS_reg_118_23_inst : DFF_X1 port map( D => n10556, CK => CLK, Q => n53680,
                           QN => n3381);
   REGS_reg_118_22_inst : DFF_X1 port map( D => n10555, CK => CLK, Q => n53681,
                           QN => n3382);
   REGS_reg_118_21_inst : DFF_X1 port map( D => n10554, CK => CLK, Q => n53682,
                           QN => n3383);
   REGS_reg_118_20_inst : DFF_X1 port map( D => n10553, CK => CLK, Q => n53683,
                           QN => n3384);
   REGS_reg_118_19_inst : DFF_X1 port map( D => n10552, CK => CLK, Q => n53684,
                           QN => n3385);
   REGS_reg_118_18_inst : DFF_X1 port map( D => n10551, CK => CLK, Q => n53685,
                           QN => n3386);
   REGS_reg_118_17_inst : DFF_X1 port map( D => n10550, CK => CLK, Q => n53686,
                           QN => n3387);
   REGS_reg_118_16_inst : DFF_X1 port map( D => n10549, CK => CLK, Q => n53687,
                           QN => n3388);
   REGS_reg_118_15_inst : DFF_X1 port map( D => n10548, CK => CLK, Q => n53688,
                           QN => n3389);
   REGS_reg_118_14_inst : DFF_X1 port map( D => n10547, CK => CLK, Q => n53689,
                           QN => n3390);
   REGS_reg_118_13_inst : DFF_X1 port map( D => n10546, CK => CLK, Q => n53690,
                           QN => n3391);
   REGS_reg_118_12_inst : DFF_X1 port map( D => n10545, CK => CLK, Q => n53691,
                           QN => n3392);
   REGS_reg_118_11_inst : DFF_X1 port map( D => n10544, CK => CLK, Q => n53692,
                           QN => n3393);
   REGS_reg_118_10_inst : DFF_X1 port map( D => n10543, CK => CLK, Q => n53693,
                           QN => n3394);
   REGS_reg_118_9_inst : DFF_X1 port map( D => n10542, CK => CLK, Q => n53694, 
                           QN => n3395);
   REGS_reg_118_8_inst : DFF_X1 port map( D => n10541, CK => CLK, Q => n53695, 
                           QN => n3396);
   REGS_reg_118_7_inst : DFF_X1 port map( D => n10540, CK => CLK, Q => n53696, 
                           QN => n3397);
   REGS_reg_118_6_inst : DFF_X1 port map( D => n10539, CK => CLK, Q => n53697, 
                           QN => n3398);
   REGS_reg_118_5_inst : DFF_X1 port map( D => n10538, CK => CLK, Q => n53698, 
                           QN => n3399);
   REGS_reg_118_4_inst : DFF_X1 port map( D => n10537, CK => CLK, Q => n53699, 
                           QN => n3400);
   REGS_reg_118_3_inst : DFF_X1 port map( D => n10536, CK => CLK, Q => n53700, 
                           QN => n3401);
   REGS_reg_118_2_inst : DFF_X1 port map( D => n10535, CK => CLK, Q => n53701, 
                           QN => n3402);
   REGS_reg_118_1_inst : DFF_X1 port map( D => n10534, CK => CLK, Q => n53702, 
                           QN => n3403);
   REGS_reg_118_0_inst : DFF_X1 port map( D => n10533, CK => CLK, Q => n53703, 
                           QN => n3404);
   REGS_reg_117_23_inst : DFF_X1 port map( D => n10588, CK => CLK, Q => n53704,
                           QN => n3405);
   REGS_reg_117_22_inst : DFF_X1 port map( D => n10587, CK => CLK, Q => n53705,
                           QN => n3406);
   REGS_reg_117_21_inst : DFF_X1 port map( D => n10586, CK => CLK, Q => n53706,
                           QN => n3407);
   REGS_reg_117_20_inst : DFF_X1 port map( D => n10585, CK => CLK, Q => n53707,
                           QN => n3408);
   REGS_reg_117_19_inst : DFF_X1 port map( D => n10584, CK => CLK, Q => n53708,
                           QN => n3457);
   REGS_reg_117_18_inst : DFF_X1 port map( D => n10583, CK => CLK, Q => n53709,
                           QN => n3458);
   REGS_reg_117_17_inst : DFF_X1 port map( D => n10582, CK => CLK, Q => n53710,
                           QN => n3459);
   REGS_reg_117_16_inst : DFF_X1 port map( D => n10581, CK => CLK, Q => n53711,
                           QN => n3460);
   REGS_reg_117_15_inst : DFF_X1 port map( D => n10580, CK => CLK, Q => n53712,
                           QN => n3461);
   REGS_reg_117_14_inst : DFF_X1 port map( D => n10579, CK => CLK, Q => n53713,
                           QN => n3462);
   REGS_reg_117_13_inst : DFF_X1 port map( D => n10578, CK => CLK, Q => n53714,
                           QN => n3463);
   REGS_reg_117_12_inst : DFF_X1 port map( D => n10577, CK => CLK, Q => n53715,
                           QN => n3464);
   REGS_reg_117_11_inst : DFF_X1 port map( D => n10576, CK => CLK, Q => n53716,
                           QN => n3465);
   REGS_reg_117_10_inst : DFF_X1 port map( D => n10575, CK => CLK, Q => n53717,
                           QN => n3466);
   REGS_reg_117_9_inst : DFF_X1 port map( D => n10574, CK => CLK, Q => n53718, 
                           QN => n3467);
   REGS_reg_117_8_inst : DFF_X1 port map( D => n10573, CK => CLK, Q => n53719, 
                           QN => n3468);
   REGS_reg_117_7_inst : DFF_X1 port map( D => n10572, CK => CLK, Q => n53720, 
                           QN => n3469);
   REGS_reg_117_6_inst : DFF_X1 port map( D => n10571, CK => CLK, Q => n53721, 
                           QN => n3470);
   REGS_reg_117_5_inst : DFF_X1 port map( D => n10570, CK => CLK, Q => n53722, 
                           QN => n3471);
   REGS_reg_117_4_inst : DFF_X1 port map( D => n10569, CK => CLK, Q => n53723, 
                           QN => n3472);
   REGS_reg_117_3_inst : DFF_X1 port map( D => n10568, CK => CLK, Q => n53724, 
                           QN => n3473);
   REGS_reg_117_2_inst : DFF_X1 port map( D => n10567, CK => CLK, Q => n53725, 
                           QN => n3474);
   REGS_reg_117_1_inst : DFF_X1 port map( D => n10566, CK => CLK, Q => n53726, 
                           QN => n3475);
   REGS_reg_117_0_inst : DFF_X1 port map( D => n10565, CK => CLK, Q => n53727, 
                           QN => n3476);
   REGS_reg_116_23_inst : DFF_X1 port map( D => n10620, CK => CLK, Q => n53728,
                           QN => n3477);
   REGS_reg_116_22_inst : DFF_X1 port map( D => n10619, CK => CLK, Q => n53729,
                           QN => n3478);
   REGS_reg_116_21_inst : DFF_X1 port map( D => n10618, CK => CLK, Q => n53730,
                           QN => n3479);
   REGS_reg_116_20_inst : DFF_X1 port map( D => n10617, CK => CLK, Q => n53731,
                           QN => n3480);
   REGS_reg_116_19_inst : DFF_X1 port map( D => n10616, CK => CLK, Q => n53732,
                           QN => n3481);
   REGS_reg_116_18_inst : DFF_X1 port map( D => n10615, CK => CLK, Q => n53733,
                           QN => n3482);
   REGS_reg_116_17_inst : DFF_X1 port map( D => n10614, CK => CLK, Q => n53734,
                           QN => n3483);
   REGS_reg_116_16_inst : DFF_X1 port map( D => n10613, CK => CLK, Q => n53735,
                           QN => n3484);
   REGS_reg_116_15_inst : DFF_X1 port map( D => n10612, CK => CLK, Q => n53736,
                           QN => n3485);
   REGS_reg_116_14_inst : DFF_X1 port map( D => n10611, CK => CLK, Q => n53737,
                           QN => n3486);
   REGS_reg_116_13_inst : DFF_X1 port map( D => n10610, CK => CLK, Q => n53738,
                           QN => n3487);
   REGS_reg_116_12_inst : DFF_X1 port map( D => n10609, CK => CLK, Q => n53739,
                           QN => n3488);
   REGS_reg_116_11_inst : DFF_X1 port map( D => n10608, CK => CLK, Q => n53740,
                           QN => n3489);
   REGS_reg_116_10_inst : DFF_X1 port map( D => n10607, CK => CLK, Q => n53741,
                           QN => n3490);
   REGS_reg_116_9_inst : DFF_X1 port map( D => n10606, CK => CLK, Q => n53742, 
                           QN => n3491);
   REGS_reg_116_8_inst : DFF_X1 port map( D => n10605, CK => CLK, Q => n53743, 
                           QN => n3492);
   REGS_reg_116_7_inst : DFF_X1 port map( D => n10604, CK => CLK, Q => n53744, 
                           QN => n3493);
   REGS_reg_116_6_inst : DFF_X1 port map( D => n10603, CK => CLK, Q => n53745, 
                           QN => n3494);
   REGS_reg_116_5_inst : DFF_X1 port map( D => n10602, CK => CLK, Q => n53746, 
                           QN => n3495);
   REGS_reg_116_4_inst : DFF_X1 port map( D => n10601, CK => CLK, Q => n53747, 
                           QN => n3496);
   REGS_reg_116_3_inst : DFF_X1 port map( D => n10600, CK => CLK, Q => n53748, 
                           QN => n3497);
   REGS_reg_116_2_inst : DFF_X1 port map( D => n10599, CK => CLK, Q => n53749, 
                           QN => n3498);
   REGS_reg_116_1_inst : DFF_X1 port map( D => n10598, CK => CLK, Q => n53750, 
                           QN => n3499);
   REGS_reg_116_0_inst : DFF_X1 port map( D => n10597, CK => CLK, Q => n53751, 
                           QN => n3500);
   REGS_reg_115_23_inst : DFF_X1 port map( D => n10652, CK => CLK, Q => n2791, 
                           QN => n3501);
   REGS_reg_115_22_inst : DFF_X1 port map( D => n10651, CK => CLK, Q => n2792, 
                           QN => n3502);
   REGS_reg_115_21_inst : DFF_X1 port map( D => n10650, CK => CLK, Q => n2793, 
                           QN => n3503);
   REGS_reg_115_20_inst : DFF_X1 port map( D => n10649, CK => CLK, Q => n2794, 
                           QN => n3504);
   REGS_reg_115_19_inst : DFF_X1 port map( D => n10648, CK => CLK, Q => n2795, 
                           QN => n3505);
   REGS_reg_115_18_inst : DFF_X1 port map( D => n10647, CK => CLK, Q => n2796, 
                           QN => n3506);
   REGS_reg_115_17_inst : DFF_X1 port map( D => n10646, CK => CLK, Q => n2797, 
                           QN => n3507);
   REGS_reg_115_16_inst : DFF_X1 port map( D => n10645, CK => CLK, Q => n2798, 
                           QN => n3508);
   REGS_reg_115_15_inst : DFF_X1 port map( D => n10644, CK => CLK, Q => n2799, 
                           QN => n3509);
   REGS_reg_115_14_inst : DFF_X1 port map( D => n10643, CK => CLK, Q => n2800, 
                           QN => n3510);
   REGS_reg_115_13_inst : DFF_X1 port map( D => n10642, CK => CLK, Q => n2801, 
                           QN => n3511);
   REGS_reg_115_12_inst : DFF_X1 port map( D => n10641, CK => CLK, Q => n2802, 
                           QN => n3512);
   REGS_reg_115_11_inst : DFF_X1 port map( D => n10640, CK => CLK, Q => n2803, 
                           QN => n3513);
   REGS_reg_115_10_inst : DFF_X1 port map( D => n10639, CK => CLK, Q => n2804, 
                           QN => n3514);
   REGS_reg_115_9_inst : DFF_X1 port map( D => n10638, CK => CLK, Q => n2805, 
                           QN => n3515);
   REGS_reg_115_8_inst : DFF_X1 port map( D => n10637, CK => CLK, Q => n2806, 
                           QN => n3516);
   REGS_reg_115_7_inst : DFF_X1 port map( D => n10636, CK => CLK, Q => n2807, 
                           QN => n3517);
   REGS_reg_115_6_inst : DFF_X1 port map( D => n10635, CK => CLK, Q => n2808, 
                           QN => n3518);
   REGS_reg_115_5_inst : DFF_X1 port map( D => n10634, CK => CLK, Q => n2809, 
                           QN => n3519);
   REGS_reg_115_4_inst : DFF_X1 port map( D => n10633, CK => CLK, Q => n2810, 
                           QN => n3520);
   REGS_reg_115_3_inst : DFF_X1 port map( D => n10632, CK => CLK, Q => n2811, 
                           QN => n3521);
   REGS_reg_115_2_inst : DFF_X1 port map( D => n10631, CK => CLK, Q => n2812, 
                           QN => n3522);
   REGS_reg_115_1_inst : DFF_X1 port map( D => n10630, CK => CLK, Q => n2813, 
                           QN => n3523);
   REGS_reg_115_0_inst : DFF_X1 port map( D => n10629, CK => CLK, Q => n2814, 
                           QN => n3524);
   REGS_reg_114_23_inst : DFF_X1 port map( D => n10684, CK => CLK, Q => n2815, 
                           QN => n3525);
   REGS_reg_114_22_inst : DFF_X1 port map( D => n10683, CK => CLK, Q => n2816, 
                           QN => n3526);
   REGS_reg_114_21_inst : DFF_X1 port map( D => n10682, CK => CLK, Q => n2817, 
                           QN => n3527);
   REGS_reg_114_20_inst : DFF_X1 port map( D => n10681, CK => CLK, Q => n2818, 
                           QN => n3528);
   REGS_reg_114_19_inst : DFF_X1 port map( D => n10680, CK => CLK, Q => n2819, 
                           QN => n3529);
   REGS_reg_114_18_inst : DFF_X1 port map( D => n10679, CK => CLK, Q => n2820, 
                           QN => n3530);
   REGS_reg_114_17_inst : DFF_X1 port map( D => n10678, CK => CLK, Q => n2821, 
                           QN => n3531);
   REGS_reg_114_16_inst : DFF_X1 port map( D => n10677, CK => CLK, Q => n2822, 
                           QN => n3532);
   REGS_reg_114_15_inst : DFF_X1 port map( D => n10676, CK => CLK, Q => n2823, 
                           QN => n3533);
   REGS_reg_114_14_inst : DFF_X1 port map( D => n10675, CK => CLK, Q => n2824, 
                           QN => n3534);
   REGS_reg_114_13_inst : DFF_X1 port map( D => n10674, CK => CLK, Q => n2825, 
                           QN => n3535);
   REGS_reg_114_12_inst : DFF_X1 port map( D => n10673, CK => CLK, Q => n2826, 
                           QN => n3536);
   REGS_reg_114_11_inst : DFF_X1 port map( D => n10672, CK => CLK, Q => n2827, 
                           QN => n3537);
   REGS_reg_114_10_inst : DFF_X1 port map( D => n10671, CK => CLK, Q => n2828, 
                           QN => n3538);
   REGS_reg_114_9_inst : DFF_X1 port map( D => n10670, CK => CLK, Q => n2829, 
                           QN => n3539);
   REGS_reg_114_8_inst : DFF_X1 port map( D => n10669, CK => CLK, Q => n2830, 
                           QN => n3540);
   REGS_reg_114_7_inst : DFF_X1 port map( D => n10668, CK => CLK, Q => n2831, 
                           QN => n3541);
   REGS_reg_114_6_inst : DFF_X1 port map( D => n10667, CK => CLK, Q => n2832, 
                           QN => n3542);
   REGS_reg_114_5_inst : DFF_X1 port map( D => n10666, CK => CLK, Q => n2833, 
                           QN => n3543);
   REGS_reg_114_4_inst : DFF_X1 port map( D => n10665, CK => CLK, Q => n2834, 
                           QN => n3544);
   REGS_reg_114_3_inst : DFF_X1 port map( D => n10664, CK => CLK, Q => n2835, 
                           QN => n3545);
   REGS_reg_114_2_inst : DFF_X1 port map( D => n10663, CK => CLK, Q => n2836, 
                           QN => n3546);
   REGS_reg_114_1_inst : DFF_X1 port map( D => n10662, CK => CLK, Q => n2837, 
                           QN => n3547);
   REGS_reg_114_0_inst : DFF_X1 port map( D => n10661, CK => CLK, Q => n2838, 
                           QN => n3548);
   REGS_reg_113_23_inst : DFF_X1 port map( D => n10716, CK => CLK, Q => n_1744,
                           QN => n3549);
   REGS_reg_113_22_inst : DFF_X1 port map( D => n10715, CK => CLK, Q => n_1745,
                           QN => n3550);
   REGS_reg_113_21_inst : DFF_X1 port map( D => n10714, CK => CLK, Q => n_1746,
                           QN => n3551);
   REGS_reg_113_20_inst : DFF_X1 port map( D => n10713, CK => CLK, Q => n_1747,
                           QN => n3552);
   REGS_reg_113_19_inst : DFF_X1 port map( D => n10712, CK => CLK, Q => n_1748,
                           QN => n3553);
   REGS_reg_113_18_inst : DFF_X1 port map( D => n10711, CK => CLK, Q => n_1749,
                           QN => n3554);
   REGS_reg_113_17_inst : DFF_X1 port map( D => n10710, CK => CLK, Q => n_1750,
                           QN => n3555);
   REGS_reg_113_16_inst : DFF_X1 port map( D => n10709, CK => CLK, Q => n_1751,
                           QN => n3556);
   REGS_reg_113_15_inst : DFF_X1 port map( D => n10708, CK => CLK, Q => n_1752,
                           QN => n3557);
   REGS_reg_113_14_inst : DFF_X1 port map( D => n10707, CK => CLK, Q => n_1753,
                           QN => n3558);
   REGS_reg_113_13_inst : DFF_X1 port map( D => n10706, CK => CLK, Q => n_1754,
                           QN => n3559);
   REGS_reg_113_12_inst : DFF_X1 port map( D => n10705, CK => CLK, Q => n_1755,
                           QN => n3560);
   REGS_reg_113_11_inst : DFF_X1 port map( D => n10704, CK => CLK, Q => n_1756,
                           QN => n3561);
   REGS_reg_113_10_inst : DFF_X1 port map( D => n10703, CK => CLK, Q => n_1757,
                           QN => n3562);
   REGS_reg_113_9_inst : DFF_X1 port map( D => n10702, CK => CLK, Q => n_1758, 
                           QN => n3563);
   REGS_reg_113_8_inst : DFF_X1 port map( D => n10701, CK => CLK, Q => n_1759, 
                           QN => n3564);
   REGS_reg_113_7_inst : DFF_X1 port map( D => n10700, CK => CLK, Q => n_1760, 
                           QN => n3565);
   REGS_reg_113_6_inst : DFF_X1 port map( D => n10699, CK => CLK, Q => n_1761, 
                           QN => n3566);
   REGS_reg_113_5_inst : DFF_X1 port map( D => n10698, CK => CLK, Q => n_1762, 
                           QN => n3567);
   REGS_reg_113_4_inst : DFF_X1 port map( D => n10697, CK => CLK, Q => n_1763, 
                           QN => n3568);
   REGS_reg_113_3_inst : DFF_X1 port map( D => n10696, CK => CLK, Q => n_1764, 
                           QN => n3569);
   REGS_reg_113_2_inst : DFF_X1 port map( D => n10695, CK => CLK, Q => n_1765, 
                           QN => n3570);
   REGS_reg_113_1_inst : DFF_X1 port map( D => n10694, CK => CLK, Q => n_1766, 
                           QN => n3571);
   REGS_reg_113_0_inst : DFF_X1 port map( D => n10693, CK => CLK, Q => n_1767, 
                           QN => n3572);
   REGS_reg_112_23_inst : DFF_X1 port map( D => n10748, CK => CLK, Q => n_1768,
                           QN => n3573);
   REGS_reg_112_22_inst : DFF_X1 port map( D => n10747, CK => CLK, Q => n_1769,
                           QN => n3574);
   REGS_reg_112_21_inst : DFF_X1 port map( D => n10746, CK => CLK, Q => n_1770,
                           QN => n3575);
   REGS_reg_112_20_inst : DFF_X1 port map( D => n10745, CK => CLK, Q => n_1771,
                           QN => n3576);
   REGS_reg_112_19_inst : DFF_X1 port map( D => n10744, CK => CLK, Q => n_1772,
                           QN => n3577);
   REGS_reg_112_18_inst : DFF_X1 port map( D => n10743, CK => CLK, Q => n_1773,
                           QN => n3578);
   REGS_reg_112_17_inst : DFF_X1 port map( D => n10742, CK => CLK, Q => n_1774,
                           QN => n3579);
   REGS_reg_112_16_inst : DFF_X1 port map( D => n10741, CK => CLK, Q => n_1775,
                           QN => n3580);
   REGS_reg_112_15_inst : DFF_X1 port map( D => n10740, CK => CLK, Q => n_1776,
                           QN => n3581);
   REGS_reg_112_14_inst : DFF_X1 port map( D => n10739, CK => CLK, Q => n_1777,
                           QN => n3582);
   REGS_reg_112_13_inst : DFF_X1 port map( D => n10738, CK => CLK, Q => n_1778,
                           QN => n3583);
   REGS_reg_112_12_inst : DFF_X1 port map( D => n10737, CK => CLK, Q => n_1779,
                           QN => n3584);
   REGS_reg_112_11_inst : DFF_X1 port map( D => n10736, CK => CLK, Q => n_1780,
                           QN => n3585);
   REGS_reg_112_10_inst : DFF_X1 port map( D => n10735, CK => CLK, Q => n_1781,
                           QN => n3586);
   REGS_reg_112_9_inst : DFF_X1 port map( D => n10734, CK => CLK, Q => n_1782, 
                           QN => n3587);
   REGS_reg_112_8_inst : DFF_X1 port map( D => n10733, CK => CLK, Q => n_1783, 
                           QN => n3588);
   REGS_reg_112_7_inst : DFF_X1 port map( D => n10732, CK => CLK, Q => n_1784, 
                           QN => n3589);
   REGS_reg_112_6_inst : DFF_X1 port map( D => n10731, CK => CLK, Q => n_1785, 
                           QN => n3590);
   REGS_reg_112_5_inst : DFF_X1 port map( D => n10730, CK => CLK, Q => n_1786, 
                           QN => n3591);
   REGS_reg_112_4_inst : DFF_X1 port map( D => n10729, CK => CLK, Q => n_1787, 
                           QN => n3592);
   REGS_reg_112_3_inst : DFF_X1 port map( D => n10728, CK => CLK, Q => n_1788, 
                           QN => n3593);
   REGS_reg_112_2_inst : DFF_X1 port map( D => n10727, CK => CLK, Q => n_1789, 
                           QN => n3594);
   REGS_reg_112_1_inst : DFF_X1 port map( D => n10726, CK => CLK, Q => n_1790, 
                           QN => n3595);
   REGS_reg_112_0_inst : DFF_X1 port map( D => n10725, CK => CLK, Q => n_1791, 
                           QN => n3596);
   REGS_reg_111_23_inst : DFF_X1 port map( D => n10780, CK => CLK, Q => n2439, 
                           QN => n5094);
   REGS_reg_111_22_inst : DFF_X1 port map( D => n10779, CK => CLK, Q => n2440, 
                           QN => n5095);
   REGS_reg_111_21_inst : DFF_X1 port map( D => n10778, CK => CLK, Q => n2441, 
                           QN => n5096);
   REGS_reg_111_20_inst : DFF_X1 port map( D => n10777, CK => CLK, Q => n2442, 
                           QN => n5097);
   REGS_reg_111_19_inst : DFF_X1 port map( D => n10776, CK => CLK, Q => n2443, 
                           QN => n5098);
   REGS_reg_111_18_inst : DFF_X1 port map( D => n10775, CK => CLK, Q => n2444, 
                           QN => n5099);
   REGS_reg_111_17_inst : DFF_X1 port map( D => n10774, CK => CLK, Q => n2445, 
                           QN => n5100);
   REGS_reg_111_16_inst : DFF_X1 port map( D => n10773, CK => CLK, Q => n2446, 
                           QN => n5101);
   REGS_reg_111_15_inst : DFF_X1 port map( D => n10772, CK => CLK, Q => n2447, 
                           QN => n5102);
   REGS_reg_111_14_inst : DFF_X1 port map( D => n10771, CK => CLK, Q => n2448, 
                           QN => n5103);
   REGS_reg_111_13_inst : DFF_X1 port map( D => n10770, CK => CLK, Q => n2449, 
                           QN => n5104);
   REGS_reg_111_12_inst : DFF_X1 port map( D => n10769, CK => CLK, Q => n2450, 
                           QN => n5105);
   REGS_reg_111_11_inst : DFF_X1 port map( D => n10768, CK => CLK, Q => n2451, 
                           QN => n5106);
   REGS_reg_111_10_inst : DFF_X1 port map( D => n10767, CK => CLK, Q => n2452, 
                           QN => n5107);
   REGS_reg_111_9_inst : DFF_X1 port map( D => n10766, CK => CLK, Q => n2453, 
                           QN => n5108);
   REGS_reg_111_8_inst : DFF_X1 port map( D => n10765, CK => CLK, Q => n2454, 
                           QN => n5109);
   REGS_reg_111_7_inst : DFF_X1 port map( D => n10764, CK => CLK, Q => n2455, 
                           QN => n5110);
   REGS_reg_111_6_inst : DFF_X1 port map( D => n10763, CK => CLK, Q => n2456, 
                           QN => n5111);
   REGS_reg_111_5_inst : DFF_X1 port map( D => n10762, CK => CLK, Q => n2457, 
                           QN => n5112);
   REGS_reg_111_4_inst : DFF_X1 port map( D => n10761, CK => CLK, Q => n2458, 
                           QN => n5113);
   REGS_reg_111_3_inst : DFF_X1 port map( D => n10760, CK => CLK, Q => n2459, 
                           QN => n5114);
   REGS_reg_111_2_inst : DFF_X1 port map( D => n10759, CK => CLK, Q => n2460, 
                           QN => n5115);
   REGS_reg_111_1_inst : DFF_X1 port map( D => n10758, CK => CLK, Q => n2461, 
                           QN => n5116);
   REGS_reg_111_0_inst : DFF_X1 port map( D => n10757, CK => CLK, Q => n2462, 
                           QN => n5117);
   REGS_reg_110_23_inst : DFF_X1 port map( D => n10812, CK => CLK, Q => n2887, 
                           QN => n3597);
   REGS_reg_110_22_inst : DFF_X1 port map( D => n10811, CK => CLK, Q => n2888, 
                           QN => n3598);
   REGS_reg_110_21_inst : DFF_X1 port map( D => n10810, CK => CLK, Q => n2889, 
                           QN => n3599);
   REGS_reg_110_20_inst : DFF_X1 port map( D => n10809, CK => CLK, Q => n2890, 
                           QN => n3600);
   REGS_reg_110_19_inst : DFF_X1 port map( D => n10808, CK => CLK, Q => n2891, 
                           QN => n3601);
   REGS_reg_110_18_inst : DFF_X1 port map( D => n10807, CK => CLK, Q => n2892, 
                           QN => n3602);
   REGS_reg_110_17_inst : DFF_X1 port map( D => n10806, CK => CLK, Q => n2893, 
                           QN => n3603);
   REGS_reg_110_16_inst : DFF_X1 port map( D => n10805, CK => CLK, Q => n2894, 
                           QN => n3604);
   REGS_reg_110_15_inst : DFF_X1 port map( D => n10804, CK => CLK, Q => n2895, 
                           QN => n3605);
   REGS_reg_110_14_inst : DFF_X1 port map( D => n10803, CK => CLK, Q => n2896, 
                           QN => n3606);
   REGS_reg_110_13_inst : DFF_X1 port map( D => n10802, CK => CLK, Q => n2897, 
                           QN => n3607);
   REGS_reg_110_12_inst : DFF_X1 port map( D => n10801, CK => CLK, Q => n2898, 
                           QN => n3608);
   REGS_reg_110_11_inst : DFF_X1 port map( D => n10800, CK => CLK, Q => n2899, 
                           QN => n3609);
   REGS_reg_110_10_inst : DFF_X1 port map( D => n10799, CK => CLK, Q => n2900, 
                           QN => n3610);
   REGS_reg_110_9_inst : DFF_X1 port map( D => n10798, CK => CLK, Q => n2901, 
                           QN => n3611);
   REGS_reg_110_8_inst : DFF_X1 port map( D => n10797, CK => CLK, Q => n2902, 
                           QN => n3612);
   REGS_reg_110_7_inst : DFF_X1 port map( D => n10796, CK => CLK, Q => n2903, 
                           QN => n3613);
   REGS_reg_110_6_inst : DFF_X1 port map( D => n10795, CK => CLK, Q => n2904, 
                           QN => n3614);
   REGS_reg_110_5_inst : DFF_X1 port map( D => n10794, CK => CLK, Q => n2905, 
                           QN => n3615);
   REGS_reg_110_4_inst : DFF_X1 port map( D => n10793, CK => CLK, Q => n2906, 
                           QN => n3616);
   REGS_reg_110_3_inst : DFF_X1 port map( D => n10792, CK => CLK, Q => n2483, 
                           QN => n5118);
   REGS_reg_110_2_inst : DFF_X1 port map( D => n10791, CK => CLK, Q => n2484, 
                           QN => n5119);
   REGS_reg_110_1_inst : DFF_X1 port map( D => n10790, CK => CLK, Q => n2485, 
                           QN => n5120);
   REGS_reg_110_0_inst : DFF_X1 port map( D => n10789, CK => CLK, Q => n2486, 
                           QN => n5121);
   REGS_reg_107_23_inst : DFF_X1 port map( D => n10908, CK => CLK, Q => n16563,
                           QN => n5122);
   REGS_reg_107_22_inst : DFF_X1 port map( D => n10907, CK => CLK, Q => n16562,
                           QN => n5123);
   REGS_reg_107_21_inst : DFF_X1 port map( D => n10906, CK => CLK, Q => n16561,
                           QN => n5124);
   REGS_reg_107_20_inst : DFF_X1 port map( D => n10905, CK => CLK, Q => n16560,
                           QN => n5125);
   REGS_reg_107_19_inst : DFF_X1 port map( D => n10904, CK => CLK, Q => n15439,
                           QN => n3617);
   REGS_reg_107_18_inst : DFF_X1 port map( D => n10903, CK => CLK, Q => n15438,
                           QN => n3618);
   REGS_reg_107_17_inst : DFF_X1 port map( D => n10902, CK => CLK, Q => n15437,
                           QN => n3619);
   REGS_reg_107_16_inst : DFF_X1 port map( D => n10901, CK => CLK, Q => n15436,
                           QN => n3620);
   REGS_reg_107_15_inst : DFF_X1 port map( D => n10900, CK => CLK, Q => n15435,
                           QN => n3645);
   REGS_reg_107_14_inst : DFF_X1 port map( D => n10899, CK => CLK, Q => n15434,
                           QN => n3646);
   REGS_reg_107_13_inst : DFF_X1 port map( D => n10898, CK => CLK, Q => n15433,
                           QN => n3647);
   REGS_reg_107_12_inst : DFF_X1 port map( D => n10897, CK => CLK, Q => n15432,
                           QN => n3648);
   REGS_reg_107_11_inst : DFF_X1 port map( D => n10896, CK => CLK, Q => n16559,
                           QN => n5126);
   REGS_reg_107_10_inst : DFF_X1 port map( D => n10895, CK => CLK, Q => n16558,
                           QN => n5127);
   REGS_reg_107_9_inst : DFF_X1 port map( D => n10894, CK => CLK, Q => n16557, 
                           QN => n5128);
   REGS_reg_107_8_inst : DFF_X1 port map( D => n10893, CK => CLK, Q => n16556, 
                           QN => n5129);
   REGS_reg_107_7_inst : DFF_X1 port map( D => n10892, CK => CLK, Q => n16555, 
                           QN => n5130);
   REGS_reg_107_6_inst : DFF_X1 port map( D => n10891, CK => CLK, Q => n16554, 
                           QN => n5131);
   REGS_reg_107_5_inst : DFF_X1 port map( D => n10890, CK => CLK, Q => n15431, 
                           QN => n3649);
   REGS_reg_107_4_inst : DFF_X1 port map( D => n10889, CK => CLK, Q => n15430, 
                           QN => n3650);
   REGS_reg_107_3_inst : DFF_X1 port map( D => n10888, CK => CLK, Q => n15429, 
                           QN => n3651);
   REGS_reg_107_2_inst : DFF_X1 port map( D => n10887, CK => CLK, Q => n15428, 
                           QN => n3652);
   REGS_reg_107_1_inst : DFF_X1 port map( D => n10886, CK => CLK, Q => n15427, 
                           QN => n3653);
   REGS_reg_107_0_inst : DFF_X1 port map( D => n10885, CK => CLK, Q => n15402, 
                           QN => n3654);
   REGS_reg_106_23_inst : DFF_X1 port map( D => n10940, CK => CLK, Q => n15706,
                           QN => n3655);
   REGS_reg_106_22_inst : DFF_X1 port map( D => n10939, CK => CLK, Q => n15703,
                           QN => n3656);
   REGS_reg_106_21_inst : DFF_X1 port map( D => n10938, CK => CLK, Q => n15700,
                           QN => n3657);
   REGS_reg_106_20_inst : DFF_X1 port map( D => n10937, CK => CLK, Q => n15697,
                           QN => n3658);
   REGS_reg_106_19_inst : DFF_X1 port map( D => n10936, CK => CLK, Q => n15401,
                           QN => n3659);
   REGS_reg_106_18_inst : DFF_X1 port map( D => n10935, CK => CLK, Q => n15400,
                           QN => n3660);
   REGS_reg_106_17_inst : DFF_X1 port map( D => n10934, CK => CLK, Q => n15399,
                           QN => n3661);
   REGS_reg_106_16_inst : DFF_X1 port map( D => n10933, CK => CLK, Q => n15398,
                           QN => n3662);
   REGS_reg_106_15_inst : DFF_X1 port map( D => n10932, CK => CLK, Q => n15397,
                           QN => n3663);
   REGS_reg_106_14_inst : DFF_X1 port map( D => n10931, CK => CLK, Q => n15396,
                           QN => n3664);
   REGS_reg_106_13_inst : DFF_X1 port map( D => n10930, CK => CLK, Q => n15395,
                           QN => n3665);
   REGS_reg_106_12_inst : DFF_X1 port map( D => n10929, CK => CLK, Q => n15386,
                           QN => n3666);
   REGS_reg_106_11_inst : DFF_X1 port map( D => n10928, CK => CLK, Q => n15694,
                           QN => n3667);
   REGS_reg_106_10_inst : DFF_X1 port map( D => n10927, CK => CLK, Q => n15691,
                           QN => n3668);
   REGS_reg_106_9_inst : DFF_X1 port map( D => n10926, CK => CLK, Q => n15688, 
                           QN => n3669);
   REGS_reg_106_8_inst : DFF_X1 port map( D => n10925, CK => CLK, Q => n15685, 
                           QN => n3670);
   REGS_reg_106_7_inst : DFF_X1 port map( D => n10924, CK => CLK, Q => n15729, 
                           QN => n3671);
   REGS_reg_106_6_inst : DFF_X1 port map( D => n10923, CK => CLK, Q => n15726, 
                           QN => n3672);
   REGS_reg_106_5_inst : DFF_X1 port map( D => n10922, CK => CLK, Q => n15385, 
                           QN => n3673);
   REGS_reg_106_4_inst : DFF_X1 port map( D => n10921, CK => CLK, Q => n15384, 
                           QN => n3674);
   REGS_reg_106_3_inst : DFF_X1 port map( D => n10920, CK => CLK, Q => n15383, 
                           QN => n3675);
   REGS_reg_106_2_inst : DFF_X1 port map( D => n10919, CK => CLK, Q => n15382, 
                           QN => n3676);
   REGS_reg_106_1_inst : DFF_X1 port map( D => n10918, CK => CLK, Q => n15381, 
                           QN => n3677);
   REGS_reg_106_0_inst : DFF_X1 port map( D => n10917, CK => CLK, Q => n15380, 
                           QN => n3678);
   REGS_reg_105_23_inst : DFF_X1 port map( D => n10972, CK => CLK, Q => n_1792,
                           QN => n3679);
   REGS_reg_105_22_inst : DFF_X1 port map( D => n10971, CK => CLK, Q => n_1793,
                           QN => n3680);
   REGS_reg_105_21_inst : DFF_X1 port map( D => n10970, CK => CLK, Q => n_1794,
                           QN => n3681);
   REGS_reg_105_20_inst : DFF_X1 port map( D => n10969, CK => CLK, Q => n_1795,
                           QN => n3682);
   REGS_reg_105_19_inst : DFF_X1 port map( D => n10968, CK => CLK, Q => n_1796,
                           QN => n3683);
   REGS_reg_105_18_inst : DFF_X1 port map( D => n10967, CK => CLK, Q => n_1797,
                           QN => n3684);
   REGS_reg_105_17_inst : DFF_X1 port map( D => n10966, CK => CLK, Q => n_1798,
                           QN => n3685);
   REGS_reg_105_16_inst : DFF_X1 port map( D => n10965, CK => CLK, Q => n_1799,
                           QN => n3686);
   REGS_reg_105_15_inst : DFF_X1 port map( D => n10964, CK => CLK, Q => n_1800,
                           QN => n3687);
   REGS_reg_105_14_inst : DFF_X1 port map( D => n10963, CK => CLK, Q => n_1801,
                           QN => n3688);
   REGS_reg_105_13_inst : DFF_X1 port map( D => n10962, CK => CLK, Q => n_1802,
                           QN => n3689);
   REGS_reg_105_12_inst : DFF_X1 port map( D => n10961, CK => CLK, Q => n_1803,
                           QN => n3690);
   REGS_reg_105_11_inst : DFF_X1 port map( D => n10960, CK => CLK, Q => n_1804,
                           QN => n3691);
   REGS_reg_105_10_inst : DFF_X1 port map( D => n10959, CK => CLK, Q => n_1805,
                           QN => n3692);
   REGS_reg_105_9_inst : DFF_X1 port map( D => n10958, CK => CLK, Q => n_1806, 
                           QN => n3693);
   REGS_reg_105_8_inst : DFF_X1 port map( D => n10957, CK => CLK, Q => n_1807, 
                           QN => n3694);
   REGS_reg_105_7_inst : DFF_X1 port map( D => n10956, CK => CLK, Q => n_1808, 
                           QN => n3695);
   REGS_reg_105_6_inst : DFF_X1 port map( D => n10955, CK => CLK, Q => n_1809, 
                           QN => n3696);
   REGS_reg_105_5_inst : DFF_X1 port map( D => n10954, CK => CLK, Q => n_1810, 
                           QN => n3697);
   REGS_reg_105_4_inst : DFF_X1 port map( D => n10953, CK => CLK, Q => n_1811, 
                           QN => n3698);
   REGS_reg_105_3_inst : DFF_X1 port map( D => n10952, CK => CLK, Q => n_1812, 
                           QN => n3699);
   REGS_reg_105_2_inst : DFF_X1 port map( D => n10951, CK => CLK, Q => n_1813, 
                           QN => n3700);
   REGS_reg_105_1_inst : DFF_X1 port map( D => n10950, CK => CLK, Q => n_1814, 
                           QN => n3701);
   REGS_reg_105_0_inst : DFF_X1 port map( D => n10949, CK => CLK, Q => n_1815, 
                           QN => n3702);
   REGS_reg_104_23_inst : DFF_X1 port map( D => n11004, CK => CLK, Q => n_1816,
                           QN => n3703);
   REGS_reg_104_22_inst : DFF_X1 port map( D => n11003, CK => CLK, Q => n_1817,
                           QN => n3704);
   REGS_reg_104_21_inst : DFF_X1 port map( D => n11002, CK => CLK, Q => n_1818,
                           QN => n3705);
   REGS_reg_104_20_inst : DFF_X1 port map( D => n11001, CK => CLK, Q => n_1819,
                           QN => n3706);
   REGS_reg_104_19_inst : DFF_X1 port map( D => n11000, CK => CLK, Q => n_1820,
                           QN => n3707);
   REGS_reg_104_18_inst : DFF_X1 port map( D => n10999, CK => CLK, Q => n_1821,
                           QN => n3708);
   REGS_reg_104_17_inst : DFF_X1 port map( D => n10998, CK => CLK, Q => n_1822,
                           QN => n3709);
   REGS_reg_104_16_inst : DFF_X1 port map( D => n10997, CK => CLK, Q => n_1823,
                           QN => n3710);
   REGS_reg_104_15_inst : DFF_X1 port map( D => n10996, CK => CLK, Q => n_1824,
                           QN => n3711);
   REGS_reg_104_14_inst : DFF_X1 port map( D => n10995, CK => CLK, Q => n_1825,
                           QN => n3712);
   REGS_reg_104_13_inst : DFF_X1 port map( D => n10994, CK => CLK, Q => n_1826,
                           QN => n3713);
   REGS_reg_104_12_inst : DFF_X1 port map( D => n10993, CK => CLK, Q => n_1827,
                           QN => n3714);
   REGS_reg_104_11_inst : DFF_X1 port map( D => n10992, CK => CLK, Q => n_1828,
                           QN => n3715);
   REGS_reg_104_10_inst : DFF_X1 port map( D => n10991, CK => CLK, Q => n_1829,
                           QN => n3716);
   REGS_reg_104_9_inst : DFF_X1 port map( D => n10990, CK => CLK, Q => n_1830, 
                           QN => n3717);
   REGS_reg_104_8_inst : DFF_X1 port map( D => n10989, CK => CLK, Q => n_1831, 
                           QN => n3718);
   REGS_reg_104_7_inst : DFF_X1 port map( D => n10988, CK => CLK, Q => n_1832, 
                           QN => n3719);
   REGS_reg_104_6_inst : DFF_X1 port map( D => n10987, CK => CLK, Q => n_1833, 
                           QN => n3720);
   REGS_reg_104_5_inst : DFF_X1 port map( D => n10986, CK => CLK, Q => n_1834, 
                           QN => n3721);
   REGS_reg_104_4_inst : DFF_X1 port map( D => n10985, CK => CLK, Q => n_1835, 
                           QN => n3722);
   REGS_reg_104_3_inst : DFF_X1 port map( D => n10984, CK => CLK, Q => n_1836, 
                           QN => n3723);
   REGS_reg_104_2_inst : DFF_X1 port map( D => n10983, CK => CLK, Q => n_1837, 
                           QN => n3724);
   REGS_reg_104_1_inst : DFF_X1 port map( D => n10982, CK => CLK, Q => n_1838, 
                           QN => n3725);
   REGS_reg_104_0_inst : DFF_X1 port map( D => n10981, CK => CLK, Q => n_1839, 
                           QN => n3726);
   REGS_reg_103_23_inst : DFF_X1 port map( D => n11036, CK => CLK, Q => n2979, 
                           QN => n3727);
   REGS_reg_103_22_inst : DFF_X1 port map( D => n11035, CK => CLK, Q => n2980, 
                           QN => n3728);
   REGS_reg_103_21_inst : DFF_X1 port map( D => n11034, CK => CLK, Q => n2981, 
                           QN => n3729);
   REGS_reg_103_20_inst : DFF_X1 port map( D => n11033, CK => CLK, Q => n2982, 
                           QN => n3730);
   REGS_reg_103_19_inst : DFF_X1 port map( D => n11032, CK => CLK, Q => n2983, 
                           QN => n3731);
   REGS_reg_103_18_inst : DFF_X1 port map( D => n11031, CK => CLK, Q => n2984, 
                           QN => n3732);
   REGS_reg_103_17_inst : DFF_X1 port map( D => n11030, CK => CLK, Q => n2985, 
                           QN => n3733);
   REGS_reg_103_16_inst : DFF_X1 port map( D => n11029, CK => CLK, Q => n2986, 
                           QN => n3734);
   REGS_reg_103_15_inst : DFF_X1 port map( D => n11028, CK => CLK, Q => n2987, 
                           QN => n3735);
   REGS_reg_103_14_inst : DFF_X1 port map( D => n11027, CK => CLK, Q => n2988, 
                           QN => n3736);
   REGS_reg_103_13_inst : DFF_X1 port map( D => n11026, CK => CLK, Q => n2989, 
                           QN => n3737);
   REGS_reg_103_12_inst : DFF_X1 port map( D => n11025, CK => CLK, Q => n2990, 
                           QN => n3738);
   REGS_reg_103_11_inst : DFF_X1 port map( D => n11024, CK => CLK, Q => n2991, 
                           QN => n3739);
   REGS_reg_103_10_inst : DFF_X1 port map( D => n11023, CK => CLK, Q => n2992, 
                           QN => n3740);
   REGS_reg_103_9_inst : DFF_X1 port map( D => n11022, CK => CLK, Q => n2993, 
                           QN => n3741);
   REGS_reg_103_8_inst : DFF_X1 port map( D => n11021, CK => CLK, Q => n2994, 
                           QN => n3742);
   REGS_reg_103_7_inst : DFF_X1 port map( D => n11020, CK => CLK, Q => n2995, 
                           QN => n3743);
   REGS_reg_103_6_inst : DFF_X1 port map( D => n11019, CK => CLK, Q => n2996, 
                           QN => n3744);
   REGS_reg_103_5_inst : DFF_X1 port map( D => n11018, CK => CLK, Q => n2997, 
                           QN => n3745);
   REGS_reg_103_4_inst : DFF_X1 port map( D => n11017, CK => CLK, Q => n2998, 
                           QN => n3746);
   REGS_reg_103_3_inst : DFF_X1 port map( D => n11016, CK => CLK, Q => n2999, 
                           QN => n3747);
   REGS_reg_103_2_inst : DFF_X1 port map( D => n11015, CK => CLK, Q => n3000, 
                           QN => n3748);
   REGS_reg_103_1_inst : DFF_X1 port map( D => n11014, CK => CLK, Q => n3001, 
                           QN => n3749);
   REGS_reg_103_0_inst : DFF_X1 port map( D => n11013, CK => CLK, Q => n3002, 
                           QN => n3750);
   REGS_reg_102_23_inst : DFF_X1 port map( D => n11068, CK => CLK, Q => n3003, 
                           QN => n3751);
   REGS_reg_102_22_inst : DFF_X1 port map( D => n11067, CK => CLK, Q => n3004, 
                           QN => n3752);
   REGS_reg_102_21_inst : DFF_X1 port map( D => n11066, CK => CLK, Q => n3005, 
                           QN => n3753);
   REGS_reg_102_20_inst : DFF_X1 port map( D => n11065, CK => CLK, Q => n3006, 
                           QN => n3754);
   REGS_reg_102_19_inst : DFF_X1 port map( D => n11064, CK => CLK, Q => n3007, 
                           QN => n3755);
   REGS_reg_102_18_inst : DFF_X1 port map( D => n11063, CK => CLK, Q => n3008, 
                           QN => n3756);
   REGS_reg_102_17_inst : DFF_X1 port map( D => n11062, CK => CLK, Q => n3009, 
                           QN => n3757);
   REGS_reg_102_16_inst : DFF_X1 port map( D => n11061, CK => CLK, Q => n3010, 
                           QN => n3758);
   REGS_reg_102_15_inst : DFF_X1 port map( D => n11060, CK => CLK, Q => n3011, 
                           QN => n3759);
   REGS_reg_102_14_inst : DFF_X1 port map( D => n11059, CK => CLK, Q => n3012, 
                           QN => n3760);
   REGS_reg_102_13_inst : DFF_X1 port map( D => n11058, CK => CLK, Q => n3013, 
                           QN => n3761);
   REGS_reg_102_12_inst : DFF_X1 port map( D => n11057, CK => CLK, Q => n3014, 
                           QN => n3762);
   REGS_reg_102_11_inst : DFF_X1 port map( D => n11056, CK => CLK, Q => n3015, 
                           QN => n3763);
   REGS_reg_102_10_inst : DFF_X1 port map( D => n11055, CK => CLK, Q => n3016, 
                           QN => n3764);
   REGS_reg_102_9_inst : DFF_X1 port map( D => n11054, CK => CLK, Q => n3017, 
                           QN => n3765);
   REGS_reg_102_8_inst : DFF_X1 port map( D => n11053, CK => CLK, Q => n3018, 
                           QN => n3766);
   REGS_reg_102_7_inst : DFF_X1 port map( D => n11052, CK => CLK, Q => n3019, 
                           QN => n3767);
   REGS_reg_102_6_inst : DFF_X1 port map( D => n11051, CK => CLK, Q => n3020, 
                           QN => n3768);
   REGS_reg_102_5_inst : DFF_X1 port map( D => n11050, CK => CLK, Q => n3021, 
                           QN => n3769);
   REGS_reg_102_4_inst : DFF_X1 port map( D => n11049, CK => CLK, Q => n3022, 
                           QN => n3770);
   REGS_reg_102_3_inst : DFF_X1 port map( D => n11048, CK => CLK, Q => n3023, 
                           QN => n3771);
   REGS_reg_102_2_inst : DFF_X1 port map( D => n11047, CK => CLK, Q => n3024, 
                           QN => n3772);
   REGS_reg_102_1_inst : DFF_X1 port map( D => n11046, CK => CLK, Q => n3025, 
                           QN => n3773);
   REGS_reg_102_0_inst : DFF_X1 port map( D => n11045, CK => CLK, Q => n3026, 
                           QN => n3774);
   REGS_reg_101_23_inst : DFF_X1 port map( D => n11100, CK => CLK, Q => n53916,
                           QN => n3775);
   REGS_reg_101_22_inst : DFF_X1 port map( D => n11099, CK => CLK, Q => n53917,
                           QN => n3776);
   REGS_reg_101_21_inst : DFF_X1 port map( D => n11098, CK => CLK, Q => n53918,
                           QN => n3777);
   REGS_reg_101_20_inst : DFF_X1 port map( D => n11097, CK => CLK, Q => n53919,
                           QN => n3778);
   REGS_reg_101_19_inst : DFF_X1 port map( D => n11096, CK => CLK, Q => n53920,
                           QN => n3779);
   REGS_reg_101_18_inst : DFF_X1 port map( D => n11095, CK => CLK, Q => n53921,
                           QN => n3780);
   REGS_reg_101_17_inst : DFF_X1 port map( D => n11094, CK => CLK, Q => n53922,
                           QN => n3781);
   REGS_reg_101_16_inst : DFF_X1 port map( D => n11093, CK => CLK, Q => n53923,
                           QN => n3782);
   REGS_reg_101_15_inst : DFF_X1 port map( D => n11092, CK => CLK, Q => n53924,
                           QN => n3783);
   REGS_reg_101_14_inst : DFF_X1 port map( D => n11091, CK => CLK, Q => n53925,
                           QN => n3784);
   REGS_reg_101_13_inst : DFF_X1 port map( D => n11090, CK => CLK, Q => n53926,
                           QN => n3785);
   REGS_reg_101_12_inst : DFF_X1 port map( D => n11089, CK => CLK, Q => n53927,
                           QN => n3786);
   REGS_reg_101_11_inst : DFF_X1 port map( D => n11088, CK => CLK, Q => n53928,
                           QN => n3787);
   REGS_reg_101_10_inst : DFF_X1 port map( D => n11087, CK => CLK, Q => n53929,
                           QN => n3788);
   REGS_reg_101_9_inst : DFF_X1 port map( D => n11086, CK => CLK, Q => n53930, 
                           QN => n3789);
   REGS_reg_101_8_inst : DFF_X1 port map( D => n11085, CK => CLK, Q => n53931, 
                           QN => n3790);
   REGS_reg_101_7_inst : DFF_X1 port map( D => n11084, CK => CLK, Q => n53932, 
                           QN => n3791);
   REGS_reg_101_6_inst : DFF_X1 port map( D => n11083, CK => CLK, Q => n53933, 
                           QN => n3792);
   REGS_reg_101_5_inst : DFF_X1 port map( D => n11082, CK => CLK, Q => n53934, 
                           QN => n3793);
   REGS_reg_101_4_inst : DFF_X1 port map( D => n11081, CK => CLK, Q => n53935, 
                           QN => n3794);
   REGS_reg_101_3_inst : DFF_X1 port map( D => n11080, CK => CLK, Q => n53936, 
                           QN => n3795);
   REGS_reg_101_2_inst : DFF_X1 port map( D => n11079, CK => CLK, Q => n53937, 
                           QN => n3796);
   REGS_reg_101_1_inst : DFF_X1 port map( D => n11078, CK => CLK, Q => n53938, 
                           QN => n3797);
   REGS_reg_101_0_inst : DFF_X1 port map( D => n11077, CK => CLK, Q => n53939, 
                           QN => n3798);
   REGS_reg_100_23_inst : DFF_X1 port map( D => n11132, CK => CLK, Q => n53940,
                           QN => n3799);
   REGS_reg_100_22_inst : DFF_X1 port map( D => n11131, CK => CLK, Q => n53941,
                           QN => n3800);
   REGS_reg_100_21_inst : DFF_X1 port map( D => n11130, CK => CLK, Q => n53942,
                           QN => n3801);
   REGS_reg_100_20_inst : DFF_X1 port map( D => n11129, CK => CLK, Q => n53943,
                           QN => n3802);
   REGS_reg_100_19_inst : DFF_X1 port map( D => n11128, CK => CLK, Q => n53944,
                           QN => n3803);
   REGS_reg_100_18_inst : DFF_X1 port map( D => n11127, CK => CLK, Q => n53945,
                           QN => n3804);
   REGS_reg_100_17_inst : DFF_X1 port map( D => n11126, CK => CLK, Q => n53946,
                           QN => n3805);
   REGS_reg_100_16_inst : DFF_X1 port map( D => n11125, CK => CLK, Q => n53947,
                           QN => n3806);
   REGS_reg_100_15_inst : DFF_X1 port map( D => n11124, CK => CLK, Q => n53948,
                           QN => n3807);
   REGS_reg_100_14_inst : DFF_X1 port map( D => n11123, CK => CLK, Q => n53949,
                           QN => n3808);
   REGS_reg_100_13_inst : DFF_X1 port map( D => n11122, CK => CLK, Q => n53950,
                           QN => n3809);
   REGS_reg_100_12_inst : DFF_X1 port map( D => n11121, CK => CLK, Q => n53951,
                           QN => n3810);
   REGS_reg_100_11_inst : DFF_X1 port map( D => n11120, CK => CLK, Q => n53952,
                           QN => n3811);
   REGS_reg_100_10_inst : DFF_X1 port map( D => n11119, CK => CLK, Q => n53953,
                           QN => n3812);
   REGS_reg_100_9_inst : DFF_X1 port map( D => n11118, CK => CLK, Q => n53954, 
                           QN => n3813);
   REGS_reg_100_8_inst : DFF_X1 port map( D => n11117, CK => CLK, Q => n53955, 
                           QN => n3814);
   REGS_reg_100_7_inst : DFF_X1 port map( D => n11116, CK => CLK, Q => n53956, 
                           QN => n3815);
   REGS_reg_100_6_inst : DFF_X1 port map( D => n11115, CK => CLK, Q => n53957, 
                           QN => n3816);
   REGS_reg_100_5_inst : DFF_X1 port map( D => n11114, CK => CLK, Q => n53958, 
                           QN => n3817);
   REGS_reg_100_4_inst : DFF_X1 port map( D => n11113, CK => CLK, Q => n53959, 
                           QN => n3818);
   REGS_reg_100_3_inst : DFF_X1 port map( D => n11112, CK => CLK, Q => n53960, 
                           QN => n3819);
   REGS_reg_100_2_inst : DFF_X1 port map( D => n11111, CK => CLK, Q => n53961, 
                           QN => n3820);
   REGS_reg_100_1_inst : DFF_X1 port map( D => n11110, CK => CLK, Q => n53962, 
                           QN => n3821);
   REGS_reg_100_0_inst : DFF_X1 port map( D => n11109, CK => CLK, Q => n53963, 
                           QN => n3822);
   REGS_reg_99_23_inst : DFF_X1 port map( D => n11164, CK => CLK, Q => n53964, 
                           QN => n3823);
   REGS_reg_99_22_inst : DFF_X1 port map( D => n11163, CK => CLK, Q => n53965, 
                           QN => n3824);
   REGS_reg_99_21_inst : DFF_X1 port map( D => n11162, CK => CLK, Q => n53966, 
                           QN => n3825);
   REGS_reg_99_20_inst : DFF_X1 port map( D => n11161, CK => CLK, Q => n53967, 
                           QN => n3826);
   REGS_reg_99_19_inst : DFF_X1 port map( D => n11160, CK => CLK, Q => n53968, 
                           QN => n3827);
   REGS_reg_99_18_inst : DFF_X1 port map( D => n11159, CK => CLK, Q => n53969, 
                           QN => n3828);
   REGS_reg_99_17_inst : DFF_X1 port map( D => n11158, CK => CLK, Q => n53970, 
                           QN => n3829);
   REGS_reg_99_16_inst : DFF_X1 port map( D => n11157, CK => CLK, Q => n53971, 
                           QN => n3830);
   REGS_reg_99_15_inst : DFF_X1 port map( D => n11156, CK => CLK, Q => n53972, 
                           QN => n3831);
   REGS_reg_99_14_inst : DFF_X1 port map( D => n11155, CK => CLK, Q => n53973, 
                           QN => n3832);
   REGS_reg_99_13_inst : DFF_X1 port map( D => n11154, CK => CLK, Q => n53974, 
                           QN => n3833);
   REGS_reg_99_12_inst : DFF_X1 port map( D => n11153, CK => CLK, Q => n53975, 
                           QN => n3834);
   REGS_reg_99_11_inst : DFF_X1 port map( D => n11152, CK => CLK, Q => n53976, 
                           QN => n3835);
   REGS_reg_99_10_inst : DFF_X1 port map( D => n11151, CK => CLK, Q => n53977, 
                           QN => n3836);
   REGS_reg_99_9_inst : DFF_X1 port map( D => n11150, CK => CLK, Q => n53978, 
                           QN => n3837);
   REGS_reg_99_8_inst : DFF_X1 port map( D => n11149, CK => CLK, Q => n53979, 
                           QN => n3838);
   REGS_reg_99_7_inst : DFF_X1 port map( D => n11148, CK => CLK, Q => n53980, 
                           QN => n3839);
   REGS_reg_99_6_inst : DFF_X1 port map( D => n11147, CK => CLK, Q => n53981, 
                           QN => n3840);
   REGS_reg_99_5_inst : DFF_X1 port map( D => n11146, CK => CLK, Q => n53982, 
                           QN => n3841);
   REGS_reg_99_4_inst : DFF_X1 port map( D => n11145, CK => CLK, Q => n53983, 
                           QN => n3842);
   REGS_reg_99_3_inst : DFF_X1 port map( D => n11144, CK => CLK, Q => n53984, 
                           QN => n3843);
   REGS_reg_99_2_inst : DFF_X1 port map( D => n11143, CK => CLK, Q => n53985, 
                           QN => n3844);
   REGS_reg_99_1_inst : DFF_X1 port map( D => n11142, CK => CLK, Q => n53986, 
                           QN => n3845);
   REGS_reg_99_0_inst : DFF_X1 port map( D => n11141, CK => CLK, Q => n53987, 
                           QN => n3846);
   REGS_reg_98_23_inst : DFF_X1 port map( D => n11196, CK => CLK, Q => n3099, 
                           QN => n3847);
   REGS_reg_98_22_inst : DFF_X1 port map( D => n11195, CK => CLK, Q => n3100, 
                           QN => n3848);
   REGS_reg_98_21_inst : DFF_X1 port map( D => n11194, CK => CLK, Q => n3101, 
                           QN => n3849);
   REGS_reg_98_20_inst : DFF_X1 port map( D => n11193, CK => CLK, Q => n3102, 
                           QN => n3850);
   REGS_reg_98_19_inst : DFF_X1 port map( D => n11192, CK => CLK, Q => n3103, 
                           QN => n3851);
   REGS_reg_98_18_inst : DFF_X1 port map( D => n11191, CK => CLK, Q => n3104, 
                           QN => n3852);
   REGS_reg_98_17_inst : DFF_X1 port map( D => n11190, CK => CLK, Q => n3105, 
                           QN => n3853);
   REGS_reg_98_16_inst : DFF_X1 port map( D => n11189, CK => CLK, Q => n3106, 
                           QN => n3854);
   REGS_reg_98_15_inst : DFF_X1 port map( D => n11188, CK => CLK, Q => n3107, 
                           QN => n3855);
   REGS_reg_98_14_inst : DFF_X1 port map( D => n11187, CK => CLK, Q => n3108, 
                           QN => n3856);
   REGS_reg_98_13_inst : DFF_X1 port map( D => n11186, CK => CLK, Q => n3109, 
                           QN => n3857);
   REGS_reg_98_12_inst : DFF_X1 port map( D => n11185, CK => CLK, Q => n3110, 
                           QN => n3858);
   REGS_reg_98_11_inst : DFF_X1 port map( D => n11184, CK => CLK, Q => n3111, 
                           QN => n3859);
   REGS_reg_98_10_inst : DFF_X1 port map( D => n11183, CK => CLK, Q => n3112, 
                           QN => n3860);
   REGS_reg_98_9_inst : DFF_X1 port map( D => n11182, CK => CLK, Q => n3113, QN
                           => n3861);
   REGS_reg_98_8_inst : DFF_X1 port map( D => n11181, CK => CLK, Q => n3114, QN
                           => n3862);
   REGS_reg_98_7_inst : DFF_X1 port map( D => n11180, CK => CLK, Q => n3115, QN
                           => n3863);
   REGS_reg_98_6_inst : DFF_X1 port map( D => n11179, CK => CLK, Q => n3116, QN
                           => n3864);
   REGS_reg_98_5_inst : DFF_X1 port map( D => n11178, CK => CLK, Q => n3117, QN
                           => n3865);
   REGS_reg_98_4_inst : DFF_X1 port map( D => n11177, CK => CLK, Q => n3118, QN
                           => n3866);
   REGS_reg_98_3_inst : DFF_X1 port map( D => n11176, CK => CLK, Q => n3119, QN
                           => n3867);
   REGS_reg_98_2_inst : DFF_X1 port map( D => n11175, CK => CLK, Q => n3120, QN
                           => n3868);
   REGS_reg_98_1_inst : DFF_X1 port map( D => n11174, CK => CLK, Q => n3121, QN
                           => n3869);
   REGS_reg_98_0_inst : DFF_X1 port map( D => n11173, CK => CLK, Q => n3122, QN
                           => n3870);
   REGS_reg_97_23_inst : DFF_X1 port map( D => n11228, CK => CLK, Q => n_1840, 
                           QN => n3871);
   REGS_reg_97_22_inst : DFF_X1 port map( D => n11227, CK => CLK, Q => n_1841, 
                           QN => n3872);
   REGS_reg_97_21_inst : DFF_X1 port map( D => n11226, CK => CLK, Q => n_1842, 
                           QN => n3873);
   REGS_reg_97_20_inst : DFF_X1 port map( D => n11225, CK => CLK, Q => n_1843, 
                           QN => n3874);
   REGS_reg_97_19_inst : DFF_X1 port map( D => n11224, CK => CLK, Q => n_1844, 
                           QN => n3875);
   REGS_reg_97_18_inst : DFF_X1 port map( D => n11223, CK => CLK, Q => n_1845, 
                           QN => n3876);
   REGS_reg_97_17_inst : DFF_X1 port map( D => n11222, CK => CLK, Q => n_1846, 
                           QN => n3877);
   REGS_reg_97_16_inst : DFF_X1 port map( D => n11221, CK => CLK, Q => n_1847, 
                           QN => n3878);
   REGS_reg_97_15_inst : DFF_X1 port map( D => n11220, CK => CLK, Q => n_1848, 
                           QN => n3879);
   REGS_reg_97_14_inst : DFF_X1 port map( D => n11219, CK => CLK, Q => n_1849, 
                           QN => n3880);
   REGS_reg_97_13_inst : DFF_X1 port map( D => n11218, CK => CLK, Q => n_1850, 
                           QN => n3881);
   REGS_reg_97_12_inst : DFF_X1 port map( D => n11217, CK => CLK, Q => n_1851, 
                           QN => n3882);
   REGS_reg_97_11_inst : DFF_X1 port map( D => n11216, CK => CLK, Q => n_1852, 
                           QN => n3883);
   REGS_reg_97_10_inst : DFF_X1 port map( D => n11215, CK => CLK, Q => n_1853, 
                           QN => n3884);
   REGS_reg_97_9_inst : DFF_X1 port map( D => n11214, CK => CLK, Q => n_1854, 
                           QN => n3885);
   REGS_reg_97_8_inst : DFF_X1 port map( D => n11213, CK => CLK, Q => n_1855, 
                           QN => n3886);
   REGS_reg_97_7_inst : DFF_X1 port map( D => n11212, CK => CLK, Q => n_1856, 
                           QN => n3887);
   REGS_reg_97_6_inst : DFF_X1 port map( D => n11211, CK => CLK, Q => n_1857, 
                           QN => n3888);
   REGS_reg_97_5_inst : DFF_X1 port map( D => n11210, CK => CLK, Q => n_1858, 
                           QN => n3889);
   REGS_reg_97_4_inst : DFF_X1 port map( D => n11209, CK => CLK, Q => n_1859, 
                           QN => n3890);
   REGS_reg_97_3_inst : DFF_X1 port map( D => n11208, CK => CLK, Q => n_1860, 
                           QN => n3891);
   REGS_reg_97_2_inst : DFF_X1 port map( D => n11207, CK => CLK, Q => n_1861, 
                           QN => n3892);
   REGS_reg_97_1_inst : DFF_X1 port map( D => n11206, CK => CLK, Q => n_1862, 
                           QN => n3893);
   REGS_reg_97_0_inst : DFF_X1 port map( D => n11205, CK => CLK, Q => n_1863, 
                           QN => n3894);
   REGS_reg_96_23_inst : DFF_X1 port map( D => n11260, CK => CLK, Q => n16106, 
                           QN => n3895);
   REGS_reg_96_22_inst : DFF_X1 port map( D => n11259, CK => CLK, Q => n16104, 
                           QN => n3896);
   REGS_reg_96_21_inst : DFF_X1 port map( D => n11258, CK => CLK, Q => n16102, 
                           QN => n3897);
   REGS_reg_96_20_inst : DFF_X1 port map( D => n11257, CK => CLK, Q => n16100, 
                           QN => n3898);
   REGS_reg_96_19_inst : DFF_X1 port map( D => n11256, CK => CLK, Q => n16118, 
                           QN => n3899);
   REGS_reg_96_18_inst : DFF_X1 port map( D => n11255, CK => CLK, Q => n16116, 
                           QN => n3900);
   REGS_reg_96_17_inst : DFF_X1 port map( D => n11254, CK => CLK, Q => n16114, 
                           QN => n3901);
   REGS_reg_96_16_inst : DFF_X1 port map( D => n11253, CK => CLK, Q => n16112, 
                           QN => n3902);
   REGS_reg_96_15_inst : DFF_X1 port map( D => n11252, CK => CLK, Q => n16110, 
                           QN => n3903);
   REGS_reg_96_14_inst : DFF_X1 port map( D => n11251, CK => CLK, Q => n16122, 
                           QN => n3904);
   REGS_reg_96_13_inst : DFF_X1 port map( D => n11250, CK => CLK, Q => n16120, 
                           QN => n3905);
   REGS_reg_96_12_inst : DFF_X1 port map( D => n11249, CK => CLK, Q => n16108, 
                           QN => n3906);
   REGS_reg_96_11_inst : DFF_X1 port map( D => n11248, CK => CLK, Q => n16136, 
                           QN => n3907);
   REGS_reg_96_10_inst : DFF_X1 port map( D => n11247, CK => CLK, Q => n16134, 
                           QN => n3908);
   REGS_reg_96_9_inst : DFF_X1 port map( D => n11246, CK => CLK, Q => n16132, 
                           QN => n3909);
   REGS_reg_96_8_inst : DFF_X1 port map( D => n11245, CK => CLK, Q => n16128, 
                           QN => n3910);
   REGS_reg_96_7_inst : DFF_X1 port map( D => n11244, CK => CLK, Q => n16130, 
                           QN => n3911);
   REGS_reg_96_6_inst : DFF_X1 port map( D => n11243, CK => CLK, Q => n16126, 
                           QN => n3912);
   REGS_reg_96_5_inst : DFF_X1 port map( D => n11242, CK => CLK, Q => n16124, 
                           QN => n3913);
   REGS_reg_96_4_inst : DFF_X1 port map( D => n11241, CK => CLK, Q => n16139, 
                           QN => n3914);
   REGS_reg_96_3_inst : DFF_X1 port map( D => n11240, CK => CLK, Q => n16138, 
                           QN => n3915);
   REGS_reg_96_2_inst : DFF_X1 port map( D => n11239, CK => CLK, Q => n16142, 
                           QN => n3916);
   REGS_reg_96_1_inst : DFF_X1 port map( D => n11238, CK => CLK, Q => n16141, 
                           QN => n3917);
   REGS_reg_96_0_inst : DFF_X1 port map( D => n11237, CK => CLK, Q => n16140, 
                           QN => n3918);
   REGS_reg_95_23_inst : DFF_X1 port map( D => n11292, CK => CLK, Q => n16107, 
                           QN => n1787);
   REGS_reg_95_22_inst : DFF_X1 port map( D => n11291, CK => CLK, Q => n16105, 
                           QN => n1788);
   REGS_reg_95_21_inst : DFF_X1 port map( D => n11290, CK => CLK, Q => n16103, 
                           QN => n1789);
   REGS_reg_95_20_inst : DFF_X1 port map( D => n11289, CK => CLK, Q => n16101, 
                           QN => n1790);
   REGS_reg_95_19_inst : DFF_X1 port map( D => n11288, CK => CLK, Q => n16119, 
                           QN => n1791);
   REGS_reg_95_18_inst : DFF_X1 port map( D => n11287, CK => CLK, Q => n16117, 
                           QN => n1792);
   REGS_reg_95_17_inst : DFF_X1 port map( D => n11286, CK => CLK, Q => n16115, 
                           QN => n1793);
   REGS_reg_95_16_inst : DFF_X1 port map( D => n11285, CK => CLK, Q => n16113, 
                           QN => n1794);
   REGS_reg_95_15_inst : DFF_X1 port map( D => n11284, CK => CLK, Q => n16111, 
                           QN => n1795);
   REGS_reg_95_14_inst : DFF_X1 port map( D => n11283, CK => CLK, Q => n16123, 
                           QN => n1796);
   REGS_reg_95_13_inst : DFF_X1 port map( D => n11282, CK => CLK, Q => n16121, 
                           QN => n1797);
   REGS_reg_95_12_inst : DFF_X1 port map( D => n11281, CK => CLK, Q => n16109, 
                           QN => n1798);
   REGS_reg_95_11_inst : DFF_X1 port map( D => n11280, CK => CLK, Q => n16137, 
                           QN => n1799);
   REGS_reg_95_10_inst : DFF_X1 port map( D => n11279, CK => CLK, Q => n16135, 
                           QN => n1800);
   REGS_reg_95_9_inst : DFF_X1 port map( D => n11278, CK => CLK, Q => n16133, 
                           QN => n1801);
   REGS_reg_95_8_inst : DFF_X1 port map( D => n11277, CK => CLK, Q => n16129, 
                           QN => n1802);
   REGS_reg_95_7_inst : DFF_X1 port map( D => n11276, CK => CLK, Q => n16131, 
                           QN => n1803);
   REGS_reg_95_6_inst : DFF_X1 port map( D => n11275, CK => CLK, Q => n16127, 
                           QN => n1804);
   REGS_reg_95_5_inst : DFF_X1 port map( D => n11274, CK => CLK, Q => n16125, 
                           QN => n1805);
   REGS_reg_95_4_inst : DFF_X1 port map( D => n11273, CK => CLK, Q => n16481, 
                           QN => n4403);
   REGS_reg_95_3_inst : DFF_X1 port map( D => n11272, CK => CLK, Q => n16480, 
                           QN => n4404);
   REGS_reg_95_2_inst : DFF_X1 port map( D => n11271, CK => CLK, Q => n16479, 
                           QN => n4405);
   REGS_reg_95_1_inst : DFF_X1 port map( D => n11270, CK => CLK, Q => n16478, 
                           QN => n4406);
   REGS_reg_95_0_inst : DFF_X1 port map( D => n11269, CK => CLK, Q => n16477, 
                           QN => n4407);
   REGS_reg_94_16_inst : DFF_X1 port map( D => n11317, CK => CLK, Q => n15723, 
                           QN => n1813);
   REGS_reg_94_15_inst : DFF_X1 port map( D => n11316, CK => CLK, Q => n15722, 
                           QN => n1814);
   REGS_reg_94_14_inst : DFF_X1 port map( D => n11315, CK => CLK, Q => n15721, 
                           QN => n1815);
   REGS_reg_94_13_inst : DFF_X1 port map( D => n11314, CK => CLK, Q => n15720, 
                           QN => n1816);
   REGS_reg_94_12_inst : DFF_X1 port map( D => n11313, CK => CLK, Q => n15719, 
                           QN => n1817);
   REGS_reg_94_11_inst : DFF_X1 port map( D => n11312, CK => CLK, Q => n15718, 
                           QN => n1818);
   REGS_reg_94_10_inst : DFF_X1 port map( D => n11311, CK => CLK, Q => n15717, 
                           QN => n1819);
   REGS_reg_94_9_inst : DFF_X1 port map( D => n11310, CK => CLK, Q => n15716, 
                           QN => n1820);
   REGS_reg_94_8_inst : DFF_X1 port map( D => n11309, CK => CLK, Q => n15715, 
                           QN => n1821);
   REGS_reg_94_7_inst : DFF_X1 port map( D => n11308, CK => CLK, Q => n15714, 
                           QN => n1822);
   REGS_reg_94_6_inst : DFF_X1 port map( D => n11307, CK => CLK, Q => n15713, 
                           QN => n1823);
   REGS_reg_94_5_inst : DFF_X1 port map( D => n11306, CK => CLK, Q => n15712, 
                           QN => n1824);
   REGS_reg_94_4_inst : DFF_X1 port map( D => n11305, CK => CLK, Q => n15711, 
                           QN => n1825);
   REGS_reg_94_3_inst : DFF_X1 port map( D => n11304, CK => CLK, Q => n15710, 
                           QN => n1826);
   REGS_reg_94_2_inst : DFF_X1 port map( D => n11303, CK => CLK, Q => n15709, 
                           QN => n1827);
   REGS_reg_94_1_inst : DFF_X1 port map( D => n11302, CK => CLK, Q => n15708, 
                           QN => n1828);
   REGS_reg_94_0_inst : DFF_X1 port map( D => n11301, CK => CLK, Q => n15707, 
                           QN => n1829);
   REGS_reg_93_23_inst : DFF_X1 port map( D => n11356, CK => CLK, Q => n15538, 
                           QN => n1830);
   REGS_reg_93_22_inst : DFF_X1 port map( D => n11355, CK => CLK, Q => n15537, 
                           QN => n1831);
   REGS_reg_93_21_inst : DFF_X1 port map( D => n11354, CK => CLK, Q => n15536, 
                           QN => n1832);
   REGS_reg_93_20_inst : DFF_X1 port map( D => n11353, CK => CLK, Q => n15535, 
                           QN => n1833);
   REGS_reg_93_19_inst : DFF_X1 port map( D => n11352, CK => CLK, Q => n15534, 
                           QN => n1834);
   REGS_reg_93_18_inst : DFF_X1 port map( D => n11351, CK => CLK, Q => n15533, 
                           QN => n1835);
   REGS_reg_93_17_inst : DFF_X1 port map( D => n11350, CK => CLK, Q => n15532, 
                           QN => n1836);
   REGS_reg_93_16_inst : DFF_X1 port map( D => n11349, CK => CLK, Q => n15531, 
                           QN => n1837);
   REGS_reg_93_15_inst : DFF_X1 port map( D => n11348, CK => CLK, Q => n15530, 
                           QN => n1838);
   REGS_reg_93_14_inst : DFF_X1 port map( D => n11347, CK => CLK, Q => n15529, 
                           QN => n1839);
   REGS_reg_93_13_inst : DFF_X1 port map( D => n11346, CK => CLK, Q => n15528, 
                           QN => n1840);
   REGS_reg_93_12_inst : DFF_X1 port map( D => n11345, CK => CLK, Q => n15527, 
                           QN => n1841);
   REGS_reg_93_11_inst : DFF_X1 port map( D => n11344, CK => CLK, Q => n15526, 
                           QN => n1842);
   REGS_reg_93_10_inst : DFF_X1 port map( D => n11343, CK => CLK, Q => n15525, 
                           QN => n1843);
   REGS_reg_93_9_inst : DFF_X1 port map( D => n11342, CK => CLK, Q => n15524, 
                           QN => n1844);
   REGS_reg_93_8_inst : DFF_X1 port map( D => n11341, CK => CLK, Q => n15523, 
                           QN => n1845);
   REGS_reg_93_7_inst : DFF_X1 port map( D => n11340, CK => CLK, Q => n15522, 
                           QN => n1846);
   REGS_reg_93_6_inst : DFF_X1 port map( D => n11339, CK => CLK, Q => n15521, 
                           QN => n1847);
   REGS_reg_93_5_inst : DFF_X1 port map( D => n11338, CK => CLK, Q => n15520, 
                           QN => n1848);
   REGS_reg_90_23_inst : DFF_X1 port map( D => n11452, CK => CLK, Q => n15871, 
                           QN => n1902);
   REGS_reg_90_22_inst : DFF_X1 port map( D => n11451, CK => CLK, Q => n15866, 
                           QN => n1903);
   REGS_reg_90_21_inst : DFF_X1 port map( D => n11450, CK => CLK, Q => n15861, 
                           QN => n1904);
   REGS_reg_90_20_inst : DFF_X1 port map( D => n11449, CK => CLK, Q => n15856, 
                           QN => n1905);
   REGS_reg_90_19_inst : DFF_X1 port map( D => n11448, CK => CLK, Q => n15851, 
                           QN => n1906);
   REGS_reg_90_18_inst : DFF_X1 port map( D => n11447, CK => CLK, Q => n15798, 
                           QN => n1907);
   REGS_reg_90_17_inst : DFF_X1 port map( D => n11446, CK => CLK, Q => n15793, 
                           QN => n1908);
   REGS_reg_90_16_inst : DFF_X1 port map( D => n11445, CK => CLK, Q => n15788, 
                           QN => n1909);
   REGS_reg_90_15_inst : DFF_X1 port map( D => n11444, CK => CLK, Q => n15783, 
                           QN => n1910);
   REGS_reg_90_14_inst : DFF_X1 port map( D => n11443, CK => CLK, Q => n15778, 
                           QN => n1911);
   REGS_reg_90_13_inst : DFF_X1 port map( D => n11442, CK => CLK, Q => n15773, 
                           QN => n1912);
   REGS_reg_90_12_inst : DFF_X1 port map( D => n11441, CK => CLK, Q => n15768, 
                           QN => n1913);
   REGS_reg_90_11_inst : DFF_X1 port map( D => n11440, CK => CLK, Q => n15763, 
                           QN => n1914);
   REGS_reg_90_10_inst : DFF_X1 port map( D => n11439, CK => CLK, Q => n15758, 
                           QN => n1915);
   REGS_reg_90_9_inst : DFF_X1 port map( D => n11438, CK => CLK, Q => n15753, 
                           QN => n1916);
   REGS_reg_90_8_inst : DFF_X1 port map( D => n11437, CK => CLK, Q => n15748, 
                           QN => n1917);
   REGS_reg_90_7_inst : DFF_X1 port map( D => n11436, CK => CLK, Q => n15909, 
                           QN => n1918);
   REGS_reg_90_6_inst : DFF_X1 port map( D => n11435, CK => CLK, Q => n15904, 
                           QN => n1919);
   REGS_reg_90_5_inst : DFF_X1 port map( D => n11434, CK => CLK, Q => n15899, 
                           QN => n1920);
   REGS_reg_90_4_inst : DFF_X1 port map( D => n11433, CK => CLK, Q => n15894, 
                           QN => n1921);
   REGS_reg_90_3_inst : DFF_X1 port map( D => n11432, CK => CLK, Q => n15889, 
                           QN => n1922);
   REGS_reg_90_2_inst : DFF_X1 port map( D => n11431, CK => CLK, Q => n15886, 
                           QN => n1923);
   REGS_reg_90_1_inst : DFF_X1 port map( D => n11430, CK => CLK, Q => n15881, 
                           QN => n1924);
   REGS_reg_90_0_inst : DFF_X1 port map( D => n11429, CK => CLK, Q => n15876, 
                           QN => n1925);
   REGS_reg_89_23_inst : DFF_X1 port map( D => n11484, CK => CLK, Q => n15872, 
                           QN => n1926);
   REGS_reg_89_22_inst : DFF_X1 port map( D => n11483, CK => CLK, Q => n15867, 
                           QN => n1927);
   REGS_reg_89_21_inst : DFF_X1 port map( D => n11482, CK => CLK, Q => n15862, 
                           QN => n1928);
   REGS_reg_89_20_inst : DFF_X1 port map( D => n11481, CK => CLK, Q => n15857, 
                           QN => n1929);
   REGS_reg_89_19_inst : DFF_X1 port map( D => n11480, CK => CLK, Q => n15852, 
                           QN => n1930);
   REGS_reg_89_18_inst : DFF_X1 port map( D => n11479, CK => CLK, Q => n15799, 
                           QN => n1931);
   REGS_reg_89_17_inst : DFF_X1 port map( D => n11478, CK => CLK, Q => n15794, 
                           QN => n1932);
   REGS_reg_89_16_inst : DFF_X1 port map( D => n11477, CK => CLK, Q => n15789, 
                           QN => n1933);
   REGS_reg_89_15_inst : DFF_X1 port map( D => n11476, CK => CLK, Q => n15784, 
                           QN => n1934);
   REGS_reg_89_14_inst : DFF_X1 port map( D => n11475, CK => CLK, Q => n15779, 
                           QN => n1935);
   REGS_reg_89_13_inst : DFF_X1 port map( D => n11474, CK => CLK, Q => n15774, 
                           QN => n1936);
   REGS_reg_89_12_inst : DFF_X1 port map( D => n11473, CK => CLK, Q => n15769, 
                           QN => n1937);
   REGS_reg_89_11_inst : DFF_X1 port map( D => n11472, CK => CLK, Q => n15764, 
                           QN => n1938);
   REGS_reg_89_10_inst : DFF_X1 port map( D => n11471, CK => CLK, Q => n15759, 
                           QN => n1939);
   REGS_reg_89_9_inst : DFF_X1 port map( D => n11470, CK => CLK, Q => n15754, 
                           QN => n1940);
   REGS_reg_89_8_inst : DFF_X1 port map( D => n11469, CK => CLK, Q => n15749, 
                           QN => n1941);
   REGS_reg_89_7_inst : DFF_X1 port map( D => n11468, CK => CLK, Q => n15910, 
                           QN => n1942);
   REGS_reg_89_6_inst : DFF_X1 port map( D => n11467, CK => CLK, Q => n15905, 
                           QN => n1943);
   REGS_reg_89_5_inst : DFF_X1 port map( D => n11466, CK => CLK, Q => n15900, 
                           QN => n1944);
   REGS_reg_89_4_inst : DFF_X1 port map( D => n11465, CK => CLK, Q => n15895, 
                           QN => n1945);
   REGS_reg_89_3_inst : DFF_X1 port map( D => n11464, CK => CLK, Q => n15890, 
                           QN => n1946);
   REGS_reg_89_2_inst : DFF_X1 port map( D => n11463, CK => CLK, Q => n15887, 
                           QN => n1947);
   REGS_reg_89_1_inst : DFF_X1 port map( D => n11462, CK => CLK, Q => n15882, 
                           QN => n1948);
   REGS_reg_89_0_inst : DFF_X1 port map( D => n11461, CK => CLK, Q => n15877, 
                           QN => n1949);
   REGS_reg_88_23_inst : DFF_X1 port map( D => n11516, CK => CLK, Q => n15873, 
                           QN => n1950);
   REGS_reg_88_22_inst : DFF_X1 port map( D => n11515, CK => CLK, Q => n15868, 
                           QN => n1951);
   REGS_reg_88_21_inst : DFF_X1 port map( D => n11514, CK => CLK, Q => n15863, 
                           QN => n1952);
   REGS_reg_88_20_inst : DFF_X1 port map( D => n11513, CK => CLK, Q => n15858, 
                           QN => n1953);
   REGS_reg_88_19_inst : DFF_X1 port map( D => n11512, CK => CLK, Q => n15853, 
                           QN => n1954);
   REGS_reg_88_18_inst : DFF_X1 port map( D => n11511, CK => CLK, Q => n15800, 
                           QN => n1955);
   REGS_reg_88_17_inst : DFF_X1 port map( D => n11510, CK => CLK, Q => n15795, 
                           QN => n1956);
   REGS_reg_88_16_inst : DFF_X1 port map( D => n11509, CK => CLK, Q => n15790, 
                           QN => n1957);
   REGS_reg_88_15_inst : DFF_X1 port map( D => n11508, CK => CLK, Q => n15785, 
                           QN => n1958);
   REGS_reg_88_14_inst : DFF_X1 port map( D => n11507, CK => CLK, Q => n15780, 
                           QN => n1959);
   REGS_reg_88_13_inst : DFF_X1 port map( D => n11506, CK => CLK, Q => n15775, 
                           QN => n1960);
   REGS_reg_88_12_inst : DFF_X1 port map( D => n11505, CK => CLK, Q => n15770, 
                           QN => n1961);
   REGS_reg_88_11_inst : DFF_X1 port map( D => n11504, CK => CLK, Q => n15765, 
                           QN => n1962);
   REGS_reg_88_10_inst : DFF_X1 port map( D => n11503, CK => CLK, Q => n15760, 
                           QN => n1963);
   REGS_reg_88_9_inst : DFF_X1 port map( D => n11502, CK => CLK, Q => n15755, 
                           QN => n1964);
   REGS_reg_88_8_inst : DFF_X1 port map( D => n11501, CK => CLK, Q => n15750, 
                           QN => n1965);
   REGS_reg_88_7_inst : DFF_X1 port map( D => n11500, CK => CLK, Q => n15911, 
                           QN => n1966);
   REGS_reg_88_6_inst : DFF_X1 port map( D => n11499, CK => CLK, Q => n15906, 
                           QN => n1967);
   REGS_reg_88_5_inst : DFF_X1 port map( D => n11498, CK => CLK, Q => n15901, 
                           QN => n1968);
   REGS_reg_88_4_inst : DFF_X1 port map( D => n11497, CK => CLK, Q => n15896, 
                           QN => n1969);
   REGS_reg_88_3_inst : DFF_X1 port map( D => n11496, CK => CLK, Q => n15891, 
                           QN => n1970);
   REGS_reg_88_2_inst : DFF_X1 port map( D => n11495, CK => CLK, Q => n15888, 
                           QN => n1971);
   REGS_reg_88_1_inst : DFF_X1 port map( D => n11494, CK => CLK, Q => n15883, 
                           QN => n1972);
   REGS_reg_88_0_inst : DFF_X1 port map( D => n11493, CK => CLK, Q => n15878, 
                           QN => n1973);
   REGS_reg_87_23_inst : DFF_X1 port map( D => n11548, CK => CLK, Q => n16553, 
                           QN => n4408);
   REGS_reg_87_22_inst : DFF_X1 port map( D => n11547, CK => CLK, Q => n16552, 
                           QN => n4409);
   REGS_reg_87_21_inst : DFF_X1 port map( D => n11546, CK => CLK, Q => n16551, 
                           QN => n4410);
   REGS_reg_87_20_inst : DFF_X1 port map( D => n11545, CK => CLK, Q => n16550, 
                           QN => n4411);
   REGS_reg_87_19_inst : DFF_X1 port map( D => n11544, CK => CLK, Q => n16549, 
                           QN => n4412);
   REGS_reg_87_18_inst : DFF_X1 port map( D => n11543, CK => CLK, Q => n16548, 
                           QN => n4413);
   REGS_reg_87_17_inst : DFF_X1 port map( D => n11542, CK => CLK, Q => n16547, 
                           QN => n4414);
   REGS_reg_87_16_inst : DFF_X1 port map( D => n11541, CK => CLK, Q => n16546, 
                           QN => n4415);
   REGS_reg_87_15_inst : DFF_X1 port map( D => n11540, CK => CLK, Q => n16545, 
                           QN => n4416);
   REGS_reg_87_14_inst : DFF_X1 port map( D => n11539, CK => CLK, Q => n16544, 
                           QN => n4417);
   REGS_reg_87_13_inst : DFF_X1 port map( D => n11538, CK => CLK, Q => n16543, 
                           QN => n4418);
   REGS_reg_87_12_inst : DFF_X1 port map( D => n11537, CK => CLK, Q => n16542, 
                           QN => n4419);
   REGS_reg_87_11_inst : DFF_X1 port map( D => n11536, CK => CLK, Q => n16541, 
                           QN => n4420);
   REGS_reg_87_10_inst : DFF_X1 port map( D => n11535, CK => CLK, Q => n16540, 
                           QN => n4421);
   REGS_reg_87_9_inst : DFF_X1 port map( D => n11534, CK => CLK, Q => n16539, 
                           QN => n4422);
   REGS_reg_87_8_inst : DFF_X1 port map( D => n11533, CK => CLK, Q => n16538, 
                           QN => n4423);
   REGS_reg_87_7_inst : DFF_X1 port map( D => n11532, CK => CLK, Q => n16537, 
                           QN => n4424);
   REGS_reg_87_6_inst : DFF_X1 port map( D => n11531, CK => CLK, Q => n16536, 
                           QN => n4425);
   REGS_reg_87_5_inst : DFF_X1 port map( D => n11530, CK => CLK, Q => n16535, 
                           QN => n4426);
   REGS_reg_87_4_inst : DFF_X1 port map( D => n11529, CK => CLK, Q => n16534, 
                           QN => n4427);
   REGS_reg_87_3_inst : DFF_X1 port map( D => n11528, CK => CLK, Q => n16533, 
                           QN => n4428);
   REGS_reg_87_2_inst : DFF_X1 port map( D => n11527, CK => CLK, Q => n16532, 
                           QN => n4429);
   REGS_reg_87_1_inst : DFF_X1 port map( D => n11526, CK => CLK, Q => n16531, 
                           QN => n4430);
   REGS_reg_87_0_inst : DFF_X1 port map( D => n11525, CK => CLK, Q => n16530, 
                           QN => n4431);
   REGS_reg_86_23_inst : DFF_X1 port map( D => n11580, CK => CLK, Q => n_1864, 
                           QN => n1974);
   REGS_reg_86_22_inst : DFF_X1 port map( D => n11579, CK => CLK, Q => n_1865, 
                           QN => n1975);
   REGS_reg_86_21_inst : DFF_X1 port map( D => n11578, CK => CLK, Q => n_1866, 
                           QN => n1976);
   REGS_reg_86_20_inst : DFF_X1 port map( D => n11577, CK => CLK, Q => n_1867, 
                           QN => n1977);
   REGS_reg_86_19_inst : DFF_X1 port map( D => n11576, CK => CLK, Q => n_1868, 
                           QN => n1978);
   REGS_reg_86_18_inst : DFF_X1 port map( D => n11575, CK => CLK, Q => n_1869, 
                           QN => n1979);
   REGS_reg_86_17_inst : DFF_X1 port map( D => n11574, CK => CLK, Q => n_1870, 
                           QN => n1980);
   REGS_reg_86_16_inst : DFF_X1 port map( D => n11573, CK => CLK, Q => n_1871, 
                           QN => n1981);
   REGS_reg_86_15_inst : DFF_X1 port map( D => n11572, CK => CLK, Q => n_1872, 
                           QN => n1982);
   REGS_reg_86_14_inst : DFF_X1 port map( D => n11571, CK => CLK, Q => n_1873, 
                           QN => n1983);
   REGS_reg_86_13_inst : DFF_X1 port map( D => n11570, CK => CLK, Q => n_1874, 
                           QN => n1984);
   REGS_reg_86_12_inst : DFF_X1 port map( D => n11569, CK => CLK, Q => n_1875, 
                           QN => n1985);
   REGS_reg_86_11_inst : DFF_X1 port map( D => n11568, CK => CLK, Q => n_1876, 
                           QN => n1986);
   REGS_reg_86_10_inst : DFF_X1 port map( D => n11567, CK => CLK, Q => n_1877, 
                           QN => n1987);
   REGS_reg_86_9_inst : DFF_X1 port map( D => n11566, CK => CLK, Q => n_1878, 
                           QN => n1988);
   REGS_reg_86_8_inst : DFF_X1 port map( D => n11565, CK => CLK, Q => n_1879, 
                           QN => n1989);
   REGS_reg_86_7_inst : DFF_X1 port map( D => n11564, CK => CLK, Q => n_1880, 
                           QN => n1990);
   REGS_reg_86_6_inst : DFF_X1 port map( D => n11563, CK => CLK, Q => n_1881, 
                           QN => n1991);
   REGS_reg_86_5_inst : DFF_X1 port map( D => n11562, CK => CLK, Q => n_1882, 
                           QN => n1992);
   REGS_reg_86_4_inst : DFF_X1 port map( D => n11561, CK => CLK, Q => n_1883, 
                           QN => n1993);
   REGS_reg_86_3_inst : DFF_X1 port map( D => n11560, CK => CLK, Q => n_1884, 
                           QN => n1994);
   REGS_reg_86_2_inst : DFF_X1 port map( D => n11559, CK => CLK, Q => n_1885, 
                           QN => n1995);
   REGS_reg_86_1_inst : DFF_X1 port map( D => n11558, CK => CLK, Q => n_1886, 
                           QN => n1996);
   REGS_reg_86_0_inst : DFF_X1 port map( D => n11557, CK => CLK, Q => n_1887, 
                           QN => n1997);
   REGS_reg_85_23_inst : DFF_X1 port map( D => n11612, CK => CLK, Q => n_1888, 
                           QN => n1998);
   REGS_reg_85_22_inst : DFF_X1 port map( D => n11611, CK => CLK, Q => n_1889, 
                           QN => n2023);
   REGS_reg_85_21_inst : DFF_X1 port map( D => n11610, CK => CLK, Q => n_1890, 
                           QN => n2024);
   REGS_reg_85_20_inst : DFF_X1 port map( D => n11609, CK => CLK, Q => n_1891, 
                           QN => n2025);
   REGS_reg_85_19_inst : DFF_X1 port map( D => n11608, CK => CLK, Q => n_1892, 
                           QN => n2026);
   REGS_reg_85_18_inst : DFF_X1 port map( D => n11607, CK => CLK, Q => n_1893, 
                           QN => n2027);
   REGS_reg_85_17_inst : DFF_X1 port map( D => n11606, CK => CLK, Q => n_1894, 
                           QN => n2028);
   REGS_reg_85_16_inst : DFF_X1 port map( D => n11605, CK => CLK, Q => n_1895, 
                           QN => n2029);
   REGS_reg_85_15_inst : DFF_X1 port map( D => n11604, CK => CLK, Q => n_1896, 
                           QN => n2030);
   REGS_reg_85_14_inst : DFF_X1 port map( D => n11603, CK => CLK, Q => n_1897, 
                           QN => n2031);
   REGS_reg_85_13_inst : DFF_X1 port map( D => n11602, CK => CLK, Q => n_1898, 
                           QN => n2032);
   REGS_reg_85_12_inst : DFF_X1 port map( D => n11601, CK => CLK, Q => n_1899, 
                           QN => n2033);
   REGS_reg_85_11_inst : DFF_X1 port map( D => n11600, CK => CLK, Q => n_1900, 
                           QN => n2034);
   REGS_reg_85_10_inst : DFF_X1 port map( D => n11599, CK => CLK, Q => n_1901, 
                           QN => n2035);
   REGS_reg_85_9_inst : DFF_X1 port map( D => n11598, CK => CLK, Q => n_1902, 
                           QN => n2036);
   REGS_reg_85_8_inst : DFF_X1 port map( D => n11597, CK => CLK, Q => n_1903, 
                           QN => n2037);
   REGS_reg_85_7_inst : DFF_X1 port map( D => n11596, CK => CLK, Q => n_1904, 
                           QN => n2038);
   REGS_reg_85_6_inst : DFF_X1 port map( D => n11595, CK => CLK, Q => n_1905, 
                           QN => n2039);
   REGS_reg_85_5_inst : DFF_X1 port map( D => n11594, CK => CLK, Q => n_1906, 
                           QN => n2040);
   REGS_reg_85_4_inst : DFF_X1 port map( D => n11593, CK => CLK, Q => n_1907, 
                           QN => n2041);
   REGS_reg_85_3_inst : DFF_X1 port map( D => n11592, CK => CLK, Q => n_1908, 
                           QN => n2042);
   REGS_reg_85_2_inst : DFF_X1 port map( D => n11591, CK => CLK, Q => n_1909, 
                           QN => n2043);
   REGS_reg_85_1_inst : DFF_X1 port map( D => n11590, CK => CLK, Q => n_1910, 
                           QN => n2044);
   REGS_reg_85_0_inst : DFF_X1 port map( D => n11589, CK => CLK, Q => n_1911, 
                           QN => n2045);
   REGS_reg_84_23_inst : DFF_X1 port map( D => n11644, CK => CLK, Q => n54156, 
                           QN => n2046);
   REGS_reg_84_22_inst : DFF_X1 port map( D => n11643, CK => CLK, Q => n54157, 
                           QN => n2047);
   REGS_reg_84_21_inst : DFF_X1 port map( D => n11642, CK => CLK, Q => n54158, 
                           QN => n2048);
   REGS_reg_84_20_inst : DFF_X1 port map( D => n11641, CK => CLK, Q => n54159, 
                           QN => n2049);
   REGS_reg_84_19_inst : DFF_X1 port map( D => n11640, CK => CLK, Q => n54160, 
                           QN => n2050);
   REGS_reg_84_18_inst : DFF_X1 port map( D => n11639, CK => CLK, Q => n54161, 
                           QN => n2051);
   REGS_reg_84_17_inst : DFF_X1 port map( D => n11638, CK => CLK, Q => n54162, 
                           QN => n2052);
   REGS_reg_84_16_inst : DFF_X1 port map( D => n11637, CK => CLK, Q => n54163, 
                           QN => n2053);
   REGS_reg_84_15_inst : DFF_X1 port map( D => n11636, CK => CLK, Q => n54164, 
                           QN => n2054);
   REGS_reg_84_14_inst : DFF_X1 port map( D => n11635, CK => CLK, Q => n54165, 
                           QN => n2055);
   REGS_reg_84_13_inst : DFF_X1 port map( D => n11634, CK => CLK, Q => n54166, 
                           QN => n2056);
   REGS_reg_84_12_inst : DFF_X1 port map( D => n11633, CK => CLK, Q => n54167, 
                           QN => n2057);
   REGS_reg_84_11_inst : DFF_X1 port map( D => n11632, CK => CLK, Q => n54168, 
                           QN => n2058);
   REGS_reg_84_10_inst : DFF_X1 port map( D => n11631, CK => CLK, Q => n54169, 
                           QN => n2059);
   REGS_reg_84_9_inst : DFF_X1 port map( D => n11630, CK => CLK, Q => n54170, 
                           QN => n2060);
   REGS_reg_84_8_inst : DFF_X1 port map( D => n11629, CK => CLK, Q => n54171, 
                           QN => n2061);
   REGS_reg_84_7_inst : DFF_X1 port map( D => n11628, CK => CLK, Q => n54172, 
                           QN => n2062);
   REGS_reg_84_6_inst : DFF_X1 port map( D => n11627, CK => CLK, Q => n54173, 
                           QN => n2063);
   REGS_reg_84_5_inst : DFF_X1 port map( D => n11626, CK => CLK, Q => n54174, 
                           QN => n2064);
   REGS_reg_84_4_inst : DFF_X1 port map( D => n11625, CK => CLK, Q => n54175, 
                           QN => n2065);
   REGS_reg_84_3_inst : DFF_X1 port map( D => n11624, CK => CLK, Q => n54176, 
                           QN => n2066);
   REGS_reg_84_2_inst : DFF_X1 port map( D => n11623, CK => CLK, Q => n54177, 
                           QN => n2067);
   REGS_reg_84_1_inst : DFF_X1 port map( D => n11622, CK => CLK, Q => n54178, 
                           QN => n2068);
   REGS_reg_84_0_inst : DFF_X1 port map( D => n11621, CK => CLK, Q => n54179, 
                           QN => n2069);
   REGS_reg_83_23_inst : DFF_X1 port map( D => n11676, CK => CLK, Q => n54180, 
                           QN => n2070);
   REGS_reg_83_22_inst : DFF_X1 port map( D => n11675, CK => CLK, Q => n54181, 
                           QN => n2071);
   REGS_reg_83_21_inst : DFF_X1 port map( D => n11674, CK => CLK, Q => n54182, 
                           QN => n2072);
   REGS_reg_83_20_inst : DFF_X1 port map( D => n11673, CK => CLK, Q => n54183, 
                           QN => n2073);
   REGS_reg_83_19_inst : DFF_X1 port map( D => n11672, CK => CLK, Q => n54184, 
                           QN => n2074);
   REGS_reg_83_18_inst : DFF_X1 port map( D => n11671, CK => CLK, Q => n54185, 
                           QN => n2079);
   REGS_reg_83_17_inst : DFF_X1 port map( D => n11670, CK => CLK, Q => n54186, 
                           QN => n2080);
   REGS_reg_83_16_inst : DFF_X1 port map( D => n11669, CK => CLK, Q => n54187, 
                           QN => n2081);
   REGS_reg_83_15_inst : DFF_X1 port map( D => n11668, CK => CLK, Q => n54188, 
                           QN => n2082);
   REGS_reg_83_14_inst : DFF_X1 port map( D => n11667, CK => CLK, Q => n54189, 
                           QN => n2083);
   REGS_reg_83_13_inst : DFF_X1 port map( D => n11666, CK => CLK, Q => n54190, 
                           QN => n2084);
   REGS_reg_83_12_inst : DFF_X1 port map( D => n11665, CK => CLK, Q => n54191, 
                           QN => n2085);
   REGS_reg_83_11_inst : DFF_X1 port map( D => n11664, CK => CLK, Q => n54192, 
                           QN => n2086);
   REGS_reg_83_10_inst : DFF_X1 port map( D => n11663, CK => CLK, Q => n54193, 
                           QN => n2087);
   REGS_reg_83_9_inst : DFF_X1 port map( D => n11662, CK => CLK, Q => n54194, 
                           QN => n2088);
   REGS_reg_83_8_inst : DFF_X1 port map( D => n11661, CK => CLK, Q => n54195, 
                           QN => n2089);
   REGS_reg_83_7_inst : DFF_X1 port map( D => n11660, CK => CLK, Q => n54196, 
                           QN => n2090);
   REGS_reg_83_6_inst : DFF_X1 port map( D => n11659, CK => CLK, Q => n54197, 
                           QN => n2091);
   REGS_reg_83_5_inst : DFF_X1 port map( D => n11658, CK => CLK, Q => n54198, 
                           QN => n2092);
   REGS_reg_83_4_inst : DFF_X1 port map( D => n11657, CK => CLK, Q => n54199, 
                           QN => n2093);
   REGS_reg_83_3_inst : DFF_X1 port map( D => n11656, CK => CLK, Q => n54200, 
                           QN => n2094);
   REGS_reg_83_2_inst : DFF_X1 port map( D => n11655, CK => CLK, Q => n54201, 
                           QN => n2095);
   REGS_reg_83_1_inst : DFF_X1 port map( D => n11654, CK => CLK, Q => n54202, 
                           QN => n2096);
   REGS_reg_83_0_inst : DFF_X1 port map( D => n11653, CK => CLK, Q => n54203, 
                           QN => n2097);
   REGS_reg_82_23_inst : DFF_X1 port map( D => n11708, CK => CLK, Q => n54204, 
                           QN => n2098);
   REGS_reg_82_22_inst : DFF_X1 port map( D => n11707, CK => CLK, Q => n54205, 
                           QN => n2099);
   REGS_reg_82_21_inst : DFF_X1 port map( D => n11706, CK => CLK, Q => n54206, 
                           QN => n2100);
   REGS_reg_82_20_inst : DFF_X1 port map( D => n11705, CK => CLK, Q => n54207, 
                           QN => n2101);
   REGS_reg_82_19_inst : DFF_X1 port map( D => n11704, CK => CLK, Q => n54208, 
                           QN => n2102);
   REGS_reg_82_18_inst : DFF_X1 port map( D => n11703, CK => CLK, Q => n54209, 
                           QN => n2103);
   REGS_reg_82_17_inst : DFF_X1 port map( D => n11702, CK => CLK, Q => n54210, 
                           QN => n2104);
   REGS_reg_82_16_inst : DFF_X1 port map( D => n11701, CK => CLK, Q => n54211, 
                           QN => n2105);
   REGS_reg_82_15_inst : DFF_X1 port map( D => n11700, CK => CLK, Q => n54212, 
                           QN => n2106);
   REGS_reg_82_14_inst : DFF_X1 port map( D => n11699, CK => CLK, Q => n54213, 
                           QN => n2107);
   REGS_reg_82_13_inst : DFF_X1 port map( D => n11698, CK => CLK, Q => n54214, 
                           QN => n2108);
   REGS_reg_82_12_inst : DFF_X1 port map( D => n11697, CK => CLK, Q => n54215, 
                           QN => n2109);
   REGS_reg_82_11_inst : DFF_X1 port map( D => n11696, CK => CLK, Q => n54216, 
                           QN => n2110);
   REGS_reg_82_10_inst : DFF_X1 port map( D => n11695, CK => CLK, Q => n54217, 
                           QN => n2111);
   REGS_reg_82_9_inst : DFF_X1 port map( D => n11694, CK => CLK, Q => n54218, 
                           QN => n2112);
   REGS_reg_82_8_inst : DFF_X1 port map( D => n11693, CK => CLK, Q => n54219, 
                           QN => n2113);
   REGS_reg_82_7_inst : DFF_X1 port map( D => n11692, CK => CLK, Q => n54220, 
                           QN => n2114);
   REGS_reg_82_6_inst : DFF_X1 port map( D => n11691, CK => CLK, Q => n54221, 
                           QN => n2115);
   REGS_reg_82_5_inst : DFF_X1 port map( D => n11690, CK => CLK, Q => n54222, 
                           QN => n2116);
   REGS_reg_82_4_inst : DFF_X1 port map( D => n11689, CK => CLK, Q => n54223, 
                           QN => n2117);
   REGS_reg_82_3_inst : DFF_X1 port map( D => n11688, CK => CLK, Q => n54224, 
                           QN => n2118);
   REGS_reg_82_2_inst : DFF_X1 port map( D => n11687, CK => CLK, Q => n54225, 
                           QN => n2119);
   REGS_reg_82_1_inst : DFF_X1 port map( D => n11686, CK => CLK, Q => n54226, 
                           QN => n2120);
   REGS_reg_82_0_inst : DFF_X1 port map( D => n11685, CK => CLK, Q => n54227, 
                           QN => n2121);
   REGS_reg_81_23_inst : DFF_X1 port map( D => n11740, CK => CLK, Q => n54521, 
                           QN => n2122);
   REGS_reg_81_22_inst : DFF_X1 port map( D => n11739, CK => CLK, Q => n54520, 
                           QN => n2123);
   REGS_reg_81_21_inst : DFF_X1 port map( D => n11738, CK => CLK, Q => n54519, 
                           QN => n2124);
   REGS_reg_81_20_inst : DFF_X1 port map( D => n11737, CK => CLK, Q => n54518, 
                           QN => n2125);
   REGS_reg_81_19_inst : DFF_X1 port map( D => n11736, CK => CLK, Q => n54517, 
                           QN => n2126);
   REGS_reg_81_18_inst : DFF_X1 port map( D => n11735, CK => CLK, Q => n54516, 
                           QN => n2127);
   REGS_reg_81_17_inst : DFF_X1 port map( D => n11734, CK => CLK, Q => n54515, 
                           QN => n2128);
   REGS_reg_81_16_inst : DFF_X1 port map( D => n11733, CK => CLK, Q => n54514, 
                           QN => n2129);
   REGS_reg_81_15_inst : DFF_X1 port map( D => n11732, CK => CLK, Q => n54513, 
                           QN => n2130);
   REGS_reg_81_14_inst : DFF_X1 port map( D => n11731, CK => CLK, Q => n54512, 
                           QN => n2131);
   REGS_reg_81_13_inst : DFF_X1 port map( D => n11730, CK => CLK, Q => n54511, 
                           QN => n2132);
   REGS_reg_81_12_inst : DFF_X1 port map( D => n11729, CK => CLK, Q => n54526, 
                           QN => n2133);
   REGS_reg_81_11_inst : DFF_X1 port map( D => n11728, CK => CLK, Q => n54525, 
                           QN => n2134);
   REGS_reg_81_10_inst : DFF_X1 port map( D => n11727, CK => CLK, Q => n54524, 
                           QN => n2135);
   REGS_reg_81_9_inst : DFF_X1 port map( D => n11726, CK => CLK, Q => n54523, 
                           QN => n2136);
   REGS_reg_81_8_inst : DFF_X1 port map( D => n11725, CK => CLK, Q => n54508, 
                           QN => n2137);
   REGS_reg_81_7_inst : DFF_X1 port map( D => n11724, CK => CLK, Q => n54522, 
                           QN => n2138);
   REGS_reg_81_6_inst : DFF_X1 port map( D => n11723, CK => CLK, Q => n54510, 
                           QN => n2139);
   REGS_reg_81_5_inst : DFF_X1 port map( D => n11722, CK => CLK, Q => n54509, 
                           QN => n2140);
   REGS_reg_81_4_inst : DFF_X1 port map( D => n11721, CK => CLK, Q => n54507, 
                           QN => n2141);
   REGS_reg_81_3_inst : DFF_X1 port map( D => n11720, CK => CLK, Q => n54506, 
                           QN => n2142);
   REGS_reg_81_2_inst : DFF_X1 port map( D => n11719, CK => CLK, Q => n54505, 
                           QN => n2143);
   REGS_reg_81_1_inst : DFF_X1 port map( D => n11718, CK => CLK, Q => n54504, 
                           QN => n2144);
   REGS_reg_81_0_inst : DFF_X1 port map( D => n11717, CK => CLK, Q => n54527, 
                           QN => n2145);
   REGS_reg_80_23_inst : DFF_X1 port map( D => n11772, CK => CLK, Q => n_1912, 
                           QN => n2146);
   REGS_reg_80_22_inst : DFF_X1 port map( D => n11771, CK => CLK, Q => n_1913, 
                           QN => n2147);
   REGS_reg_80_21_inst : DFF_X1 port map( D => n11770, CK => CLK, Q => n_1914, 
                           QN => n2148);
   REGS_reg_80_20_inst : DFF_X1 port map( D => n11769, CK => CLK, Q => n_1915, 
                           QN => n2149);
   REGS_reg_80_19_inst : DFF_X1 port map( D => n11768, CK => CLK, Q => n_1916, 
                           QN => n2150);
   REGS_reg_80_18_inst : DFF_X1 port map( D => n11767, CK => CLK, Q => n_1917, 
                           QN => n2151);
   REGS_reg_80_17_inst : DFF_X1 port map( D => n11766, CK => CLK, Q => n_1918, 
                           QN => n2152);
   REGS_reg_80_16_inst : DFF_X1 port map( D => n11765, CK => CLK, Q => n_1919, 
                           QN => n2153);
   REGS_reg_80_15_inst : DFF_X1 port map( D => n11764, CK => CLK, Q => n_1920, 
                           QN => n2154);
   REGS_reg_80_14_inst : DFF_X1 port map( D => n11763, CK => CLK, Q => n_1921, 
                           QN => n2155);
   REGS_reg_80_13_inst : DFF_X1 port map( D => n11762, CK => CLK, Q => n_1922, 
                           QN => n2156);
   REGS_reg_80_12_inst : DFF_X1 port map( D => n11761, CK => CLK, Q => n_1923, 
                           QN => n2157);
   REGS_reg_80_11_inst : DFF_X1 port map( D => n11760, CK => CLK, Q => n_1924, 
                           QN => n2158);
   REGS_reg_80_10_inst : DFF_X1 port map( D => n11759, CK => CLK, Q => n_1925, 
                           QN => n2159);
   REGS_reg_80_9_inst : DFF_X1 port map( D => n11758, CK => CLK, Q => n_1926, 
                           QN => n2160);
   REGS_reg_80_8_inst : DFF_X1 port map( D => n11757, CK => CLK, Q => n_1927, 
                           QN => n2161);
   REGS_reg_80_7_inst : DFF_X1 port map( D => n11756, CK => CLK, Q => n_1928, 
                           QN => n2162);
   REGS_reg_80_6_inst : DFF_X1 port map( D => n11755, CK => CLK, Q => n_1929, 
                           QN => n2163);
   REGS_reg_80_5_inst : DFF_X1 port map( D => n11754, CK => CLK, Q => n_1930, 
                           QN => n2164);
   REGS_reg_80_4_inst : DFF_X1 port map( D => n11753, CK => CLK, Q => n_1931, 
                           QN => n2165);
   REGS_reg_80_3_inst : DFF_X1 port map( D => n11752, CK => CLK, Q => n_1932, 
                           QN => n2166);
   REGS_reg_80_2_inst : DFF_X1 port map( D => n11751, CK => CLK, Q => n_1933, 
                           QN => n2167);
   REGS_reg_80_1_inst : DFF_X1 port map( D => n11750, CK => CLK, Q => n_1934, 
                           QN => n2168);
   REGS_reg_80_0_inst : DFF_X1 port map( D => n11749, CK => CLK, Q => n_1935, 
                           QN => n2169);
   REGS_reg_79_23_inst : DFF_X1 port map( D => n11804, CK => CLK, Q => n54228, 
                           QN => n2170);
   REGS_reg_79_22_inst : DFF_X1 port map( D => n11803, CK => CLK, Q => n54229, 
                           QN => n2171);
   REGS_reg_79_21_inst : DFF_X1 port map( D => n11802, CK => CLK, Q => n54230, 
                           QN => n2172);
   REGS_reg_79_20_inst : DFF_X1 port map( D => n11801, CK => CLK, Q => n54231, 
                           QN => n2173);
   REGS_reg_79_19_inst : DFF_X1 port map( D => n11800, CK => CLK, Q => n54232, 
                           QN => n2174);
   REGS_reg_79_18_inst : DFF_X1 port map( D => n11799, CK => CLK, Q => n54233, 
                           QN => n2175);
   REGS_reg_79_17_inst : DFF_X1 port map( D => n11798, CK => CLK, Q => n54234, 
                           QN => n2176);
   REGS_reg_79_16_inst : DFF_X1 port map( D => n11797, CK => CLK, Q => n54235, 
                           QN => n2177);
   REGS_reg_79_15_inst : DFF_X1 port map( D => n11796, CK => CLK, Q => n54236, 
                           QN => n2178);
   REGS_reg_79_14_inst : DFF_X1 port map( D => n11795, CK => CLK, Q => n54237, 
                           QN => n2179);
   REGS_reg_79_13_inst : DFF_X1 port map( D => n11794, CK => CLK, Q => n54238, 
                           QN => n2180);
   REGS_reg_79_12_inst : DFF_X1 port map( D => n11793, CK => CLK, Q => n54239, 
                           QN => n2181);
   REGS_reg_79_11_inst : DFF_X1 port map( D => n11792, CK => CLK, Q => n54240, 
                           QN => n2182);
   REGS_reg_79_10_inst : DFF_X1 port map( D => n11791, CK => CLK, Q => n54241, 
                           QN => n2183);
   REGS_reg_79_9_inst : DFF_X1 port map( D => n11790, CK => CLK, Q => n54242, 
                           QN => n2184);
   REGS_reg_79_8_inst : DFF_X1 port map( D => n11789, CK => CLK, Q => n54243, 
                           QN => n2185);
   REGS_reg_79_7_inst : DFF_X1 port map( D => n11788, CK => CLK, Q => n54244, 
                           QN => n2186);
   REGS_reg_79_6_inst : DFF_X1 port map( D => n11787, CK => CLK, Q => n54245, 
                           QN => n2187);
   REGS_reg_79_5_inst : DFF_X1 port map( D => n11786, CK => CLK, Q => n54246, 
                           QN => n2188);
   REGS_reg_79_4_inst : DFF_X1 port map( D => n11785, CK => CLK, Q => n54247, 
                           QN => n2189);
   REGS_reg_79_3_inst : DFF_X1 port map( D => n11784, CK => CLK, Q => n54248, 
                           QN => n2190);
   REGS_reg_79_2_inst : DFF_X1 port map( D => n11783, CK => CLK, Q => n54249, 
                           QN => n2191);
   REGS_reg_79_1_inst : DFF_X1 port map( D => n11782, CK => CLK, Q => n54250, 
                           QN => n2192);
   REGS_reg_79_0_inst : DFF_X1 port map( D => n11781, CK => CLK, Q => n54251, 
                           QN => n2193);
   REGS_reg_78_23_inst : DFF_X1 port map( D => n11836, CK => CLK, Q => n54252, 
                           QN => n2194);
   REGS_reg_78_22_inst : DFF_X1 port map( D => n11835, CK => CLK, Q => n54253, 
                           QN => n2195);
   REGS_reg_78_21_inst : DFF_X1 port map( D => n11834, CK => CLK, Q => n54254, 
                           QN => n2196);
   REGS_reg_78_20_inst : DFF_X1 port map( D => n11833, CK => CLK, Q => n54255, 
                           QN => n2197);
   REGS_reg_78_19_inst : DFF_X1 port map( D => n11832, CK => CLK, Q => n54256, 
                           QN => n2198);
   REGS_reg_78_18_inst : DFF_X1 port map( D => n11831, CK => CLK, Q => n54257, 
                           QN => n2199);
   REGS_reg_78_17_inst : DFF_X1 port map( D => n11830, CK => CLK, Q => n54258, 
                           QN => n2200);
   REGS_reg_78_16_inst : DFF_X1 port map( D => n11829, CK => CLK, Q => n54259, 
                           QN => n2201);
   REGS_reg_78_15_inst : DFF_X1 port map( D => n11828, CK => CLK, Q => n54260, 
                           QN => n2202);
   REGS_reg_78_14_inst : DFF_X1 port map( D => n11827, CK => CLK, Q => n54261, 
                           QN => n2203);
   REGS_reg_78_13_inst : DFF_X1 port map( D => n11826, CK => CLK, Q => n54262, 
                           QN => n2204);
   REGS_reg_78_12_inst : DFF_X1 port map( D => n11825, CK => CLK, Q => n54263, 
                           QN => n2205);
   REGS_reg_78_11_inst : DFF_X1 port map( D => n11824, CK => CLK, Q => n54264, 
                           QN => n2206);
   REGS_reg_78_10_inst : DFF_X1 port map( D => n11823, CK => CLK, Q => n54265, 
                           QN => n2207);
   REGS_reg_78_9_inst : DFF_X1 port map( D => n11822, CK => CLK, Q => n54266, 
                           QN => n2208);
   REGS_reg_78_8_inst : DFF_X1 port map( D => n11821, CK => CLK, Q => n54267, 
                           QN => n2209);
   REGS_reg_78_7_inst : DFF_X1 port map( D => n11820, CK => CLK, Q => n54268, 
                           QN => n2210);
   REGS_reg_78_6_inst : DFF_X1 port map( D => n11819, CK => CLK, Q => n54269, 
                           QN => n2211);
   REGS_reg_78_5_inst : DFF_X1 port map( D => n11818, CK => CLK, Q => n54270, 
                           QN => n2212);
   REGS_reg_78_4_inst : DFF_X1 port map( D => n11817, CK => CLK, Q => n54271, 
                           QN => n2221);
   REGS_reg_78_3_inst : DFF_X1 port map( D => n11816, CK => CLK, Q => n54272, 
                           QN => n2222);
   REGS_reg_78_2_inst : DFF_X1 port map( D => n11815, CK => CLK, Q => n54273, 
                           QN => n2223);
   REGS_reg_78_1_inst : DFF_X1 port map( D => n11814, CK => CLK, Q => n54274, 
                           QN => n2224);
   REGS_reg_78_0_inst : DFF_X1 port map( D => n11813, CK => CLK, Q => n54275, 
                           QN => n2225);
   REGS_reg_77_23_inst : DFF_X1 port map( D => n11868, CK => CLK, Q => n_1936, 
                           QN => n2226);
   REGS_reg_77_22_inst : DFF_X1 port map( D => n11867, CK => CLK, Q => n_1937, 
                           QN => n2227);
   REGS_reg_77_21_inst : DFF_X1 port map( D => n11866, CK => CLK, Q => n_1938, 
                           QN => n2228);
   REGS_reg_77_20_inst : DFF_X1 port map( D => n11865, CK => CLK, Q => n_1939, 
                           QN => n2229);
   REGS_reg_77_19_inst : DFF_X1 port map( D => n11864, CK => CLK, Q => n_1940, 
                           QN => n2230);
   REGS_reg_77_18_inst : DFF_X1 port map( D => n11863, CK => CLK, Q => n_1941, 
                           QN => n2231);
   REGS_reg_77_17_inst : DFF_X1 port map( D => n11862, CK => CLK, Q => n_1942, 
                           QN => n2232);
   REGS_reg_77_16_inst : DFF_X1 port map( D => n11861, CK => CLK, Q => n_1943, 
                           QN => n2233);
   REGS_reg_77_15_inst : DFF_X1 port map( D => n11860, CK => CLK, Q => n_1944, 
                           QN => n2234);
   REGS_reg_77_14_inst : DFF_X1 port map( D => n11859, CK => CLK, Q => n_1945, 
                           QN => n2271);
   REGS_reg_77_13_inst : DFF_X1 port map( D => n11858, CK => CLK, Q => n_1946, 
                           QN => n2272);
   REGS_reg_77_12_inst : DFF_X1 port map( D => n11857, CK => CLK, Q => n_1947, 
                           QN => n2273);
   REGS_reg_77_11_inst : DFF_X1 port map( D => n11856, CK => CLK, Q => n_1948, 
                           QN => n2274);
   REGS_reg_77_10_inst : DFF_X1 port map( D => n11855, CK => CLK, Q => n_1949, 
                           QN => n2275);
   REGS_reg_77_9_inst : DFF_X1 port map( D => n11854, CK => CLK, Q => n_1950, 
                           QN => n2276);
   REGS_reg_77_8_inst : DFF_X1 port map( D => n11853, CK => CLK, Q => n_1951, 
                           QN => n2277);
   REGS_reg_77_7_inst : DFF_X1 port map( D => n11852, CK => CLK, Q => n_1952, 
                           QN => n2278);
   REGS_reg_77_6_inst : DFF_X1 port map( D => n11851, CK => CLK, Q => n_1953, 
                           QN => n2279);
   REGS_reg_77_5_inst : DFF_X1 port map( D => n11850, CK => CLK, Q => n_1954, 
                           QN => n2280);
   REGS_reg_77_4_inst : DFF_X1 port map( D => n11849, CK => CLK, Q => n_1955, 
                           QN => n2281);
   REGS_reg_77_3_inst : DFF_X1 port map( D => n11848, CK => CLK, Q => n_1956, 
                           QN => n2282);
   REGS_reg_77_2_inst : DFF_X1 port map( D => n11847, CK => CLK, Q => n_1957, 
                           QN => n2283);
   REGS_reg_77_1_inst : DFF_X1 port map( D => n11846, CK => CLK, Q => n_1958, 
                           QN => n2284);
   REGS_reg_77_0_inst : DFF_X1 port map( D => n11845, CK => CLK, Q => n_1959, 
                           QN => n2285);
   REGS_reg_76_23_inst : DFF_X1 port map( D => n11900, CK => CLK, Q => n_1960, 
                           QN => n2286);
   REGS_reg_76_22_inst : DFF_X1 port map( D => n11899, CK => CLK, Q => n_1961, 
                           QN => n2287);
   REGS_reg_76_21_inst : DFF_X1 port map( D => n11898, CK => CLK, Q => n_1962, 
                           QN => n2288);
   REGS_reg_76_20_inst : DFF_X1 port map( D => n11897, CK => CLK, Q => n_1963, 
                           QN => n2289);
   REGS_reg_76_19_inst : DFF_X1 port map( D => n11896, CK => CLK, Q => n_1964, 
                           QN => n2290);
   REGS_reg_76_18_inst : DFF_X1 port map( D => n11895, CK => CLK, Q => n_1965, 
                           QN => n2291);
   REGS_reg_76_17_inst : DFF_X1 port map( D => n11894, CK => CLK, Q => n_1966, 
                           QN => n2292);
   REGS_reg_76_16_inst : DFF_X1 port map( D => n11893, CK => CLK, Q => n_1967, 
                           QN => n2293);
   REGS_reg_76_15_inst : DFF_X1 port map( D => n11892, CK => CLK, Q => n_1968, 
                           QN => n2294);
   REGS_reg_76_14_inst : DFF_X1 port map( D => n11891, CK => CLK, Q => n_1969, 
                           QN => n2295);
   REGS_reg_76_13_inst : DFF_X1 port map( D => n11890, CK => CLK, Q => n_1970, 
                           QN => n2296);
   REGS_reg_76_12_inst : DFF_X1 port map( D => n11889, CK => CLK, Q => n_1971, 
                           QN => n2297);
   REGS_reg_76_11_inst : DFF_X1 port map( D => n11888, CK => CLK, Q => n_1972, 
                           QN => n2298);
   REGS_reg_76_10_inst : DFF_X1 port map( D => n11887, CK => CLK, Q => n_1973, 
                           QN => n2391);
   REGS_reg_76_9_inst : DFF_X1 port map( D => n11886, CK => CLK, Q => n_1974, 
                           QN => n2392);
   REGS_reg_76_8_inst : DFF_X1 port map( D => n11885, CK => CLK, Q => n_1975, 
                           QN => n2393);
   REGS_reg_76_7_inst : DFF_X1 port map( D => n11884, CK => CLK, Q => n_1976, 
                           QN => n2394);
   REGS_reg_76_6_inst : DFF_X1 port map( D => n11883, CK => CLK, Q => n_1977, 
                           QN => n2395);
   REGS_reg_76_5_inst : DFF_X1 port map( D => n11882, CK => CLK, Q => n_1978, 
                           QN => n2396);
   REGS_reg_76_4_inst : DFF_X1 port map( D => n11881, CK => CLK, Q => n_1979, 
                           QN => n2397);
   REGS_reg_76_3_inst : DFF_X1 port map( D => n11880, CK => CLK, Q => n_1980, 
                           QN => n2398);
   REGS_reg_76_2_inst : DFF_X1 port map( D => n11879, CK => CLK, Q => n_1981, 
                           QN => n2399);
   REGS_reg_76_1_inst : DFF_X1 port map( D => n11878, CK => CLK, Q => n_1982, 
                           QN => n2400);
   REGS_reg_76_0_inst : DFF_X1 port map( D => n11877, CK => CLK, Q => n_1983, 
                           QN => n2401);
   REGS_reg_75_23_inst : DFF_X1 port map( D => n11932, CK => CLK, Q => n54638, 
                           QN => n2402);
   REGS_reg_75_22_inst : DFF_X1 port map( D => n11931, CK => CLK, Q => n54637, 
                           QN => n2403);
   REGS_reg_75_21_inst : DFF_X1 port map( D => n11930, CK => CLK, Q => n54636, 
                           QN => n2404);
   REGS_reg_75_20_inst : DFF_X1 port map( D => n11929, CK => CLK, Q => n54635, 
                           QN => n2405);
   REGS_reg_75_19_inst : DFF_X1 port map( D => n11928, CK => CLK, Q => n54634, 
                           QN => n2406);
   REGS_reg_75_18_inst : DFF_X1 port map( D => n11927, CK => CLK, Q => n54633, 
                           QN => n2407);
   REGS_reg_75_17_inst : DFF_X1 port map( D => n11926, CK => CLK, Q => n54632, 
                           QN => n2408);
   REGS_reg_75_16_inst : DFF_X1 port map( D => n11925, CK => CLK, Q => n54631, 
                           QN => n2409);
   REGS_reg_75_15_inst : DFF_X1 port map( D => n11924, CK => CLK, Q => n54630, 
                           QN => n2410);
   REGS_reg_75_14_inst : DFF_X1 port map( D => n11923, CK => CLK, Q => n54629, 
                           QN => n2411);
   REGS_reg_75_13_inst : DFF_X1 port map( D => n11922, CK => CLK, Q => n54628, 
                           QN => n2412);
   REGS_reg_75_12_inst : DFF_X1 port map( D => n11921, CK => CLK, Q => n54627, 
                           QN => n2413);
   REGS_reg_75_11_inst : DFF_X1 port map( D => n11920, CK => CLK, Q => n54626, 
                           QN => n2414);
   REGS_reg_75_10_inst : DFF_X1 port map( D => n11919, CK => CLK, Q => n54625, 
                           QN => n2415);
   REGS_reg_75_9_inst : DFF_X1 port map( D => n11918, CK => CLK, Q => n54624, 
                           QN => n2416);
   REGS_reg_75_8_inst : DFF_X1 port map( D => n11917, CK => CLK, Q => n54623, 
                           QN => n2417);
   REGS_reg_75_7_inst : DFF_X1 port map( D => n11916, CK => CLK, Q => n54646, 
                           QN => n2418);
   REGS_reg_75_6_inst : DFF_X1 port map( D => n11915, CK => CLK, Q => n54645, 
                           QN => n2419);
   REGS_reg_75_5_inst : DFF_X1 port map( D => n11914, CK => CLK, Q => n54644, 
                           QN => n2420);
   REGS_reg_75_4_inst : DFF_X1 port map( D => n11913, CK => CLK, Q => n54643, 
                           QN => n2421);
   REGS_reg_75_3_inst : DFF_X1 port map( D => n11912, CK => CLK, Q => n54642, 
                           QN => n2422);
   REGS_reg_75_2_inst : DFF_X1 port map( D => n11911, CK => CLK, Q => n54641, 
                           QN => n2423);
   REGS_reg_75_1_inst : DFF_X1 port map( D => n11910, CK => CLK, Q => n54640, 
                           QN => n2424);
   REGS_reg_75_0_inst : DFF_X1 port map( D => n11909, CK => CLK, Q => n54639, 
                           QN => n2425);
   REGS_reg_74_23_inst : DFF_X1 port map( D => n11964, CK => CLK, Q => n54494, 
                           QN => n2426);
   REGS_reg_74_22_inst : DFF_X1 port map( D => n11963, CK => CLK, Q => n54493, 
                           QN => n2427);
   REGS_reg_74_21_inst : DFF_X1 port map( D => n11962, CK => CLK, Q => n54492, 
                           QN => n2428);
   REGS_reg_74_20_inst : DFF_X1 port map( D => n11961, CK => CLK, Q => n54491, 
                           QN => n2429);
   REGS_reg_74_19_inst : DFF_X1 port map( D => n11960, CK => CLK, Q => n54490, 
                           QN => n2430);
   REGS_reg_74_18_inst : DFF_X1 port map( D => n11959, CK => CLK, Q => n54489, 
                           QN => n2431);
   REGS_reg_74_17_inst : DFF_X1 port map( D => n11958, CK => CLK, Q => n54488, 
                           QN => n2432);
   REGS_reg_74_16_inst : DFF_X1 port map( D => n11957, CK => CLK, Q => n54487, 
                           QN => n2433);
   REGS_reg_74_15_inst : DFF_X1 port map( D => n11956, CK => CLK, Q => n54486, 
                           QN => n2434);
   REGS_reg_74_14_inst : DFF_X1 port map( D => n11955, CK => CLK, Q => n54485, 
                           QN => n2435);
   REGS_reg_74_13_inst : DFF_X1 port map( D => n11954, CK => CLK, Q => n54484, 
                           QN => n2436);
   REGS_reg_74_12_inst : DFF_X1 port map( D => n11953, CK => CLK, Q => n54483, 
                           QN => n2437);
   REGS_reg_74_11_inst : DFF_X1 port map( D => n11952, CK => CLK, Q => n54482, 
                           QN => n2438);
   REGS_reg_74_10_inst : DFF_X1 port map( D => n11951, CK => CLK, Q => n54481, 
                           QN => n2463);
   REGS_reg_74_9_inst : DFF_X1 port map( D => n11950, CK => CLK, Q => n54480, 
                           QN => n2464);
   REGS_reg_74_8_inst : DFF_X1 port map( D => n11949, CK => CLK, Q => n54479, 
                           QN => n2465);
   REGS_reg_74_7_inst : DFF_X1 port map( D => n11948, CK => CLK, Q => n54502, 
                           QN => n2466);
   REGS_reg_74_6_inst : DFF_X1 port map( D => n11947, CK => CLK, Q => n54501, 
                           QN => n2467);
   REGS_reg_74_5_inst : DFF_X1 port map( D => n11946, CK => CLK, Q => n54500, 
                           QN => n2468);
   REGS_reg_74_4_inst : DFF_X1 port map( D => n11945, CK => CLK, Q => n54499, 
                           QN => n2469);
   REGS_reg_74_3_inst : DFF_X1 port map( D => n11944, CK => CLK, Q => n54498, 
                           QN => n2470);
   REGS_reg_74_2_inst : DFF_X1 port map( D => n11943, CK => CLK, Q => n54497, 
                           QN => n2471);
   REGS_reg_74_1_inst : DFF_X1 port map( D => n11942, CK => CLK, Q => n54496, 
                           QN => n2472);
   REGS_reg_74_0_inst : DFF_X1 port map( D => n11941, CK => CLK, Q => n54495, 
                           QN => n2473);
   REGS_reg_73_23_inst : DFF_X1 port map( D => n11996, CK => CLK, Q => n_1984, 
                           QN => n2474);
   REGS_reg_73_22_inst : DFF_X1 port map( D => n11995, CK => CLK, Q => n_1985, 
                           QN => n2475);
   REGS_reg_73_21_inst : DFF_X1 port map( D => n11994, CK => CLK, Q => n_1986, 
                           QN => n2476);
   REGS_reg_73_20_inst : DFF_X1 port map( D => n11993, CK => CLK, Q => n_1987, 
                           QN => n2477);
   REGS_reg_73_19_inst : DFF_X1 port map( D => n11992, CK => CLK, Q => n_1988, 
                           QN => n2478);
   REGS_reg_73_18_inst : DFF_X1 port map( D => n11991, CK => CLK, Q => n_1989, 
                           QN => n2479);
   REGS_reg_73_17_inst : DFF_X1 port map( D => n11990, CK => CLK, Q => n_1990, 
                           QN => n2480);
   REGS_reg_73_16_inst : DFF_X1 port map( D => n11989, CK => CLK, Q => n_1991, 
                           QN => n2481);
   REGS_reg_73_15_inst : DFF_X1 port map( D => n11988, CK => CLK, Q => n_1992, 
                           QN => n2482);
   REGS_reg_73_14_inst : DFF_X1 port map( D => n11987, CK => CLK, Q => n_1993, 
                           QN => n2511);
   REGS_reg_73_13_inst : DFF_X1 port map( D => n11986, CK => CLK, Q => n_1994, 
                           QN => n2512);
   REGS_reg_73_12_inst : DFF_X1 port map( D => n11985, CK => CLK, Q => n_1995, 
                           QN => n2513);
   REGS_reg_73_11_inst : DFF_X1 port map( D => n11984, CK => CLK, Q => n_1996, 
                           QN => n2514);
   REGS_reg_73_10_inst : DFF_X1 port map( D => n11983, CK => CLK, Q => n_1997, 
                           QN => n2515);
   REGS_reg_73_9_inst : DFF_X1 port map( D => n11982, CK => CLK, Q => n_1998, 
                           QN => n2516);
   REGS_reg_73_8_inst : DFF_X1 port map( D => n11981, CK => CLK, Q => n_1999, 
                           QN => n2517);
   REGS_reg_73_7_inst : DFF_X1 port map( D => n11980, CK => CLK, Q => n_2000, 
                           QN => n2518);
   REGS_reg_73_6_inst : DFF_X1 port map( D => n11979, CK => CLK, Q => n_2001, 
                           QN => n2519);
   REGS_reg_73_5_inst : DFF_X1 port map( D => n11978, CK => CLK, Q => n_2002, 
                           QN => n2520);
   REGS_reg_73_4_inst : DFF_X1 port map( D => n11977, CK => CLK, Q => n_2003, 
                           QN => n2521);
   REGS_reg_73_3_inst : DFF_X1 port map( D => n11976, CK => CLK, Q => n_2004, 
                           QN => n2522);
   REGS_reg_73_2_inst : DFF_X1 port map( D => n11975, CK => CLK, Q => n_2005, 
                           QN => n2523);
   REGS_reg_73_1_inst : DFF_X1 port map( D => n11974, CK => CLK, Q => n_2006, 
                           QN => n2524);
   REGS_reg_73_0_inst : DFF_X1 port map( D => n11973, CK => CLK, Q => n_2007, 
                           QN => n2525);
   REGS_reg_72_23_inst : DFF_X1 port map( D => n12028, CK => CLK, Q => n_2008, 
                           QN => n2526);
   REGS_reg_72_22_inst : DFF_X1 port map( D => n12027, CK => CLK, Q => n_2009, 
                           QN => n2527);
   REGS_reg_72_21_inst : DFF_X1 port map( D => n12026, CK => CLK, Q => n_2010, 
                           QN => n2528);
   REGS_reg_72_20_inst : DFF_X1 port map( D => n12025, CK => CLK, Q => n_2011, 
                           QN => n2529);
   REGS_reg_72_19_inst : DFF_X1 port map( D => n12024, CK => CLK, Q => n_2012, 
                           QN => n2530);
   REGS_reg_72_18_inst : DFF_X1 port map( D => n12023, CK => CLK, Q => n_2013, 
                           QN => n2531);
   REGS_reg_72_17_inst : DFF_X1 port map( D => n12022, CK => CLK, Q => n_2014, 
                           QN => n2532);
   REGS_reg_72_16_inst : DFF_X1 port map( D => n12021, CK => CLK, Q => n_2015, 
                           QN => n2533);
   REGS_reg_72_15_inst : DFF_X1 port map( D => n12020, CK => CLK, Q => n_2016, 
                           QN => n2534);
   REGS_reg_72_14_inst : DFF_X1 port map( D => n12019, CK => CLK, Q => n_2017, 
                           QN => n2535);
   REGS_reg_72_13_inst : DFF_X1 port map( D => n12018, CK => CLK, Q => n_2018, 
                           QN => n2536);
   REGS_reg_72_12_inst : DFF_X1 port map( D => n12017, CK => CLK, Q => n_2019, 
                           QN => n2537);
   REGS_reg_72_11_inst : DFF_X1 port map( D => n12016, CK => CLK, Q => n_2020, 
                           QN => n2538);
   REGS_reg_72_10_inst : DFF_X1 port map( D => n12015, CK => CLK, Q => n_2021, 
                           QN => n2539);
   REGS_reg_72_9_inst : DFF_X1 port map( D => n12014, CK => CLK, Q => n_2022, 
                           QN => n2540);
   REGS_reg_72_8_inst : DFF_X1 port map( D => n12013, CK => CLK, Q => n_2023, 
                           QN => n2541);
   REGS_reg_72_7_inst : DFF_X1 port map( D => n12012, CK => CLK, Q => n_2024, 
                           QN => n2542);
   REGS_reg_72_6_inst : DFF_X1 port map( D => n12011, CK => CLK, Q => n_2025, 
                           QN => n2543);
   REGS_reg_72_5_inst : DFF_X1 port map( D => n12010, CK => CLK, Q => n_2026, 
                           QN => n2544);
   REGS_reg_72_4_inst : DFF_X1 port map( D => n12009, CK => CLK, Q => n_2027, 
                           QN => n2545);
   REGS_reg_72_3_inst : DFF_X1 port map( D => n12008, CK => CLK, Q => n_2028, 
                           QN => n2546);
   REGS_reg_72_2_inst : DFF_X1 port map( D => n12007, CK => CLK, Q => n_2029, 
                           QN => n2547);
   REGS_reg_72_1_inst : DFF_X1 port map( D => n12006, CK => CLK, Q => n_2030, 
                           QN => n2548);
   REGS_reg_72_0_inst : DFF_X1 port map( D => n12005, CK => CLK, Q => n_2031, 
                           QN => n2549);
   REGS_reg_71_23_inst : DFF_X1 port map( D => n12060, CK => CLK, Q => n54324, 
                           QN => n2550);
   REGS_reg_71_22_inst : DFF_X1 port map( D => n12059, CK => CLK, Q => n54325, 
                           QN => n2551);
   REGS_reg_71_21_inst : DFF_X1 port map( D => n12058, CK => CLK, Q => n54326, 
                           QN => n2552);
   REGS_reg_71_20_inst : DFF_X1 port map( D => n12057, CK => CLK, Q => n54327, 
                           QN => n2553);
   REGS_reg_71_19_inst : DFF_X1 port map( D => n12056, CK => CLK, Q => n54328, 
                           QN => n2554);
   REGS_reg_71_18_inst : DFF_X1 port map( D => n12055, CK => CLK, Q => n54329, 
                           QN => n2555);
   REGS_reg_71_17_inst : DFF_X1 port map( D => n12054, CK => CLK, Q => n54330, 
                           QN => n2556);
   REGS_reg_71_16_inst : DFF_X1 port map( D => n12053, CK => CLK, Q => n54331, 
                           QN => n2557);
   REGS_reg_71_15_inst : DFF_X1 port map( D => n12052, CK => CLK, Q => n54332, 
                           QN => n2558);
   REGS_reg_71_14_inst : DFF_X1 port map( D => n12051, CK => CLK, Q => n54333, 
                           QN => n2559);
   REGS_reg_71_13_inst : DFF_X1 port map( D => n12050, CK => CLK, Q => n54334, 
                           QN => n2560);
   REGS_reg_71_12_inst : DFF_X1 port map( D => n12049, CK => CLK, Q => n54335, 
                           QN => n2561);
   REGS_reg_71_11_inst : DFF_X1 port map( D => n12048, CK => CLK, Q => n54336, 
                           QN => n2562);
   REGS_reg_71_10_inst : DFF_X1 port map( D => n12047, CK => CLK, Q => n54337, 
                           QN => n2563);
   REGS_reg_71_9_inst : DFF_X1 port map( D => n12046, CK => CLK, Q => n54338, 
                           QN => n2564);
   REGS_reg_71_8_inst : DFF_X1 port map( D => n12045, CK => CLK, Q => n54339, 
                           QN => n2565);
   REGS_reg_71_7_inst : DFF_X1 port map( D => n12044, CK => CLK, Q => n54340, 
                           QN => n2566);
   REGS_reg_71_6_inst : DFF_X1 port map( D => n12043, CK => CLK, Q => n54341, 
                           QN => n2567);
   REGS_reg_71_5_inst : DFF_X1 port map( D => n12042, CK => CLK, Q => n54342, 
                           QN => n2568);
   REGS_reg_71_4_inst : DFF_X1 port map( D => n12041, CK => CLK, Q => n54343, 
                           QN => n2569);
   REGS_reg_71_3_inst : DFF_X1 port map( D => n12040, CK => CLK, Q => n54344, 
                           QN => n2570);
   REGS_reg_71_2_inst : DFF_X1 port map( D => n12039, CK => CLK, Q => n54345, 
                           QN => n2571);
   REGS_reg_71_1_inst : DFF_X1 port map( D => n12038, CK => CLK, Q => n54346, 
                           QN => n2572);
   REGS_reg_71_0_inst : DFF_X1 port map( D => n12037, CK => CLK, Q => n54347, 
                           QN => n2573);
   REGS_reg_70_23_inst : DFF_X1 port map( D => n12092, CK => CLK, Q => n54348, 
                           QN => n2574);
   REGS_reg_70_22_inst : DFF_X1 port map( D => n12091, CK => CLK, Q => n54349, 
                           QN => n2575);
   REGS_reg_70_21_inst : DFF_X1 port map( D => n12090, CK => CLK, Q => n54350, 
                           QN => n2576);
   REGS_reg_70_20_inst : DFF_X1 port map( D => n12089, CK => CLK, Q => n54351, 
                           QN => n2577);
   REGS_reg_70_19_inst : DFF_X1 port map( D => n12088, CK => CLK, Q => n54352, 
                           QN => n2578);
   REGS_reg_70_18_inst : DFF_X1 port map( D => n12087, CK => CLK, Q => n54353, 
                           QN => n2579);
   REGS_reg_70_17_inst : DFF_X1 port map( D => n12086, CK => CLK, Q => n54354, 
                           QN => n2580);
   REGS_reg_70_16_inst : DFF_X1 port map( D => n12085, CK => CLK, Q => n54355, 
                           QN => n2581);
   REGS_reg_70_15_inst : DFF_X1 port map( D => n12084, CK => CLK, Q => n54356, 
                           QN => n2582);
   REGS_reg_70_14_inst : DFF_X1 port map( D => n12083, CK => CLK, Q => n54357, 
                           QN => n2583);
   REGS_reg_70_13_inst : DFF_X1 port map( D => n12082, CK => CLK, Q => n54358, 
                           QN => n2584);
   REGS_reg_70_12_inst : DFF_X1 port map( D => n12081, CK => CLK, Q => n54359, 
                           QN => n2585);
   REGS_reg_70_11_inst : DFF_X1 port map( D => n12080, CK => CLK, Q => n54360, 
                           QN => n2586);
   REGS_reg_70_10_inst : DFF_X1 port map( D => n12079, CK => CLK, Q => n54361, 
                           QN => n2587);
   REGS_reg_70_9_inst : DFF_X1 port map( D => n12078, CK => CLK, Q => n54362, 
                           QN => n2588);
   REGS_reg_70_8_inst : DFF_X1 port map( D => n12077, CK => CLK, Q => n54363, 
                           QN => n2589);
   REGS_reg_70_7_inst : DFF_X1 port map( D => n12076, CK => CLK, Q => n54364, 
                           QN => n2590);
   REGS_reg_70_6_inst : DFF_X1 port map( D => n12075, CK => CLK, Q => n54365, 
                           QN => n2591);
   REGS_reg_70_5_inst : DFF_X1 port map( D => n12074, CK => CLK, Q => n54366, 
                           QN => n2592);
   REGS_reg_70_4_inst : DFF_X1 port map( D => n12073, CK => CLK, Q => n54367, 
                           QN => n2593);
   REGS_reg_70_3_inst : DFF_X1 port map( D => n12072, CK => CLK, Q => n54368, 
                           QN => n2594);
   REGS_reg_70_2_inst : DFF_X1 port map( D => n12071, CK => CLK, Q => n54369, 
                           QN => n2595);
   REGS_reg_70_1_inst : DFF_X1 port map( D => n12070, CK => CLK, Q => n54370, 
                           QN => n2596);
   REGS_reg_70_0_inst : DFF_X1 port map( D => n12069, CK => CLK, Q => n54371, 
                           QN => n2597);
   REGS_reg_69_23_inst : DFF_X1 port map( D => n12124, CK => CLK, Q => n_2032, 
                           QN => n2598);
   REGS_reg_69_22_inst : DFF_X1 port map( D => n12123, CK => CLK, Q => n_2033, 
                           QN => n2599);
   REGS_reg_69_21_inst : DFF_X1 port map( D => n12122, CK => CLK, Q => n_2034, 
                           QN => n2600);
   REGS_reg_69_20_inst : DFF_X1 port map( D => n12121, CK => CLK, Q => n_2035, 
                           QN => n2601);
   REGS_reg_69_19_inst : DFF_X1 port map( D => n12120, CK => CLK, Q => n_2036, 
                           QN => n2602);
   REGS_reg_69_18_inst : DFF_X1 port map( D => n12119, CK => CLK, Q => n_2037, 
                           QN => n2603);
   REGS_reg_69_17_inst : DFF_X1 port map( D => n12118, CK => CLK, Q => n_2038, 
                           QN => n2604);
   REGS_reg_69_16_inst : DFF_X1 port map( D => n12117, CK => CLK, Q => n_2039, 
                           QN => n2605);
   REGS_reg_69_15_inst : DFF_X1 port map( D => n12116, CK => CLK, Q => n_2040, 
                           QN => n2606);
   REGS_reg_69_14_inst : DFF_X1 port map( D => n12115, CK => CLK, Q => n_2041, 
                           QN => n2607);
   REGS_reg_69_13_inst : DFF_X1 port map( D => n12114, CK => CLK, Q => n_2042, 
                           QN => n2608);
   REGS_reg_69_12_inst : DFF_X1 port map( D => n12113, CK => CLK, Q => n_2043, 
                           QN => n2609);
   REGS_reg_69_11_inst : DFF_X1 port map( D => n12112, CK => CLK, Q => n_2044, 
                           QN => n2610);
   REGS_reg_69_10_inst : DFF_X1 port map( D => n12111, CK => CLK, Q => n_2045, 
                           QN => n2611);
   REGS_reg_69_9_inst : DFF_X1 port map( D => n12110, CK => CLK, Q => n_2046, 
                           QN => n2612);
   REGS_reg_69_8_inst : DFF_X1 port map( D => n12109, CK => CLK, Q => n_2047, 
                           QN => n2613);
   REGS_reg_69_7_inst : DFF_X1 port map( D => n12108, CK => CLK, Q => n_2048, 
                           QN => n2614);
   REGS_reg_69_6_inst : DFF_X1 port map( D => n12107, CK => CLK, Q => n_2049, 
                           QN => n2615);
   REGS_reg_69_5_inst : DFF_X1 port map( D => n12106, CK => CLK, Q => n_2050, 
                           QN => n2616);
   REGS_reg_69_4_inst : DFF_X1 port map( D => n12105, CK => CLK, Q => n_2051, 
                           QN => n2617);
   REGS_reg_69_3_inst : DFF_X1 port map( D => n12104, CK => CLK, Q => n_2052, 
                           QN => n2618);
   REGS_reg_69_2_inst : DFF_X1 port map( D => n12103, CK => CLK, Q => n_2053, 
                           QN => n2619);
   REGS_reg_69_1_inst : DFF_X1 port map( D => n12102, CK => CLK, Q => n_2054, 
                           QN => n2620);
   REGS_reg_69_0_inst : DFF_X1 port map( D => n12101, CK => CLK, Q => n_2055, 
                           QN => n2621);
   REGS_reg_68_23_inst : DFF_X1 port map( D => n12156, CK => CLK, Q => n_2056, 
                           QN => n2622);
   REGS_reg_68_22_inst : DFF_X1 port map( D => n12155, CK => CLK, Q => n_2057, 
                           QN => n2623);
   REGS_reg_68_21_inst : DFF_X1 port map( D => n12154, CK => CLK, Q => n_2058, 
                           QN => n2624);
   REGS_reg_68_20_inst : DFF_X1 port map( D => n12153, CK => CLK, Q => n_2059, 
                           QN => n2625);
   REGS_reg_68_19_inst : DFF_X1 port map( D => n12152, CK => CLK, Q => n_2060, 
                           QN => n2626);
   REGS_reg_68_18_inst : DFF_X1 port map( D => n12151, CK => CLK, Q => n_2061, 
                           QN => n2627);
   REGS_reg_68_17_inst : DFF_X1 port map( D => n12150, CK => CLK, Q => n_2062, 
                           QN => n2628);
   REGS_reg_68_16_inst : DFF_X1 port map( D => n12149, CK => CLK, Q => n_2063, 
                           QN => n2629);
   REGS_reg_68_15_inst : DFF_X1 port map( D => n12148, CK => CLK, Q => n_2064, 
                           QN => n2630);
   REGS_reg_68_14_inst : DFF_X1 port map( D => n12147, CK => CLK, Q => n_2065, 
                           QN => n2631);
   REGS_reg_68_13_inst : DFF_X1 port map( D => n12146, CK => CLK, Q => n_2066, 
                           QN => n2632);
   REGS_reg_68_12_inst : DFF_X1 port map( D => n12145, CK => CLK, Q => n_2067, 
                           QN => n2633);
   REGS_reg_68_11_inst : DFF_X1 port map( D => n12144, CK => CLK, Q => n_2068, 
                           QN => n2634);
   REGS_reg_68_10_inst : DFF_X1 port map( D => n12143, CK => CLK, Q => n_2069, 
                           QN => n2635);
   REGS_reg_68_9_inst : DFF_X1 port map( D => n12142, CK => CLK, Q => n_2070, 
                           QN => n2636);
   REGS_reg_68_8_inst : DFF_X1 port map( D => n12141, CK => CLK, Q => n_2071, 
                           QN => n2637);
   REGS_reg_68_7_inst : DFF_X1 port map( D => n12140, CK => CLK, Q => n_2072, 
                           QN => n2638);
   REGS_reg_68_6_inst : DFF_X1 port map( D => n12139, CK => CLK, Q => n_2073, 
                           QN => n2639);
   REGS_reg_68_5_inst : DFF_X1 port map( D => n12138, CK => CLK, Q => n_2074, 
                           QN => n2640);
   REGS_reg_68_4_inst : DFF_X1 port map( D => n12137, CK => CLK, Q => n_2075, 
                           QN => n2641);
   REGS_reg_68_3_inst : DFF_X1 port map( D => n12136, CK => CLK, Q => n_2076, 
                           QN => n2642);
   REGS_reg_68_2_inst : DFF_X1 port map( D => n12135, CK => CLK, Q => n_2077, 
                           QN => n2643);
   REGS_reg_68_1_inst : DFF_X1 port map( D => n12134, CK => CLK, Q => n_2078, 
                           QN => n2644);
   REGS_reg_68_0_inst : DFF_X1 port map( D => n12133, CK => CLK, Q => n_2079, 
                           QN => n2652);
   REGS_reg_67_23_inst : DFF_X1 port map( D => n12188, CK => CLK, Q => n54372, 
                           QN => n2653);
   REGS_reg_67_22_inst : DFF_X1 port map( D => n12187, CK => CLK, Q => n54373, 
                           QN => n2654);
   REGS_reg_67_21_inst : DFF_X1 port map( D => n12186, CK => CLK, Q => n54374, 
                           QN => n2655);
   REGS_reg_67_20_inst : DFF_X1 port map( D => n12185, CK => CLK, Q => n54375, 
                           QN => n2656);
   REGS_reg_67_19_inst : DFF_X1 port map( D => n12184, CK => CLK, Q => n54376, 
                           QN => n2657);
   REGS_reg_67_18_inst : DFF_X1 port map( D => n12183, CK => CLK, Q => n54377, 
                           QN => n2658);
   REGS_reg_67_17_inst : DFF_X1 port map( D => n12182, CK => CLK, Q => n54378, 
                           QN => n2659);
   REGS_reg_67_16_inst : DFF_X1 port map( D => n12181, CK => CLK, Q => n54379, 
                           QN => n2660);
   REGS_reg_67_15_inst : DFF_X1 port map( D => n12180, CK => CLK, Q => n54380, 
                           QN => n2661);
   REGS_reg_67_14_inst : DFF_X1 port map( D => n12179, CK => CLK, Q => n54381, 
                           QN => n2662);
   REGS_reg_67_13_inst : DFF_X1 port map( D => n12178, CK => CLK, Q => n54382, 
                           QN => n2663);
   REGS_reg_67_12_inst : DFF_X1 port map( D => n12177, CK => CLK, Q => n54383, 
                           QN => n2664);
   REGS_reg_67_11_inst : DFF_X1 port map( D => n12176, CK => CLK, Q => n54384, 
                           QN => n2665);
   REGS_reg_67_10_inst : DFF_X1 port map( D => n12175, CK => CLK, Q => n54385, 
                           QN => n2666);
   REGS_reg_67_9_inst : DFF_X1 port map( D => n12174, CK => CLK, Q => n54386, 
                           QN => n2667);
   REGS_reg_67_8_inst : DFF_X1 port map( D => n12173, CK => CLK, Q => n54387, 
                           QN => n2668);
   REGS_reg_67_7_inst : DFF_X1 port map( D => n12172, CK => CLK, Q => n54388, 
                           QN => n2669);
   REGS_reg_67_6_inst : DFF_X1 port map( D => n12171, CK => CLK, Q => n54389, 
                           QN => n2670);
   REGS_reg_67_5_inst : DFF_X1 port map( D => n12170, CK => CLK, Q => n54390, 
                           QN => n2671);
   REGS_reg_67_4_inst : DFF_X1 port map( D => n12169, CK => CLK, Q => n54391, 
                           QN => n2672);
   REGS_reg_67_3_inst : DFF_X1 port map( D => n12168, CK => CLK, Q => n54392, 
                           QN => n2673);
   REGS_reg_67_2_inst : DFF_X1 port map( D => n12167, CK => CLK, Q => n54393, 
                           QN => n2674);
   REGS_reg_67_1_inst : DFF_X1 port map( D => n12166, CK => CLK, Q => n54394, 
                           QN => n2675);
   REGS_reg_67_0_inst : DFF_X1 port map( D => n12165, CK => CLK, Q => n54395, 
                           QN => n2676);
   REGS_reg_66_23_inst : DFF_X1 port map( D => n12220, CK => CLK, Q => n54553, 
                           QN => n2677);
   REGS_reg_66_22_inst : DFF_X1 port map( D => n12219, CK => CLK, Q => n54552, 
                           QN => n2678);
   REGS_reg_66_21_inst : DFF_X1 port map( D => n12218, CK => CLK, Q => n54551, 
                           QN => n2679);
   REGS_reg_66_20_inst : DFF_X1 port map( D => n12217, CK => CLK, Q => n54550, 
                           QN => n2680);
   REGS_reg_66_19_inst : DFF_X1 port map( D => n12216, CK => CLK, Q => n54549, 
                           QN => n2681);
   REGS_reg_66_18_inst : DFF_X1 port map( D => n12215, CK => CLK, Q => n54548, 
                           QN => n2682);
   REGS_reg_66_17_inst : DFF_X1 port map( D => n12214, CK => CLK, Q => n54547, 
                           QN => n2683);
   REGS_reg_66_16_inst : DFF_X1 port map( D => n12213, CK => CLK, Q => n54546, 
                           QN => n2684);
   REGS_reg_66_15_inst : DFF_X1 port map( D => n12212, CK => CLK, Q => n54545, 
                           QN => n2685);
   REGS_reg_66_14_inst : DFF_X1 port map( D => n12211, CK => CLK, Q => n54544, 
                           QN => n2686);
   REGS_reg_66_13_inst : DFF_X1 port map( D => n12210, CK => CLK, Q => n54543, 
                           QN => n2687);
   REGS_reg_66_12_inst : DFF_X1 port map( D => n12209, CK => CLK, Q => n54558, 
                           QN => n2688);
   REGS_reg_65_23_inst : DFF_X1 port map( D => n12252, CK => CLK, Q => n54396, 
                           QN => n2701);
   REGS_reg_65_22_inst : DFF_X1 port map( D => n12251, CK => CLK, Q => n54397, 
                           QN => n2702);
   REGS_reg_65_21_inst : DFF_X1 port map( D => n12250, CK => CLK, Q => n54398, 
                           QN => n2703);
   REGS_reg_65_20_inst : DFF_X1 port map( D => n12249, CK => CLK, Q => n54399, 
                           QN => n2704);
   REGS_reg_65_19_inst : DFF_X1 port map( D => n12248, CK => CLK, Q => n54400, 
                           QN => n2705);
   REGS_reg_65_18_inst : DFF_X1 port map( D => n12247, CK => CLK, Q => n54401, 
                           QN => n2706);
   REGS_reg_65_17_inst : DFF_X1 port map( D => n12246, CK => CLK, Q => n54402, 
                           QN => n2707);
   REGS_reg_65_16_inst : DFF_X1 port map( D => n12245, CK => CLK, Q => n54403, 
                           QN => n2708);
   REGS_reg_65_15_inst : DFF_X1 port map( D => n12244, CK => CLK, Q => n54404, 
                           QN => n2709);
   REGS_reg_65_14_inst : DFF_X1 port map( D => n12243, CK => CLK, Q => n54405, 
                           QN => n2710);
   REGS_reg_65_13_inst : DFF_X1 port map( D => n12242, CK => CLK, Q => n54406, 
                           QN => n2711);
   REGS_reg_65_12_inst : DFF_X1 port map( D => n12241, CK => CLK, Q => n54407, 
                           QN => n2712);
   REGS_reg_65_11_inst : DFF_X1 port map( D => n12240, CK => CLK, Q => n54408, 
                           QN => n2713);
   REGS_reg_65_10_inst : DFF_X1 port map( D => n12239, CK => CLK, Q => n54409, 
                           QN => n2714);
   REGS_reg_65_9_inst : DFF_X1 port map( D => n12238, CK => CLK, Q => n54410, 
                           QN => n2715);
   REGS_reg_65_8_inst : DFF_X1 port map( D => n12237, CK => CLK, Q => n54411, 
                           QN => n2716);
   REGS_reg_65_7_inst : DFF_X1 port map( D => n12236, CK => CLK, Q => n54412, 
                           QN => n2717);
   REGS_reg_65_6_inst : DFF_X1 port map( D => n12235, CK => CLK, Q => n54413, 
                           QN => n2718);
   REGS_reg_65_5_inst : DFF_X1 port map( D => n12234, CK => CLK, Q => n54414, 
                           QN => n2719);
   REGS_reg_65_4_inst : DFF_X1 port map( D => n12233, CK => CLK, Q => n54415, 
                           QN => n2720);
   REGS_reg_65_3_inst : DFF_X1 port map( D => n12232, CK => CLK, Q => n54416, 
                           QN => n2721);
   REGS_reg_65_2_inst : DFF_X1 port map( D => n12231, CK => CLK, Q => n54417, 
                           QN => n2722);
   REGS_reg_65_1_inst : DFF_X1 port map( D => n12230, CK => CLK, Q => n54418, 
                           QN => n2723);
   REGS_reg_65_0_inst : DFF_X1 port map( D => n12229, CK => CLK, Q => n54419, 
                           QN => n2724);
   REGS_reg_134_2_inst : DFF_X1 port map( D => n10023, CK => CLK, Q => n54564, 
                           QN => n3927);
   REGS_reg_134_1_inst : DFF_X1 port map( D => n10022, CK => CLK, Q => n54563, 
                           QN => n3928);
   REGS_reg_134_0_inst : DFF_X1 port map( D => n10021, CK => CLK, Q => n54575, 
                           QN => n3929);
   REGS_reg_134_23_inst : DFF_X1 port map( D => n10044, CK => CLK, Q => n54574,
                           QN => n3930);
   REGS_reg_134_22_inst : DFF_X1 port map( D => n10043, CK => CLK, Q => n54573,
                           QN => n3931);
   REGS_reg_134_21_inst : DFF_X1 port map( D => n10042, CK => CLK, Q => n54572,
                           QN => n3932);
   REGS_reg_134_20_inst : DFF_X1 port map( D => n10041, CK => CLK, Q => n54571,
                           QN => n3933);
   REGS_reg_134_19_inst : DFF_X1 port map( D => n10040, CK => CLK, Q => n54570,
                           QN => n3934);
   REGS_reg_133_28_inst : DFF_X1 port map( D => n10081, CK => CLK, Q => n3935, 
                           QN => n52239);
   REGS_reg_133_27_inst : DFF_X1 port map( D => n10080, CK => CLK, Q => n3936, 
                           QN => n52240);
   REGS_reg_133_26_inst : DFF_X1 port map( D => n10079, CK => CLK, Q => n3937, 
                           QN => n52241);
   REGS_reg_133_25_inst : DFF_X1 port map( D => n10078, CK => CLK, Q => n3938, 
                           QN => n52242);
   REGS_reg_133_24_inst : DFF_X1 port map( D => n10077, CK => CLK, Q => n3939, 
                           QN => n52243);
   REGS_reg_63_31_inst : DFF_X1 port map( D => n12324, CK => CLK, Q => n_2080, 
                           QN => n474);
   REGS_reg_63_30_inst : DFF_X1 port map( D => n12323, CK => CLK, Q => n_2081, 
                           QN => n475);
   REGS_reg_63_29_inst : DFF_X1 port map( D => n12322, CK => CLK, Q => n_2082, 
                           QN => n500);
   REGS_reg_63_28_inst : DFF_X1 port map( D => n12321, CK => CLK, Q => n_2083, 
                           QN => n501);
   REGS_reg_63_27_inst : DFF_X1 port map( D => n12320, CK => CLK, Q => n_2084, 
                           QN => n502);
   REGS_reg_63_26_inst : DFF_X1 port map( D => n12319, CK => CLK, Q => n_2085, 
                           QN => n503);
   REGS_reg_63_25_inst : DFF_X1 port map( D => n12318, CK => CLK, Q => n_2086, 
                           QN => n504);
   REGS_reg_63_24_inst : DFF_X1 port map( D => n12317, CK => CLK, Q => n_2087, 
                           QN => n505);
   REGS_reg_54_31_inst : DFF_X1 port map( D => n12612, CK => CLK, Q => n771, QN
                           => n539);
   REGS_reg_54_30_inst : DFF_X1 port map( D => n12611, CK => CLK, Q => n772, QN
                           => n540);
   REGS_reg_54_29_inst : DFF_X1 port map( D => n12610, CK => CLK, Q => n773, QN
                           => n541);
   REGS_reg_54_28_inst : DFF_X1 port map( D => n12609, CK => CLK, Q => n774, QN
                           => n542);
   REGS_reg_54_27_inst : DFF_X1 port map( D => n12608, CK => CLK, Q => n775, QN
                           => n543);
   REGS_reg_54_26_inst : DFF_X1 port map( D => n12607, CK => CLK, Q => n784, QN
                           => n544);
   REGS_reg_54_25_inst : DFF_X1 port map( D => n12606, CK => CLK, Q => n785, QN
                           => n545);
   REGS_reg_54_24_inst : DFF_X1 port map( D => n12605, CK => CLK, Q => n786, QN
                           => n546);
   REGS_reg_39_31_inst : DFF_X1 port map( D => n13092, CK => CLK, Q => n4257, 
                           QN => n9779);
   REGS_reg_39_30_inst : DFF_X1 port map( D => n13091, CK => CLK, Q => n4258, 
                           QN => n9780);
   REGS_reg_39_29_inst : DFF_X1 port map( D => n13090, CK => CLK, Q => n4259, 
                           QN => n9781);
   REGS_reg_39_28_inst : DFF_X1 port map( D => n13089, CK => CLK, Q => n4260, 
                           QN => n9782);
   REGS_reg_39_27_inst : DFF_X1 port map( D => n13088, CK => CLK, Q => n4261, 
                           QN => n9783);
   REGS_reg_39_26_inst : DFF_X1 port map( D => n13087, CK => CLK, Q => n4262, 
                           QN => n9784);
   REGS_reg_39_25_inst : DFF_X1 port map( D => n13086, CK => CLK, Q => n4263, 
                           QN => n9785);
   REGS_reg_39_24_inst : DFF_X1 port map( D => n13085, CK => CLK, Q => n4264, 
                           QN => n9786);
   REGS_reg_38_31_inst : DFF_X1 port map( D => n13124, CK => CLK, Q => n4265, 
                           QN => n9747);
   REGS_reg_38_30_inst : DFF_X1 port map( D => n13123, CK => CLK, Q => n4266, 
                           QN => n9748);
   REGS_reg_38_29_inst : DFF_X1 port map( D => n13122, CK => CLK, Q => n4267, 
                           QN => n9749);
   REGS_reg_38_28_inst : DFF_X1 port map( D => n13121, CK => CLK, Q => n4268, 
                           QN => n9750);
   REGS_reg_38_27_inst : DFF_X1 port map( D => n13120, CK => CLK, Q => n4269, 
                           QN => n9751);
   REGS_reg_38_26_inst : DFF_X1 port map( D => n13119, CK => CLK, Q => n4270, 
                           QN => n9752);
   REGS_reg_38_25_inst : DFF_X1 port map( D => n13118, CK => CLK, Q => n4271, 
                           QN => n9753);
   REGS_reg_38_24_inst : DFF_X1 port map( D => n13117, CK => CLK, Q => n4272, 
                           QN => n9754);
   REGS_reg_28_31_inst : DFF_X1 port map( D => n13444, CK => CLK, Q => n3956, 
                           QN => n9611);
   REGS_reg_28_30_inst : DFF_X1 port map( D => n13443, CK => CLK, Q => n3957, 
                           QN => n9612);
   REGS_reg_28_29_inst : DFF_X1 port map( D => n13442, CK => CLK, Q => n3958, 
                           QN => n9613);
   REGS_reg_28_28_inst : DFF_X1 port map( D => n13441, CK => CLK, Q => n3959, 
                           QN => n9614);
   REGS_reg_28_27_inst : DFF_X1 port map( D => n13440, CK => CLK, Q => n3960, 
                           QN => n9615);
   REGS_reg_28_26_inst : DFF_X1 port map( D => n13439, CK => CLK, Q => n3961, 
                           QN => n9616);
   REGS_reg_28_25_inst : DFF_X1 port map( D => n13438, CK => CLK, Q => n3962, 
                           QN => n9617);
   REGS_reg_28_24_inst : DFF_X1 port map( D => n13437, CK => CLK, Q => n3963, 
                           QN => n9618);
   REGS_reg_27_31_inst : DFF_X1 port map( D => n13476, CK => CLK, Q => n3964, 
                           QN => n9603);
   REGS_reg_27_30_inst : DFF_X1 port map( D => n13475, CK => CLK, Q => n3965, 
                           QN => n9604);
   REGS_reg_27_29_inst : DFF_X1 port map( D => n13474, CK => CLK, Q => n3966, 
                           QN => n9605);
   REGS_reg_27_28_inst : DFF_X1 port map( D => n13473, CK => CLK, Q => n3991, 
                           QN => n9606);
   REGS_reg_27_27_inst : DFF_X1 port map( D => n13472, CK => CLK, Q => n3992, 
                           QN => n9607);
   REGS_reg_27_26_inst : DFF_X1 port map( D => n13471, CK => CLK, Q => n3993, 
                           QN => n9608);
   REGS_reg_27_25_inst : DFF_X1 port map( D => n13470, CK => CLK, Q => n3994, 
                           QN => n9609);
   REGS_reg_27_24_inst : DFF_X1 port map( D => n13469, CK => CLK, Q => n3995, 
                           QN => n9610);
   REGS_reg_22_31_inst : DFF_X1 port map( D => n13636, CK => CLK, Q => n104, QN
                           => n816);
   REGS_reg_22_30_inst : DFF_X1 port map( D => n13635, CK => CLK, Q => n105, QN
                           => n817);
   REGS_reg_22_29_inst : DFF_X1 port map( D => n13634, CK => CLK, Q => n106, QN
                           => n818);
   REGS_reg_22_28_inst : DFF_X1 port map( D => n13633, CK => CLK, Q => n107, QN
                           => n819);
   REGS_reg_22_27_inst : DFF_X1 port map( D => n13632, CK => CLK, Q => n108, QN
                           => n820);
   REGS_reg_22_26_inst : DFF_X1 port map( D => n13631, CK => CLK, Q => n109, QN
                           => n821);
   REGS_reg_22_25_inst : DFF_X1 port map( D => n13630, CK => CLK, Q => n110, QN
                           => n822);
   REGS_reg_22_24_inst : DFF_X1 port map( D => n13629, CK => CLK, Q => n111, QN
                           => n823);
   REGS_reg_21_31_inst : DFF_X1 port map( D => n13668, CK => CLK, Q => n_2088, 
                           QN => n824);
   REGS_reg_21_30_inst : DFF_X1 port map( D => n13667, CK => CLK, Q => n_2089, 
                           QN => n825);
   REGS_reg_21_29_inst : DFF_X1 port map( D => n13666, CK => CLK, Q => n_2090, 
                           QN => n826);
   REGS_reg_21_28_inst : DFF_X1 port map( D => n13665, CK => CLK, Q => n_2091, 
                           QN => n827);
   REGS_reg_21_27_inst : DFF_X1 port map( D => n13664, CK => CLK, Q => n_2092, 
                           QN => n828);
   REGS_reg_21_26_inst : DFF_X1 port map( D => n13663, CK => CLK, Q => n_2093, 
                           QN => n829);
   REGS_reg_21_25_inst : DFF_X1 port map( D => n13662, CK => CLK, Q => n_2094, 
                           QN => n830);
   REGS_reg_21_24_inst : DFF_X1 port map( D => n13661, CK => CLK, Q => n_2095, 
                           QN => n831);
   REGS_reg_20_31_inst : DFF_X1 port map( D => n13700, CK => CLK, Q => n112, QN
                           => n2909);
   REGS_reg_20_30_inst : DFF_X1 port map( D => n13699, CK => CLK, Q => n113, QN
                           => n2910);
   REGS_reg_20_29_inst : DFF_X1 port map( D => n13698, CK => CLK, Q => n114, QN
                           => n2911);
   REGS_reg_20_28_inst : DFF_X1 port map( D => n13697, CK => CLK, Q => n115, QN
                           => n2912);
   REGS_reg_20_27_inst : DFF_X1 port map( D => n13696, CK => CLK, Q => n116, QN
                           => n2913);
   REGS_reg_20_26_inst : DFF_X1 port map( D => n13695, CK => CLK, Q => n117, QN
                           => n2914);
   REGS_reg_20_25_inst : DFF_X1 port map( D => n13694, CK => CLK, Q => n118, QN
                           => n2915);
   REGS_reg_20_24_inst : DFF_X1 port map( D => n13693, CK => CLK, Q => n119, QN
                           => n2916);
   REGS_reg_19_31_inst : DFF_X1 port map( D => n13732, CK => CLK, Q => n120, QN
                           => n2917);
   REGS_reg_19_30_inst : DFF_X1 port map( D => n13731, CK => CLK, Q => n121, QN
                           => n2918);
   REGS_reg_19_29_inst : DFF_X1 port map( D => n13730, CK => CLK, Q => n122, QN
                           => n2919);
   REGS_reg_19_28_inst : DFF_X1 port map( D => n13729, CK => CLK, Q => n123, QN
                           => n2920);
   REGS_reg_19_27_inst : DFF_X1 port map( D => n13728, CK => CLK, Q => n124, QN
                           => n2921);
   REGS_reg_19_26_inst : DFF_X1 port map( D => n13727, CK => CLK, Q => n125, QN
                           => n2922);
   REGS_reg_19_25_inst : DFF_X1 port map( D => n13726, CK => CLK, Q => n126, QN
                           => n2923);
   REGS_reg_19_24_inst : DFF_X1 port map( D => n13725, CK => CLK, Q => n127, QN
                           => n2924);
   REGS_reg_3_31_inst : DFF_X1 port map( D => n14244, CK => CLK, Q => n4164, QN
                           => n51632);
   REGS_reg_3_30_inst : DFF_X1 port map( D => n14243, CK => CLK, Q => n4165, QN
                           => n51633);
   REGS_reg_3_29_inst : DFF_X1 port map( D => n14242, CK => CLK, Q => n4166, QN
                           => n51634);
   REGS_reg_3_28_inst : DFF_X1 port map( D => n14241, CK => CLK, Q => n4167, QN
                           => n51635);
   REGS_reg_3_27_inst : DFF_X1 port map( D => n14240, CK => CLK, Q => n4168, QN
                           => n51636);
   REGS_reg_3_26_inst : DFF_X1 port map( D => n14239, CK => CLK, Q => n4169, QN
                           => n51637);
   REGS_reg_3_25_inst : DFF_X1 port map( D => n14238, CK => CLK, Q => n4170, QN
                           => n51638);
   REGS_reg_3_24_inst : DFF_X1 port map( D => n14237, CK => CLK, Q => n4171, QN
                           => n51639);
   REGS_reg_2_31_inst : DFF_X1 port map( D => n14276, CK => CLK, Q => n4172, QN
                           => n51640);
   REGS_reg_2_30_inst : DFF_X1 port map( D => n14275, CK => CLK, Q => n4173, QN
                           => n51641);
   REGS_reg_2_29_inst : DFF_X1 port map( D => n14274, CK => CLK, Q => n4174, QN
                           => n51642);
   REGS_reg_2_28_inst : DFF_X1 port map( D => n14273, CK => CLK, Q => n4175, QN
                           => n51643);
   REGS_reg_2_27_inst : DFF_X1 port map( D => n14272, CK => CLK, Q => n4176, QN
                           => n51644);
   REGS_reg_2_26_inst : DFF_X1 port map( D => n14271, CK => CLK, Q => n4177, QN
                           => n51645);
   REGS_reg_2_25_inst : DFF_X1 port map( D => n14270, CK => CLK, Q => n4178, QN
                           => n51646);
   REGS_reg_2_24_inst : DFF_X1 port map( D => n14269, CK => CLK, Q => n4179, QN
                           => n51647);
   REGS_reg_126_31_inst : DFF_X1 port map( D => n10308, CK => CLK, Q => n4289, 
                           QN => n15331);
   REGS_reg_126_30_inst : DFF_X1 port map( D => n10307, CK => CLK, Q => n4290, 
                           QN => n15332);
   REGS_reg_126_29_inst : DFF_X1 port map( D => n10306, CK => CLK, Q => n4291, 
                           QN => n15333);
   REGS_reg_126_28_inst : DFF_X1 port map( D => n10305, CK => CLK, Q => n4292, 
                           QN => n15334);
   REGS_reg_126_27_inst : DFF_X1 port map( D => n10304, CK => CLK, Q => n4293, 
                           QN => n15335);
   REGS_reg_126_26_inst : DFF_X1 port map( D => n10303, CK => CLK, Q => n4294, 
                           QN => n15336);
   REGS_reg_126_25_inst : DFF_X1 port map( D => n10302, CK => CLK, Q => n4295, 
                           QN => n15337);
   REGS_reg_126_24_inst : DFF_X1 port map( D => n10301, CK => CLK, Q => n4296, 
                           QN => n15338);
   REGS_reg_125_31_inst : DFF_X1 port map( D => n10340, CK => CLK, Q => n4297, 
                           QN => n15299);
   REGS_reg_125_30_inst : DFF_X1 port map( D => n10339, CK => CLK, Q => n4298, 
                           QN => n15300);
   REGS_reg_125_29_inst : DFF_X1 port map( D => n10338, CK => CLK, Q => n4299, 
                           QN => n15301);
   REGS_reg_125_28_inst : DFF_X1 port map( D => n10337, CK => CLK, Q => n4300, 
                           QN => n15302);
   REGS_reg_125_27_inst : DFF_X1 port map( D => n10336, CK => CLK, Q => n4301, 
                           QN => n15303);
   REGS_reg_125_26_inst : DFF_X1 port map( D => n10335, CK => CLK, Q => n4302, 
                           QN => n15304);
   REGS_reg_125_25_inst : DFF_X1 port map( D => n10334, CK => CLK, Q => n4303, 
                           QN => n15305);
   REGS_reg_125_24_inst : DFF_X1 port map( D => n10333, CK => CLK, Q => n4304, 
                           QN => n15306);
   REGS_reg_122_31_inst : DFF_X1 port map( D => n10436, CK => CLK, Q => n4305, 
                           QN => n52496);
   REGS_reg_122_30_inst : DFF_X1 port map( D => n10435, CK => CLK, Q => n4306, 
                           QN => n52497);
   REGS_reg_122_29_inst : DFF_X1 port map( D => n10434, CK => CLK, Q => n4307, 
                           QN => n52498);
   REGS_reg_122_28_inst : DFF_X1 port map( D => n10433, CK => CLK, Q => n4308, 
                           QN => n52499);
   REGS_reg_122_27_inst : DFF_X1 port map( D => n10432, CK => CLK, Q => n4309, 
                           QN => n52500);
   REGS_reg_122_26_inst : DFF_X1 port map( D => n10431, CK => CLK, Q => n4310, 
                           QN => n52501);
   REGS_reg_122_25_inst : DFF_X1 port map( D => n10430, CK => CLK, Q => n4311, 
                           QN => n52502);
   REGS_reg_122_24_inst : DFF_X1 port map( D => n10429, CK => CLK, Q => n4312, 
                           QN => n52503);
   REGS_reg_121_31_inst : DFF_X1 port map( D => n10468, CK => CLK, Q => n4313, 
                           QN => n52504);
   REGS_reg_121_30_inst : DFF_X1 port map( D => n10467, CK => CLK, Q => n4314, 
                           QN => n52505);
   REGS_reg_121_29_inst : DFF_X1 port map( D => n10466, CK => CLK, Q => n4315, 
                           QN => n52506);
   REGS_reg_121_28_inst : DFF_X1 port map( D => n10465, CK => CLK, Q => n4316, 
                           QN => n52507);
   REGS_reg_115_31_inst : DFF_X1 port map( D => n10660, CK => CLK, Q => n4317, 
                           QN => n15203);
   REGS_reg_115_30_inst : DFF_X1 port map( D => n10659, CK => CLK, Q => n4318, 
                           QN => n15204);
   REGS_reg_115_29_inst : DFF_X1 port map( D => n10658, CK => CLK, Q => n4319, 
                           QN => n15205);
   REGS_reg_115_28_inst : DFF_X1 port map( D => n10657, CK => CLK, Q => n4320, 
                           QN => n15206);
   REGS_reg_115_27_inst : DFF_X1 port map( D => n10656, CK => CLK, Q => n4321, 
                           QN => n15207);
   REGS_reg_115_26_inst : DFF_X1 port map( D => n10655, CK => CLK, Q => n4322, 
                           QN => n15208);
   REGS_reg_115_25_inst : DFF_X1 port map( D => n10654, CK => CLK, Q => n4323, 
                           QN => n15209);
   REGS_reg_115_24_inst : DFF_X1 port map( D => n10653, CK => CLK, Q => n4324, 
                           QN => n15210);
   REGS_reg_114_31_inst : DFF_X1 port map( D => n10692, CK => CLK, Q => n4325, 
                           QN => n15171);
   REGS_reg_114_30_inst : DFF_X1 port map( D => n10691, CK => CLK, Q => n4326, 
                           QN => n15172);
   REGS_reg_114_29_inst : DFF_X1 port map( D => n10690, CK => CLK, Q => n4327, 
                           QN => n15173);
   REGS_reg_114_28_inst : DFF_X1 port map( D => n10689, CK => CLK, Q => n4328, 
                           QN => n15174);
   REGS_reg_114_27_inst : DFF_X1 port map( D => n10688, CK => CLK, Q => n4329, 
                           QN => n15175);
   REGS_reg_114_26_inst : DFF_X1 port map( D => n10687, CK => CLK, Q => n4330, 
                           QN => n15176);
   REGS_reg_114_25_inst : DFF_X1 port map( D => n10686, CK => CLK, Q => n4331, 
                           QN => n15177);
   REGS_reg_83_31_inst : DFF_X1 port map( D => n11684, CK => CLK, Q => n4028, 
                           QN => n52664);
   REGS_reg_83_30_inst : DFF_X1 port map( D => n11683, CK => CLK, Q => n4029, 
                           QN => n52665);
   REGS_reg_83_29_inst : DFF_X1 port map( D => n11682, CK => CLK, Q => n4030, 
                           QN => n52666);
   REGS_reg_83_28_inst : DFF_X1 port map( D => n11681, CK => CLK, Q => n4031, 
                           QN => n52667);
   REGS_reg_83_27_inst : DFF_X1 port map( D => n11680, CK => CLK, Q => n4032, 
                           QN => n52668);
   REGS_reg_83_26_inst : DFF_X1 port map( D => n11679, CK => CLK, Q => n4033, 
                           QN => n52669);
   REGS_reg_83_25_inst : DFF_X1 port map( D => n11678, CK => CLK, Q => n4034, 
                           QN => n52670);
   REGS_reg_83_24_inst : DFF_X1 port map( D => n11677, CK => CLK, Q => n4035, 
                           QN => n52671);
   REGS_reg_82_31_inst : DFF_X1 port map( D => n11716, CK => CLK, Q => n4036, 
                           QN => n52672);
   REGS_reg_82_30_inst : DFF_X1 port map( D => n11715, CK => CLK, Q => n4037, 
                           QN => n52673);
   REGS_reg_82_29_inst : DFF_X1 port map( D => n11714, CK => CLK, Q => n4038, 
                           QN => n52674);
   REGS_reg_82_28_inst : DFF_X1 port map( D => n11713, CK => CLK, Q => n4039, 
                           QN => n52675);
   REGS_reg_82_27_inst : DFF_X1 port map( D => n11712, CK => CLK, Q => n4040, 
                           QN => n52676);
   REGS_reg_82_26_inst : DFF_X1 port map( D => n11711, CK => CLK, Q => n4041, 
                           QN => n52677);
   REGS_reg_82_25_inst : DFF_X1 port map( D => n11710, CK => CLK, Q => n4042, 
                           QN => n52678);
   REGS_reg_82_24_inst : DFF_X1 port map( D => n11709, CK => CLK, Q => n4043, 
                           QN => n52679);
   REGS_reg_67_31_inst : DFF_X1 port map( D => n12196, CK => CLK, Q => n4076, 
                           QN => n52728);
   REGS_reg_67_30_inst : DFF_X1 port map( D => n12195, CK => CLK, Q => n4077, 
                           QN => n52729);
   REGS_reg_67_29_inst : DFF_X1 port map( D => n12194, CK => CLK, Q => n4078, 
                           QN => n52730);
   REGS_reg_67_28_inst : DFF_X1 port map( D => n12193, CK => CLK, Q => n4079, 
                           QN => n52731);
   REGS_reg_67_27_inst : DFF_X1 port map( D => n12192, CK => CLK, Q => n4080, 
                           QN => n52732);
   REGS_reg_67_26_inst : DFF_X1 port map( D => n12191, CK => CLK, Q => n4081, 
                           QN => n52733);
   REGS_reg_67_25_inst : DFF_X1 port map( D => n12190, CK => CLK, Q => n4082, 
                           QN => n52734);
   REGS_reg_67_24_inst : DFF_X1 port map( D => n12189, CK => CLK, Q => n4083, 
                           QN => n52735);
   REGS_reg_66_31_inst : DFF_X1 port map( D => n12228, CK => CLK, Q => n4084, 
                           QN => n52736);
   REGS_reg_66_30_inst : DFF_X1 port map( D => n12227, CK => CLK, Q => n4085, 
                           QN => n52737);
   REGS_reg_66_29_inst : DFF_X1 port map( D => n12226, CK => CLK, Q => n4086, 
                           QN => n52738);
   REGS_reg_66_28_inst : DFF_X1 port map( D => n12225, CK => CLK, Q => n4087, 
                           QN => n52739);
   REGS_reg_66_27_inst : DFF_X1 port map( D => n12224, CK => CLK, Q => n4088, 
                           QN => n52740);
   REGS_reg_66_26_inst : DFF_X1 port map( D => n12223, CK => CLK, Q => n4089, 
                           QN => n52741);
   REGS_reg_66_25_inst : DFF_X1 port map( D => n12222, CK => CLK, Q => n4090, 
                           QN => n52742);
   REGS_reg_66_24_inst : DFF_X1 port map( D => n12221, CK => CLK, Q => n4091, 
                           QN => n52743);
   REGS_reg_65_31_inst : DFF_X1 port map( D => n12260, CK => CLK, Q => n4092, 
                           QN => n52744);
   REGS_reg_65_30_inst : DFF_X1 port map( D => n12259, CK => CLK, Q => n4093, 
                           QN => n52745);
   REGS_reg_65_29_inst : DFF_X1 port map( D => n12258, CK => CLK, Q => n4094, 
                           QN => n52746);
   REGS_reg_65_28_inst : DFF_X1 port map( D => n12257, CK => CLK, Q => n4095, 
                           QN => n52747);
   REGS_reg_65_27_inst : DFF_X1 port map( D => n12256, CK => CLK, Q => n4096, 
                           QN => n52748);
   REGS_reg_65_26_inst : DFF_X1 port map( D => n12255, CK => CLK, Q => n4097, 
                           QN => n52749);
   REGS_reg_65_25_inst : DFF_X1 port map( D => n12254, CK => CLK, Q => n4098, 
                           QN => n52750);
   REGS_reg_65_24_inst : DFF_X1 port map( D => n12253, CK => CLK, Q => n4099, 
                           QN => n52751);
   REGS_reg_28_23_inst : DFF_X1 port map( D => n13436, CK => CLK, Q => n4332, 
                           QN => n52928);
   REGS_reg_28_22_inst : DFF_X1 port map( D => n13435, CK => CLK, Q => n4333, 
                           QN => n52929);
   REGS_reg_28_21_inst : DFF_X1 port map( D => n13434, CK => CLK, Q => n4334, 
                           QN => n52930);
   REGS_reg_28_20_inst : DFF_X1 port map( D => n13433, CK => CLK, Q => n4335, 
                           QN => n52931);
   REGS_reg_28_19_inst : DFF_X1 port map( D => n13432, CK => CLK, Q => n4336, 
                           QN => n52932);
   REGS_reg_28_18_inst : DFF_X1 port map( D => n13431, CK => CLK, Q => n4337, 
                           QN => n52933);
   REGS_reg_28_17_inst : DFF_X1 port map( D => n13430, CK => CLK, Q => n4338, 
                           QN => n52934);
   REGS_reg_28_16_inst : DFF_X1 port map( D => n13429, CK => CLK, Q => n4339, 
                           QN => n52935);
   REGS_reg_28_15_inst : DFF_X1 port map( D => n13428, CK => CLK, Q => n4340, 
                           QN => n52936);
   REGS_reg_28_14_inst : DFF_X1 port map( D => n13427, CK => CLK, Q => n4341, 
                           QN => n52937);
   REGS_reg_28_13_inst : DFF_X1 port map( D => n13426, CK => CLK, Q => n4342, 
                           QN => n52938);
   REGS_reg_28_12_inst : DFF_X1 port map( D => n13425, CK => CLK, Q => n4343, 
                           QN => n52939);
   REGS_reg_28_11_inst : DFF_X1 port map( D => n13424, CK => CLK, Q => n4344, 
                           QN => n52940);
   REGS_reg_28_10_inst : DFF_X1 port map( D => n13423, CK => CLK, Q => n4345, 
                           QN => n52941);
   REGS_reg_28_9_inst : DFF_X1 port map( D => n13422, CK => CLK, Q => n4346, QN
                           => n52942);
   REGS_reg_28_8_inst : DFF_X1 port map( D => n13421, CK => CLK, Q => n4347, QN
                           => n52943);
   REGS_reg_28_7_inst : DFF_X1 port map( D => n13420, CK => CLK, Q => n4348, QN
                           => n52944);
   REGS_reg_28_6_inst : DFF_X1 port map( D => n13419, CK => CLK, Q => n4349, QN
                           => n52945);
   REGS_reg_28_5_inst : DFF_X1 port map( D => n13418, CK => CLK, Q => n4350, QN
                           => n52946);
   REGS_reg_28_4_inst : DFF_X1 port map( D => n13417, CK => CLK, Q => n4351, QN
                           => n52947);
   REGS_reg_28_3_inst : DFF_X1 port map( D => n13416, CK => CLK, Q => n4352, QN
                           => n52948);
   REGS_reg_28_2_inst : DFF_X1 port map( D => n13415, CK => CLK, Q => n4353, QN
                           => n52949);
   REGS_reg_28_1_inst : DFF_X1 port map( D => n13414, CK => CLK, Q => n4354, QN
                           => n52950);
   REGS_reg_28_0_inst : DFF_X1 port map( D => n13413, CK => CLK, Q => n4355, QN
                           => n52951);
   REGS_reg_27_23_inst : DFF_X1 port map( D => n13468, CK => CLK, Q => n4356, 
                           QN => n51808);
   REGS_reg_27_22_inst : DFF_X1 port map( D => n13467, CK => CLK, Q => n4357, 
                           QN => n51809);
   REGS_reg_27_21_inst : DFF_X1 port map( D => n13466, CK => CLK, Q => n4358, 
                           QN => n51810);
   REGS_reg_27_20_inst : DFF_X1 port map( D => n13465, CK => CLK, Q => n4359, 
                           QN => n51811);
   REGS_reg_27_19_inst : DFF_X1 port map( D => n13464, CK => CLK, Q => n4360, 
                           QN => n51812);
   REGS_reg_27_18_inst : DFF_X1 port map( D => n13463, CK => CLK, Q => n4361, 
                           QN => n51813);
   REGS_reg_27_17_inst : DFF_X1 port map( D => n13462, CK => CLK, Q => n4362, 
                           QN => n51814);
   REGS_reg_27_16_inst : DFF_X1 port map( D => n13461, CK => CLK, Q => n4363, 
                           QN => n51815);
   REGS_reg_27_15_inst : DFF_X1 port map( D => n13460, CK => CLK, Q => n4364, 
                           QN => n51816);
   REGS_reg_27_14_inst : DFF_X1 port map( D => n13459, CK => CLK, Q => n4365, 
                           QN => n51817);
   REGS_reg_27_13_inst : DFF_X1 port map( D => n13458, CK => CLK, Q => n4366, 
                           QN => n51818);
   REGS_reg_27_12_inst : DFF_X1 port map( D => n13457, CK => CLK, Q => n4367, 
                           QN => n51819);
   REGS_reg_27_11_inst : DFF_X1 port map( D => n13456, CK => CLK, Q => n4368, 
                           QN => n51820);
   REGS_reg_27_10_inst : DFF_X1 port map( D => n13455, CK => CLK, Q => n4369, 
                           QN => n51821);
   REGS_reg_27_9_inst : DFF_X1 port map( D => n13454, CK => CLK, Q => n4370, QN
                           => n51822);
   REGS_reg_27_8_inst : DFF_X1 port map( D => n13453, CK => CLK, Q => n4371, QN
                           => n51823);
   REGS_reg_27_7_inst : DFF_X1 port map( D => n13452, CK => CLK, Q => n4372, QN
                           => n51824);
   REGS_reg_27_6_inst : DFF_X1 port map( D => n13451, CK => CLK, Q => n4373, QN
                           => n51825);
   REGS_reg_27_5_inst : DFF_X1 port map( D => n13450, CK => CLK, Q => n4374, QN
                           => n51826);
   REGS_reg_27_3_inst : DFF_X1 port map( D => n13448, CK => CLK, Q => n4375, QN
                           => n52952);
   REGS_reg_27_2_inst : DFF_X1 port map( D => n13447, CK => CLK, Q => n4376, QN
                           => n52953);
   REGS_reg_27_1_inst : DFF_X1 port map( D => n13446, CK => CLK, Q => n4377, QN
                           => n52954);
   REGS_reg_27_0_inst : DFF_X1 port map( D => n13445, CK => CLK, Q => n4378, QN
                           => n52955);
   REGS_reg_21_13_inst : DFF_X1 port map( D => n13650, CK => CLK, Q => n_2096, 
                           QN => n1575);
   REGS_reg_21_12_inst : DFF_X1 port map( D => n13649, CK => CLK, Q => n_2097, 
                           QN => n1576);
   REGS_reg_21_11_inst : DFF_X1 port map( D => n13648, CK => CLK, Q => n_2098, 
                           QN => n1577);
   REGS_reg_21_10_inst : DFF_X1 port map( D => n13647, CK => CLK, Q => n_2099, 
                           QN => n1578);
   REGS_reg_21_9_inst : DFF_X1 port map( D => n13646, CK => CLK, Q => n_2100, 
                           QN => n1579);
   REGS_reg_21_8_inst : DFF_X1 port map( D => n13645, CK => CLK, Q => n_2101, 
                           QN => n1580);
   REGS_reg_21_7_inst : DFF_X1 port map( D => n13644, CK => CLK, Q => n_2102, 
                           QN => n1581);
   REGS_reg_21_6_inst : DFF_X1 port map( D => n13643, CK => CLK, Q => n_2103, 
                           QN => n1582);
   REGS_reg_21_5_inst : DFF_X1 port map( D => n13642, CK => CLK, Q => n_2104, 
                           QN => n1583);
   REGS_reg_21_4_inst : DFF_X1 port map( D => n13641, CK => CLK, Q => n_2105, 
                           QN => n1584);
   REGS_reg_21_3_inst : DFF_X1 port map( D => n13640, CK => CLK, Q => n_2106, 
                           QN => n1585);
   REGS_reg_21_2_inst : DFF_X1 port map( D => n13639, CK => CLK, Q => n_2107, 
                           QN => n1586);
   REGS_reg_21_1_inst : DFF_X1 port map( D => n13638, CK => CLK, Q => n_2108, 
                           QN => n1587);
   REGS_reg_21_0_inst : DFF_X1 port map( D => n13637, CK => CLK, Q => n_2109, 
                           QN => n1588);
   REGS_reg_20_23_inst : DFF_X1 port map( D => n13692, CK => CLK, Q => n1739, 
                           QN => n3409);
   REGS_reg_20_22_inst : DFF_X1 port map( D => n13691, CK => CLK, Q => n1740, 
                           QN => n3410);
   REGS_reg_20_21_inst : DFF_X1 port map( D => n13690, CK => CLK, Q => n1741, 
                           QN => n3411);
   REGS_reg_20_20_inst : DFF_X1 port map( D => n13689, CK => CLK, Q => n1742, 
                           QN => n3412);
   REGS_reg_20_19_inst : DFF_X1 port map( D => n13688, CK => CLK, Q => n1743, 
                           QN => n3413);
   REGS_reg_20_18_inst : DFF_X1 port map( D => n13687, CK => CLK, Q => n1744, 
                           QN => n3414);
   REGS_reg_20_17_inst : DFF_X1 port map( D => n13686, CK => CLK, Q => n1745, 
                           QN => n3415);
   REGS_reg_20_16_inst : DFF_X1 port map( D => n13685, CK => CLK, Q => n1746, 
                           QN => n3416);
   REGS_reg_20_15_inst : DFF_X1 port map( D => n13684, CK => CLK, Q => n1747, 
                           QN => n3417);
   REGS_reg_20_14_inst : DFF_X1 port map( D => n13683, CK => CLK, Q => n1748, 
                           QN => n3418);
   REGS_reg_20_13_inst : DFF_X1 port map( D => n13682, CK => CLK, Q => n1749, 
                           QN => n3419);
   REGS_reg_20_12_inst : DFF_X1 port map( D => n13681, CK => CLK, Q => n1750, 
                           QN => n3420);
   REGS_reg_20_11_inst : DFF_X1 port map( D => n13680, CK => CLK, Q => n1751, 
                           QN => n3421);
   REGS_reg_20_10_inst : DFF_X1 port map( D => n13679, CK => CLK, Q => n1752, 
                           QN => n3422);
   REGS_reg_20_9_inst : DFF_X1 port map( D => n13678, CK => CLK, Q => n1753, QN
                           => n3423);
   REGS_reg_20_8_inst : DFF_X1 port map( D => n13677, CK => CLK, Q => n1754, QN
                           => n3424);
   REGS_reg_20_7_inst : DFF_X1 port map( D => n13676, CK => CLK, Q => n1755, QN
                           => n3425);
   REGS_reg_20_6_inst : DFF_X1 port map( D => n13675, CK => CLK, Q => n1756, QN
                           => n3426);
   REGS_reg_20_5_inst : DFF_X1 port map( D => n13674, CK => CLK, Q => n1757, QN
                           => n3427);
   REGS_reg_20_4_inst : DFF_X1 port map( D => n13673, CK => CLK, Q => n1758, QN
                           => n3428);
   REGS_reg_20_3_inst : DFF_X1 port map( D => n13672, CK => CLK, Q => n1759, QN
                           => n3429);
   REGS_reg_20_2_inst : DFF_X1 port map( D => n13671, CK => CLK, Q => n1760, QN
                           => n3430);
   REGS_reg_20_1_inst : DFF_X1 port map( D => n13670, CK => CLK, Q => n1761, QN
                           => n3431);
   REGS_reg_20_0_inst : DFF_X1 port map( D => n13669, CK => CLK, Q => n1762, QN
                           => n3432);
   REGS_reg_19_23_inst : DFF_X1 port map( D => n13724, CK => CLK, Q => n1763, 
                           QN => n3433);
   REGS_reg_19_22_inst : DFF_X1 port map( D => n13723, CK => CLK, Q => n1764, 
                           QN => n3434);
   REGS_reg_19_21_inst : DFF_X1 port map( D => n13722, CK => CLK, Q => n1765, 
                           QN => n3435);
   REGS_reg_19_20_inst : DFF_X1 port map( D => n13721, CK => CLK, Q => n1766, 
                           QN => n3436);
   REGS_reg_19_19_inst : DFF_X1 port map( D => n13720, CK => CLK, Q => n1767, 
                           QN => n3437);
   REGS_reg_19_18_inst : DFF_X1 port map( D => n13719, CK => CLK, Q => n1768, 
                           QN => n3438);
   REGS_reg_19_17_inst : DFF_X1 port map( D => n13718, CK => CLK, Q => n1769, 
                           QN => n3439);
   REGS_reg_19_16_inst : DFF_X1 port map( D => n13717, CK => CLK, Q => n1770, 
                           QN => n3440);
   REGS_reg_19_15_inst : DFF_X1 port map( D => n13716, CK => CLK, Q => n1771, 
                           QN => n3441);
   REGS_reg_19_14_inst : DFF_X1 port map( D => n13715, CK => CLK, Q => n1772, 
                           QN => n3442);
   REGS_reg_19_13_inst : DFF_X1 port map( D => n13714, CK => CLK, Q => n1773, 
                           QN => n3443);
   REGS_reg_19_12_inst : DFF_X1 port map( D => n13713, CK => CLK, Q => n1774, 
                           QN => n3444);
   REGS_reg_19_11_inst : DFF_X1 port map( D => n13712, CK => CLK, Q => n1775, 
                           QN => n3445);
   REGS_reg_19_10_inst : DFF_X1 port map( D => n13711, CK => CLK, Q => n1776, 
                           QN => n3446);
   REGS_reg_19_9_inst : DFF_X1 port map( D => n13710, CK => CLK, Q => n1777, QN
                           => n3447);
   REGS_reg_19_8_inst : DFF_X1 port map( D => n13709, CK => CLK, Q => n1778, QN
                           => n3448);
   REGS_reg_19_7_inst : DFF_X1 port map( D => n13708, CK => CLK, Q => n1779, QN
                           => n3449);
   REGS_reg_19_6_inst : DFF_X1 port map( D => n13707, CK => CLK, Q => n1780, QN
                           => n3450);
   REGS_reg_19_5_inst : DFF_X1 port map( D => n13706, CK => CLK, Q => n1781, QN
                           => n3451);
   REGS_reg_19_4_inst : DFF_X1 port map( D => n13705, CK => CLK, Q => n1782, QN
                           => n3452);
   REGS_reg_19_3_inst : DFF_X1 port map( D => n13704, CK => CLK, Q => n1783, QN
                           => n3453);
   REGS_reg_19_2_inst : DFF_X1 port map( D => n13703, CK => CLK, Q => n1784, QN
                           => n3454);
   REGS_reg_19_1_inst : DFF_X1 port map( D => n13702, CK => CLK, Q => n1785, QN
                           => n3455);
   REGS_reg_19_0_inst : DFF_X1 port map( D => n13701, CK => CLK, Q => n1786, QN
                           => n3456);
   REGS_reg_18_23_inst : DFF_X1 port map( D => n13756, CK => CLK, Q => n_2110, 
                           QN => n52956);
   REGS_reg_18_22_inst : DFF_X1 port map( D => n13755, CK => CLK, Q => n_2111, 
                           QN => n52957);
   REGS_reg_18_21_inst : DFF_X1 port map( D => n13754, CK => CLK, Q => n_2112, 
                           QN => n52958);
   REGS_reg_18_20_inst : DFF_X1 port map( D => n13753, CK => CLK, Q => n_2113, 
                           QN => n52959);
   REGS_reg_18_19_inst : DFF_X1 port map( D => n13752, CK => CLK, Q => n_2114, 
                           QN => n52960);
   REGS_reg_18_18_inst : DFF_X1 port map( D => n13751, CK => CLK, Q => n_2115, 
                           QN => n52961);
   REGS_reg_18_17_inst : DFF_X1 port map( D => n13750, CK => CLK, Q => n_2116, 
                           QN => n52962);
   REGS_reg_18_16_inst : DFF_X1 port map( D => n13749, CK => CLK, Q => n_2117, 
                           QN => n52963);
   REGS_reg_18_15_inst : DFF_X1 port map( D => n13748, CK => CLK, Q => n_2118, 
                           QN => n52964);
   REGS_reg_18_14_inst : DFF_X1 port map( D => n13747, CK => CLK, Q => n_2119, 
                           QN => n52965);
   REGS_reg_18_13_inst : DFF_X1 port map( D => n13746, CK => CLK, Q => n_2120, 
                           QN => n52966);
   REGS_reg_18_12_inst : DFF_X1 port map( D => n13745, CK => CLK, Q => n_2121, 
                           QN => n52967);
   REGS_reg_18_11_inst : DFF_X1 port map( D => n13744, CK => CLK, Q => n_2122, 
                           QN => n52968);
   REGS_reg_18_10_inst : DFF_X1 port map( D => n13743, CK => CLK, Q => n_2123, 
                           QN => n52969);
   REGS_reg_18_9_inst : DFF_X1 port map( D => n13742, CK => CLK, Q => n_2124, 
                           QN => n52970);
   REGS_reg_18_8_inst : DFF_X1 port map( D => n13741, CK => CLK, Q => n_2125, 
                           QN => n52971);
   REGS_reg_18_7_inst : DFF_X1 port map( D => n13740, CK => CLK, Q => n_2126, 
                           QN => n52972);
   REGS_reg_18_6_inst : DFF_X1 port map( D => n13739, CK => CLK, Q => n_2127, 
                           QN => n52973);
   REGS_reg_18_5_inst : DFF_X1 port map( D => n13738, CK => CLK, Q => n_2128, 
                           QN => n52974);
   REGS_reg_18_4_inst : DFF_X1 port map( D => n13737, CK => CLK, Q => n_2129, 
                           QN => n52975);
   REGS_reg_18_3_inst : DFF_X1 port map( D => n13736, CK => CLK, Q => n_2130, 
                           QN => n52976);
   REGS_reg_18_2_inst : DFF_X1 port map( D => n13735, CK => CLK, Q => n_2131, 
                           QN => n52977);
   REGS_reg_18_1_inst : DFF_X1 port map( D => n13734, CK => CLK, Q => n_2132, 
                           QN => n52978);
   REGS_reg_18_0_inst : DFF_X1 port map( D => n13733, CK => CLK, Q => n_2133, 
                           QN => n52979);
   REGS_reg_17_23_inst : DFF_X1 port map( D => n13788, CK => CLK, Q => n_2134, 
                           QN => n52980);
   REGS_reg_17_22_inst : DFF_X1 port map( D => n13787, CK => CLK, Q => n_2135, 
                           QN => n52981);
   REGS_reg_17_21_inst : DFF_X1 port map( D => n13786, CK => CLK, Q => n_2136, 
                           QN => n52982);
   REGS_reg_17_20_inst : DFF_X1 port map( D => n13785, CK => CLK, Q => n_2137, 
                           QN => n52983);
   REGS_reg_17_19_inst : DFF_X1 port map( D => n13784, CK => CLK, Q => n_2138, 
                           QN => n52984);
   REGS_reg_17_18_inst : DFF_X1 port map( D => n13783, CK => CLK, Q => n_2139, 
                           QN => n52985);
   REGS_reg_17_17_inst : DFF_X1 port map( D => n13782, CK => CLK, Q => n_2140, 
                           QN => n52986);
   REGS_reg_17_16_inst : DFF_X1 port map( D => n13781, CK => CLK, Q => n_2141, 
                           QN => n52987);
   REGS_reg_17_15_inst : DFF_X1 port map( D => n13780, CK => CLK, Q => n_2142, 
                           QN => n52988);
   REGS_reg_17_14_inst : DFF_X1 port map( D => n13779, CK => CLK, Q => n_2143, 
                           QN => n52989);
   REGS_reg_17_13_inst : DFF_X1 port map( D => n13778, CK => CLK, Q => n_2144, 
                           QN => n52990);
   REGS_reg_17_12_inst : DFF_X1 port map( D => n13777, CK => CLK, Q => n_2145, 
                           QN => n52991);
   REGS_reg_17_11_inst : DFF_X1 port map( D => n13776, CK => CLK, Q => n_2146, 
                           QN => n52992);
   REGS_reg_17_10_inst : DFF_X1 port map( D => n13775, CK => CLK, Q => n_2147, 
                           QN => n52993);
   REGS_reg_17_9_inst : DFF_X1 port map( D => n13774, CK => CLK, Q => n_2148, 
                           QN => n52994);
   REGS_reg_17_8_inst : DFF_X1 port map( D => n13773, CK => CLK, Q => n_2149, 
                           QN => n52995);
   REGS_reg_17_7_inst : DFF_X1 port map( D => n13772, CK => CLK, Q => n_2150, 
                           QN => n52996);
   REGS_reg_17_6_inst : DFF_X1 port map( D => n13771, CK => CLK, Q => n_2151, 
                           QN => n52997);
   REGS_reg_17_5_inst : DFF_X1 port map( D => n13770, CK => CLK, Q => n_2152, 
                           QN => n52998);
   REGS_reg_17_4_inst : DFF_X1 port map( D => n13769, CK => CLK, Q => n_2153, 
                           QN => n52999);
   REGS_reg_17_3_inst : DFF_X1 port map( D => n13768, CK => CLK, Q => n_2154, 
                           QN => n53000);
   REGS_reg_17_2_inst : DFF_X1 port map( D => n13767, CK => CLK, Q => n_2155, 
                           QN => n53001);
   REGS_reg_17_1_inst : DFF_X1 port map( D => n13766, CK => CLK, Q => n_2156, 
                           QN => n53002);
   REGS_reg_17_0_inst : DFF_X1 port map( D => n13765, CK => CLK, Q => n_2157, 
                           QN => n53003);
   REGS_reg_16_23_inst : DFF_X1 port map( D => n13820, CK => CLK, Q => n4379, 
                           QN => n568);
   REGS_reg_16_22_inst : DFF_X1 port map( D => n13819, CK => CLK, Q => n4380, 
                           QN => n569);
   REGS_reg_16_21_inst : DFF_X1 port map( D => n13818, CK => CLK, Q => n4381, 
                           QN => n570);
   REGS_reg_16_20_inst : DFF_X1 port map( D => n13817, CK => CLK, Q => n4382, 
                           QN => n571);
   REGS_reg_16_19_inst : DFF_X1 port map( D => n13816, CK => CLK, Q => n4383, 
                           QN => n572);
   REGS_reg_16_18_inst : DFF_X1 port map( D => n13815, CK => CLK, Q => n4384, 
                           QN => n573);
   REGS_reg_16_17_inst : DFF_X1 port map( D => n13814, CK => CLK, Q => n4385, 
                           QN => n574);
   REGS_reg_16_16_inst : DFF_X1 port map( D => n13813, CK => CLK, Q => n4386, 
                           QN => n575);
   REGS_reg_16_15_inst : DFF_X1 port map( D => n13812, CK => CLK, Q => n4387, 
                           QN => n576);
   REGS_reg_16_14_inst : DFF_X1 port map( D => n13811, CK => CLK, Q => n4388, 
                           QN => n577);
   REGS_reg_16_13_inst : DFF_X1 port map( D => n13810, CK => CLK, Q => n4389, 
                           QN => n578);
   REGS_reg_16_12_inst : DFF_X1 port map( D => n13809, CK => CLK, Q => n4390, 
                           QN => n579);
   REGS_reg_16_11_inst : DFF_X1 port map( D => n13808, CK => CLK, Q => n4391, 
                           QN => n580);
   REGS_reg_16_10_inst : DFF_X1 port map( D => n13807, CK => CLK, Q => n4392, 
                           QN => n581);
   REGS_reg_16_9_inst : DFF_X1 port map( D => n13806, CK => CLK, Q => n4393, QN
                           => n582);
   REGS_reg_16_8_inst : DFF_X1 port map( D => n13805, CK => CLK, Q => n4394, QN
                           => n583);
   REGS_reg_16_7_inst : DFF_X1 port map( D => n13804, CK => CLK, Q => n4395, QN
                           => n584);
   REGS_reg_16_6_inst : DFF_X1 port map( D => n13803, CK => CLK, Q => n4396, QN
                           => n585);
   REGS_reg_16_5_inst : DFF_X1 port map( D => n13802, CK => CLK, Q => n4397, QN
                           => n586);
   REGS_reg_16_4_inst : DFF_X1 port map( D => n13801, CK => CLK, Q => n4398, QN
                           => n587);
   REGS_reg_16_3_inst : DFF_X1 port map( D => n13800, CK => CLK, Q => n4399, QN
                           => n588);
   REGS_reg_16_2_inst : DFF_X1 port map( D => n13799, CK => CLK, Q => n4400, QN
                           => n589);
   REGS_reg_16_1_inst : DFF_X1 port map( D => n13798, CK => CLK, Q => n4401, QN
                           => n590);
   REGS_reg_16_0_inst : DFF_X1 port map( D => n13797, CK => CLK, Q => n4402, QN
                           => n591);
   REGS_reg_63_23_inst : DFF_X1 port map( D => n12316, CK => CLK, Q => n_2158, 
                           QN => n1669);
   REGS_reg_63_22_inst : DFF_X1 port map( D => n12315, CK => CLK, Q => n_2159, 
                           QN => n1670);
   REGS_reg_63_21_inst : DFF_X1 port map( D => n12314, CK => CLK, Q => n_2160, 
                           QN => n1671);
   REGS_reg_63_20_inst : DFF_X1 port map( D => n12313, CK => CLK, Q => n_2161, 
                           QN => n1672);
   REGS_reg_63_19_inst : DFF_X1 port map( D => n12312, CK => CLK, Q => n_2162, 
                           QN => n1673);
   REGS_reg_63_18_inst : DFF_X1 port map( D => n12311, CK => CLK, Q => n_2163, 
                           QN => n1674);
   REGS_reg_63_17_inst : DFF_X1 port map( D => n12310, CK => CLK, Q => n_2164, 
                           QN => n1675);
   REGS_reg_63_16_inst : DFF_X1 port map( D => n12309, CK => CLK, Q => n_2165, 
                           QN => n1676);
   REGS_reg_63_15_inst : DFF_X1 port map( D => n12308, CK => CLK, Q => n_2166, 
                           QN => n1677);
   REGS_reg_63_14_inst : DFF_X1 port map( D => n12307, CK => CLK, Q => n_2167, 
                           QN => n1678);
   REGS_reg_63_13_inst : DFF_X1 port map( D => n12306, CK => CLK, Q => n_2168, 
                           QN => n1679);
   REGS_reg_63_12_inst : DFF_X1 port map( D => n12305, CK => CLK, Q => n_2169, 
                           QN => n1680);
   REGS_reg_63_11_inst : DFF_X1 port map( D => n12304, CK => CLK, Q => n_2170, 
                           QN => n1681);
   REGS_reg_63_10_inst : DFF_X1 port map( D => n12303, CK => CLK, Q => n_2171, 
                           QN => n1682);
   REGS_reg_63_9_inst : DFF_X1 port map( D => n12302, CK => CLK, Q => n_2172, 
                           QN => n1683);
   REGS_reg_63_8_inst : DFF_X1 port map( D => n12301, CK => CLK, Q => n_2173, 
                           QN => n1684);
   REGS_reg_63_7_inst : DFF_X1 port map( D => n12300, CK => CLK, Q => n_2174, 
                           QN => n1685);
   REGS_reg_63_6_inst : DFF_X1 port map( D => n12299, CK => CLK, Q => n_2175, 
                           QN => n1686);
   REGS_reg_63_5_inst : DFF_X1 port map( D => n12298, CK => CLK, Q => n_2176, 
                           QN => n1687);
   REGS_reg_63_4_inst : DFF_X1 port map( D => n12297, CK => CLK, Q => n_2177, 
                           QN => n1688);
   REGS_reg_63_3_inst : DFF_X1 port map( D => n12296, CK => CLK, Q => n_2178, 
                           QN => n1689);
   REGS_reg_63_2_inst : DFF_X1 port map( D => n12295, CK => CLK, Q => n_2179, 
                           QN => n1690);
   REGS_reg_63_1_inst : DFF_X1 port map( D => n12294, CK => CLK, Q => n_2180, 
                           QN => n1691);
   REGS_reg_63_0_inst : DFF_X1 port map( D => n12293, CK => CLK, Q => n_2181, 
                           QN => n1692);
   REGS_reg_60_23_inst : DFF_X1 port map( D => n12412, CK => CLK, Q => n_2182, 
                           QN => n53028);
   REGS_reg_60_22_inst : DFF_X1 port map( D => n12411, CK => CLK, Q => n_2183, 
                           QN => n53029);
   REGS_reg_60_21_inst : DFF_X1 port map( D => n12410, CK => CLK, Q => n_2184, 
                           QN => n53030);
   REGS_reg_60_20_inst : DFF_X1 port map( D => n12409, CK => CLK, Q => n_2185, 
                           QN => n53031);
   REGS_reg_60_19_inst : DFF_X1 port map( D => n12408, CK => CLK, Q => n_2186, 
                           QN => n53032);
   REGS_reg_60_18_inst : DFF_X1 port map( D => n12407, CK => CLK, Q => n_2187, 
                           QN => n53033);
   REGS_reg_60_17_inst : DFF_X1 port map( D => n12406, CK => CLK, Q => n_2188, 
                           QN => n53034);
   REGS_reg_60_16_inst : DFF_X1 port map( D => n12405, CK => CLK, Q => n_2189, 
                           QN => n53035);
   REGS_reg_60_15_inst : DFF_X1 port map( D => n12404, CK => CLK, Q => n_2190, 
                           QN => n53036);
   REGS_reg_60_14_inst : DFF_X1 port map( D => n12403, CK => CLK, Q => n_2191, 
                           QN => n53037);
   REGS_reg_60_13_inst : DFF_X1 port map( D => n12402, CK => CLK, Q => n_2192, 
                           QN => n53038);
   REGS_reg_60_12_inst : DFF_X1 port map( D => n12401, CK => CLK, Q => n_2193, 
                           QN => n53039);
   REGS_reg_60_11_inst : DFF_X1 port map( D => n12400, CK => CLK, Q => n_2194, 
                           QN => n53040);
   REGS_reg_60_10_inst : DFF_X1 port map( D => n12399, CK => CLK, Q => n_2195, 
                           QN => n53041);
   REGS_reg_60_9_inst : DFF_X1 port map( D => n12398, CK => CLK, Q => n_2196, 
                           QN => n53042);
   REGS_reg_60_8_inst : DFF_X1 port map( D => n12397, CK => CLK, Q => n_2197, 
                           QN => n53043);
   REGS_reg_60_7_inst : DFF_X1 port map( D => n12396, CK => CLK, Q => n_2198, 
                           QN => n53044);
   REGS_reg_60_6_inst : DFF_X1 port map( D => n12395, CK => CLK, Q => n_2199, 
                           QN => n53045);
   REGS_reg_60_5_inst : DFF_X1 port map( D => n12394, CK => CLK, Q => n_2200, 
                           QN => n53046);
   REGS_reg_60_4_inst : DFF_X1 port map( D => n12393, CK => CLK, Q => n_2201, 
                           QN => n53047);
   REGS_reg_60_3_inst : DFF_X1 port map( D => n12392, CK => CLK, Q => n_2202, 
                           QN => n53048);
   REGS_reg_60_2_inst : DFF_X1 port map( D => n12391, CK => CLK, Q => n_2203, 
                           QN => n53049);
   REGS_reg_60_1_inst : DFF_X1 port map( D => n12390, CK => CLK, Q => n_2204, 
                           QN => n53050);
   REGS_reg_60_0_inst : DFF_X1 port map( D => n12389, CK => CLK, Q => n_2205, 
                           QN => n53051);
   REGS_reg_49_23_inst : DFF_X1 port map( D => n12764, CK => CLK, Q => n4786, 
                           QN => n53148);
   REGS_reg_49_22_inst : DFF_X1 port map( D => n12763, CK => CLK, Q => n4787, 
                           QN => n53149);
   REGS_reg_49_21_inst : DFF_X1 port map( D => n12762, CK => CLK, Q => n4788, 
                           QN => n53150);
   REGS_reg_49_20_inst : DFF_X1 port map( D => n12761, CK => CLK, Q => n4789, 
                           QN => n53151);
   REGS_reg_49_19_inst : DFF_X1 port map( D => n12760, CK => CLK, Q => n4790, 
                           QN => n53152);
   REGS_reg_49_18_inst : DFF_X1 port map( D => n12759, CK => CLK, Q => n4791, 
                           QN => n53153);
   REGS_reg_49_17_inst : DFF_X1 port map( D => n12758, CK => CLK, Q => n4792, 
                           QN => n53154);
   REGS_reg_49_16_inst : DFF_X1 port map( D => n12757, CK => CLK, Q => n4793, 
                           QN => n53155);
   REGS_reg_49_15_inst : DFF_X1 port map( D => n12756, CK => CLK, Q => n4794, 
                           QN => n53156);
   REGS_reg_49_14_inst : DFF_X1 port map( D => n12755, CK => CLK, Q => n4795, 
                           QN => n53157);
   REGS_reg_49_13_inst : DFF_X1 port map( D => n12754, CK => CLK, Q => n4796, 
                           QN => n53158);
   REGS_reg_49_12_inst : DFF_X1 port map( D => n12753, CK => CLK, Q => n4797, 
                           QN => n53159);
   REGS_reg_49_11_inst : DFF_X1 port map( D => n12752, CK => CLK, Q => n4798, 
                           QN => n53160);
   REGS_reg_49_10_inst : DFF_X1 port map( D => n12751, CK => CLK, Q => n4799, 
                           QN => n53161);
   REGS_reg_49_9_inst : DFF_X1 port map( D => n12750, CK => CLK, Q => n4800, QN
                           => n53162);
   REGS_reg_49_8_inst : DFF_X1 port map( D => n12749, CK => CLK, Q => n4801, QN
                           => n53163);
   REGS_reg_49_7_inst : DFF_X1 port map( D => n12748, CK => CLK, Q => n4802, QN
                           => n53164);
   REGS_reg_49_6_inst : DFF_X1 port map( D => n12747, CK => CLK, Q => n4803, QN
                           => n53165);
   REGS_reg_49_5_inst : DFF_X1 port map( D => n12746, CK => CLK, Q => n4804, QN
                           => n53166);
   REGS_reg_49_4_inst : DFF_X1 port map( D => n12745, CK => CLK, Q => n4805, QN
                           => n53167);
   REGS_reg_49_3_inst : DFF_X1 port map( D => n12744, CK => CLK, Q => n4806, QN
                           => n53168);
   REGS_reg_49_2_inst : DFF_X1 port map( D => n12743, CK => CLK, Q => n4807, QN
                           => n53169);
   REGS_reg_49_1_inst : DFF_X1 port map( D => n12742, CK => CLK, Q => n4808, QN
                           => n53170);
   REGS_reg_49_0_inst : DFF_X1 port map( D => n12741, CK => CLK, Q => n4809, QN
                           => n53171);
   REGS_reg_48_23_inst : DFF_X1 port map( D => n12796, CK => CLK, Q => n4810, 
                           QN => n53172);
   REGS_reg_48_22_inst : DFF_X1 port map( D => n12795, CK => CLK, Q => n4811, 
                           QN => n53173);
   REGS_reg_48_21_inst : DFF_X1 port map( D => n12794, CK => CLK, Q => n4812, 
                           QN => n53174);
   REGS_reg_48_20_inst : DFF_X1 port map( D => n12793, CK => CLK, Q => n4813, 
                           QN => n53175);
   REGS_reg_48_19_inst : DFF_X1 port map( D => n12792, CK => CLK, Q => n4814, 
                           QN => n53176);
   REGS_reg_48_18_inst : DFF_X1 port map( D => n12791, CK => CLK, Q => n4815, 
                           QN => n53177);
   REGS_reg_48_17_inst : DFF_X1 port map( D => n12790, CK => CLK, Q => n4816, 
                           QN => n53178);
   REGS_reg_48_16_inst : DFF_X1 port map( D => n12789, CK => CLK, Q => n4817, 
                           QN => n53179);
   REGS_reg_48_15_inst : DFF_X1 port map( D => n12788, CK => CLK, Q => n4818, 
                           QN => n53180);
   REGS_reg_48_14_inst : DFF_X1 port map( D => n12787, CK => CLK, Q => n4819, 
                           QN => n53181);
   REGS_reg_48_13_inst : DFF_X1 port map( D => n12786, CK => CLK, Q => n4820, 
                           QN => n53182);
   REGS_reg_48_12_inst : DFF_X1 port map( D => n12785, CK => CLK, Q => n4821, 
                           QN => n53183);
   REGS_reg_48_11_inst : DFF_X1 port map( D => n12784, CK => CLK, Q => n4822, 
                           QN => n53184);
   REGS_reg_48_10_inst : DFF_X1 port map( D => n12783, CK => CLK, Q => n4823, 
                           QN => n53185);
   REGS_reg_44_23_inst : DFF_X1 port map( D => n12924, CK => CLK, Q => n_2206, 
                           QN => n53244);
   REGS_reg_44_22_inst : DFF_X1 port map( D => n12923, CK => CLK, Q => n_2207, 
                           QN => n53245);
   REGS_reg_44_21_inst : DFF_X1 port map( D => n12922, CK => CLK, Q => n_2208, 
                           QN => n53246);
   REGS_reg_44_20_inst : DFF_X1 port map( D => n12921, CK => CLK, Q => n_2209, 
                           QN => n53247);
   REGS_reg_44_19_inst : DFF_X1 port map( D => n12920, CK => CLK, Q => n_2210, 
                           QN => n53248);
   REGS_reg_44_18_inst : DFF_X1 port map( D => n12919, CK => CLK, Q => n_2211, 
                           QN => n53249);
   REGS_reg_44_17_inst : DFF_X1 port map( D => n12918, CK => CLK, Q => n_2212, 
                           QN => n53250);
   REGS_reg_44_16_inst : DFF_X1 port map( D => n12917, CK => CLK, Q => n_2213, 
                           QN => n53251);
   REGS_reg_44_15_inst : DFF_X1 port map( D => n12916, CK => CLK, Q => n_2214, 
                           QN => n53252);
   REGS_reg_44_14_inst : DFF_X1 port map( D => n12915, CK => CLK, Q => n_2215, 
                           QN => n53253);
   REGS_reg_44_13_inst : DFF_X1 port map( D => n12914, CK => CLK, Q => n_2216, 
                           QN => n53254);
   REGS_reg_44_12_inst : DFF_X1 port map( D => n12913, CK => CLK, Q => n_2217, 
                           QN => n53255);
   REGS_reg_44_11_inst : DFF_X1 port map( D => n12912, CK => CLK, Q => n_2218, 
                           QN => n53256);
   REGS_reg_44_10_inst : DFF_X1 port map( D => n12911, CK => CLK, Q => n_2219, 
                           QN => n53257);
   REGS_reg_39_23_inst : DFF_X1 port map( D => n13084, CK => CLK, Q => n4906, 
                           QN => n9787);
   REGS_reg_39_22_inst : DFF_X1 port map( D => n13083, CK => CLK, Q => n4907, 
                           QN => n9788);
   REGS_reg_39_21_inst : DFF_X1 port map( D => n13082, CK => CLK, Q => n4908, 
                           QN => n9789);
   REGS_reg_39_20_inst : DFF_X1 port map( D => n13081, CK => CLK, Q => n4909, 
                           QN => n9790);
   REGS_reg_39_19_inst : DFF_X1 port map( D => n13080, CK => CLK, Q => n4910, 
                           QN => n9791);
   REGS_reg_39_18_inst : DFF_X1 port map( D => n13079, CK => CLK, Q => n4911, 
                           QN => n9792);
   REGS_reg_39_17_inst : DFF_X1 port map( D => n13078, CK => CLK, Q => n4912, 
                           QN => n9793);
   REGS_reg_39_16_inst : DFF_X1 port map( D => n13077, CK => CLK, Q => n4913, 
                           QN => n9794);
   REGS_reg_39_15_inst : DFF_X1 port map( D => n13076, CK => CLK, Q => n4914, 
                           QN => n9795);
   REGS_reg_39_14_inst : DFF_X1 port map( D => n13075, CK => CLK, Q => n4915, 
                           QN => n9796);
   REGS_reg_39_13_inst : DFF_X1 port map( D => n13074, CK => CLK, Q => n4916, 
                           QN => n9797);
   REGS_reg_39_12_inst : DFF_X1 port map( D => n13073, CK => CLK, Q => n4917, 
                           QN => n9798);
   REGS_reg_39_11_inst : DFF_X1 port map( D => n13072, CK => CLK, Q => n4918, 
                           QN => n9799);
   REGS_reg_39_10_inst : DFF_X1 port map( D => n13071, CK => CLK, Q => n4919, 
                           QN => n9800);
   REGS_reg_39_9_inst : DFF_X1 port map( D => n13070, CK => CLK, Q => n4920, QN
                           => n9801);
   REGS_reg_39_8_inst : DFF_X1 port map( D => n13069, CK => CLK, Q => n4921, QN
                           => n9802);
   REGS_reg_39_7_inst : DFF_X1 port map( D => n13068, CK => CLK, Q => n4922, QN
                           => n9803);
   REGS_reg_39_6_inst : DFF_X1 port map( D => n13067, CK => CLK, Q => n4923, QN
                           => n9804);
   REGS_reg_39_5_inst : DFF_X1 port map( D => n13066, CK => CLK, Q => n4924, QN
                           => n9805);
   REGS_reg_39_4_inst : DFF_X1 port map( D => n13065, CK => CLK, Q => n4925, QN
                           => n9806);
   REGS_reg_39_3_inst : DFF_X1 port map( D => n13064, CK => CLK, Q => n4926, QN
                           => n9807);
   REGS_reg_39_2_inst : DFF_X1 port map( D => n13063, CK => CLK, Q => n4927, QN
                           => n9808);
   REGS_reg_39_1_inst : DFF_X1 port map( D => n13062, CK => CLK, Q => n4928, QN
                           => n9809);
   REGS_reg_39_0_inst : DFF_X1 port map( D => n13061, CK => CLK, Q => n4929, QN
                           => n9810);
   REGS_reg_38_23_inst : DFF_X1 port map( D => n13116, CK => CLK, Q => n4930, 
                           QN => n9755);
   REGS_reg_38_22_inst : DFF_X1 port map( D => n13115, CK => CLK, Q => n4931, 
                           QN => n9756);
   REGS_reg_38_21_inst : DFF_X1 port map( D => n13114, CK => CLK, Q => n4932, 
                           QN => n9757);
   REGS_reg_38_20_inst : DFF_X1 port map( D => n13113, CK => CLK, Q => n4933, 
                           QN => n9758);
   REGS_reg_38_19_inst : DFF_X1 port map( D => n13112, CK => CLK, Q => n4934, 
                           QN => n9759);
   REGS_reg_38_18_inst : DFF_X1 port map( D => n13111, CK => CLK, Q => n4935, 
                           QN => n9760);
   REGS_reg_38_17_inst : DFF_X1 port map( D => n13110, CK => CLK, Q => n4936, 
                           QN => n9761);
   REGS_reg_38_16_inst : DFF_X1 port map( D => n13109, CK => CLK, Q => n4937, 
                           QN => n9762);
   REGS_reg_38_15_inst : DFF_X1 port map( D => n13108, CK => CLK, Q => n4938, 
                           QN => n9763);
   REGS_reg_38_14_inst : DFF_X1 port map( D => n13107, CK => CLK, Q => n4939, 
                           QN => n9764);
   REGS_reg_38_13_inst : DFF_X1 port map( D => n13106, CK => CLK, Q => n4940, 
                           QN => n9765);
   REGS_reg_38_12_inst : DFF_X1 port map( D => n13105, CK => CLK, Q => n4941, 
                           QN => n9766);
   REGS_reg_38_11_inst : DFF_X1 port map( D => n13104, CK => CLK, Q => n4942, 
                           QN => n9767);
   REGS_reg_38_10_inst : DFF_X1 port map( D => n13103, CK => CLK, Q => n4943, 
                           QN => n9768);
   REGS_reg_38_9_inst : DFF_X1 port map( D => n13102, CK => CLK, Q => n4944, QN
                           => n9769);
   REGS_reg_38_8_inst : DFF_X1 port map( D => n13101, CK => CLK, Q => n4945, QN
                           => n9770);
   REGS_reg_38_7_inst : DFF_X1 port map( D => n13100, CK => CLK, Q => n4946, QN
                           => n9771);
   REGS_reg_38_6_inst : DFF_X1 port map( D => n13099, CK => CLK, Q => n4947, QN
                           => n9772);
   REGS_reg_38_5_inst : DFF_X1 port map( D => n13098, CK => CLK, Q => n4948, QN
                           => n9773);
   REGS_reg_38_4_inst : DFF_X1 port map( D => n13097, CK => CLK, Q => n4949, QN
                           => n9774);
   REGS_reg_38_3_inst : DFF_X1 port map( D => n13096, CK => CLK, Q => n4950, QN
                           => n9775);
   REGS_reg_38_2_inst : DFF_X1 port map( D => n13095, CK => CLK, Q => n4951, QN
                           => n9776);
   REGS_reg_38_1_inst : DFF_X1 port map( D => n13094, CK => CLK, Q => n4952, QN
                           => n9777);
   REGS_reg_38_0_inst : DFF_X1 port map( D => n13093, CK => CLK, Q => n4953, QN
                           => n9778);
   REGS_reg_37_23_inst : DFF_X1 port map( D => n13148, CK => CLK, Q => n_2220, 
                           QN => n3621);
   REGS_reg_37_22_inst : DFF_X1 port map( D => n13147, CK => CLK, Q => n_2221, 
                           QN => n3622);
   REGS_reg_37_21_inst : DFF_X1 port map( D => n13146, CK => CLK, Q => n_2222, 
                           QN => n3623);
   REGS_reg_37_20_inst : DFF_X1 port map( D => n13145, CK => CLK, Q => n_2223, 
                           QN => n3624);
   REGS_reg_37_19_inst : DFF_X1 port map( D => n13144, CK => CLK, Q => n_2224, 
                           QN => n3625);
   REGS_reg_37_18_inst : DFF_X1 port map( D => n13143, CK => CLK, Q => n_2225, 
                           QN => n3626);
   REGS_reg_37_17_inst : DFF_X1 port map( D => n13142, CK => CLK, Q => n_2226, 
                           QN => n3627);
   REGS_reg_37_16_inst : DFF_X1 port map( D => n13141, CK => CLK, Q => n_2227, 
                           QN => n3628);
   REGS_reg_37_15_inst : DFF_X1 port map( D => n13140, CK => CLK, Q => n_2228, 
                           QN => n3629);
   REGS_reg_37_14_inst : DFF_X1 port map( D => n13139, CK => CLK, Q => n_2229, 
                           QN => n3630);
   REGS_reg_37_13_inst : DFF_X1 port map( D => n13138, CK => CLK, Q => n_2230, 
                           QN => n3631);
   REGS_reg_37_12_inst : DFF_X1 port map( D => n13137, CK => CLK, Q => n_2231, 
                           QN => n3632);
   REGS_reg_37_11_inst : DFF_X1 port map( D => n13136, CK => CLK, Q => n_2232, 
                           QN => n3633);
   REGS_reg_37_10_inst : DFF_X1 port map( D => n13135, CK => CLK, Q => n_2233, 
                           QN => n3634);
   REGS_reg_37_9_inst : DFF_X1 port map( D => n13134, CK => CLK, Q => n_2234, 
                           QN => n3635);
   REGS_reg_37_8_inst : DFF_X1 port map( D => n13133, CK => CLK, Q => n_2235, 
                           QN => n3636);
   REGS_reg_37_7_inst : DFF_X1 port map( D => n13132, CK => CLK, Q => n_2236, 
                           QN => n3637);
   REGS_reg_37_6_inst : DFF_X1 port map( D => n13131, CK => CLK, Q => n_2237, 
                           QN => n3638);
   REGS_reg_37_5_inst : DFF_X1 port map( D => n13130, CK => CLK, Q => n_2238, 
                           QN => n3639);
   REGS_reg_37_4_inst : DFF_X1 port map( D => n13129, CK => CLK, Q => n_2239, 
                           QN => n3640);
   REGS_reg_37_3_inst : DFF_X1 port map( D => n13128, CK => CLK, Q => n_2240, 
                           QN => n3641);
   REGS_reg_37_2_inst : DFF_X1 port map( D => n13127, CK => CLK, Q => n_2241, 
                           QN => n3642);
   REGS_reg_37_1_inst : DFF_X1 port map( D => n13126, CK => CLK, Q => n_2242, 
                           QN => n3643);
   REGS_reg_37_0_inst : DFF_X1 port map( D => n13125, CK => CLK, Q => n_2243, 
                           QN => n3644);
   REGS_reg_36_23_inst : DFF_X1 port map( D => n13180, CK => CLK, Q => n_2244, 
                           QN => n1999);
   REGS_reg_36_22_inst : DFF_X1 port map( D => n13179, CK => CLK, Q => n_2245, 
                           QN => n2000);
   REGS_reg_36_21_inst : DFF_X1 port map( D => n13178, CK => CLK, Q => n_2246, 
                           QN => n2001);
   REGS_reg_36_20_inst : DFF_X1 port map( D => n13177, CK => CLK, Q => n_2247, 
                           QN => n2002);
   REGS_reg_36_19_inst : DFF_X1 port map( D => n13176, CK => CLK, Q => n_2248, 
                           QN => n2003);
   REGS_reg_36_18_inst : DFF_X1 port map( D => n13175, CK => CLK, Q => n_2249, 
                           QN => n2004);
   REGS_reg_36_17_inst : DFF_X1 port map( D => n13174, CK => CLK, Q => n_2250, 
                           QN => n2005);
   REGS_reg_36_16_inst : DFF_X1 port map( D => n13173, CK => CLK, Q => n_2251, 
                           QN => n2006);
   REGS_reg_36_15_inst : DFF_X1 port map( D => n13172, CK => CLK, Q => n_2252, 
                           QN => n2007);
   REGS_reg_36_14_inst : DFF_X1 port map( D => n13171, CK => CLK, Q => n_2253, 
                           QN => n2008);
   REGS_reg_36_13_inst : DFF_X1 port map( D => n13170, CK => CLK, Q => n_2254, 
                           QN => n2009);
   REGS_reg_36_12_inst : DFF_X1 port map( D => n13169, CK => CLK, Q => n_2255, 
                           QN => n2010);
   REGS_reg_36_11_inst : DFF_X1 port map( D => n13168, CK => CLK, Q => n_2256, 
                           QN => n2011);
   REGS_reg_36_10_inst : DFF_X1 port map( D => n13167, CK => CLK, Q => n_2257, 
                           QN => n2012);
   REGS_reg_36_9_inst : DFF_X1 port map( D => n13166, CK => CLK, Q => n_2258, 
                           QN => n2013);
   REGS_reg_36_8_inst : DFF_X1 port map( D => n13165, CK => CLK, Q => n_2259, 
                           QN => n2014);
   REGS_reg_36_7_inst : DFF_X1 port map( D => n13164, CK => CLK, Q => n_2260, 
                           QN => n2015);
   REGS_reg_36_6_inst : DFF_X1 port map( D => n13163, CK => CLK, Q => n_2261, 
                           QN => n2016);
   REGS_reg_36_5_inst : DFF_X1 port map( D => n13162, CK => CLK, Q => n_2262, 
                           QN => n2017);
   REGS_reg_36_4_inst : DFF_X1 port map( D => n13161, CK => CLK, Q => n_2263, 
                           QN => n2018);
   REGS_reg_36_3_inst : DFF_X1 port map( D => n13160, CK => CLK, Q => n_2264, 
                           QN => n2019);
   REGS_reg_36_2_inst : DFF_X1 port map( D => n13159, CK => CLK, Q => n_2265, 
                           QN => n2020);
   REGS_reg_36_1_inst : DFF_X1 port map( D => n13158, CK => CLK, Q => n_2266, 
                           QN => n2021);
   REGS_reg_36_0_inst : DFF_X1 port map( D => n13157, CK => CLK, Q => n_2267, 
                           QN => n2022);
   REGS_reg_33_23_inst : DFF_X1 port map( D => n13276, CK => CLK, Q => n5002, 
                           QN => n53356);
   REGS_reg_33_22_inst : DFF_X1 port map( D => n13275, CK => CLK, Q => n5003, 
                           QN => n53357);
   REGS_reg_33_21_inst : DFF_X1 port map( D => n13274, CK => CLK, Q => n5004, 
                           QN => n53358);
   REGS_reg_33_20_inst : DFF_X1 port map( D => n13273, CK => CLK, Q => n5005, 
                           QN => n53359);
   REGS_reg_33_19_inst : DFF_X1 port map( D => n13272, CK => CLK, Q => n5006, 
                           QN => n53360);
   REGS_reg_33_18_inst : DFF_X1 port map( D => n13271, CK => CLK, Q => n5007, 
                           QN => n53361);
   REGS_reg_33_17_inst : DFF_X1 port map( D => n13270, CK => CLK, Q => n5008, 
                           QN => n53362);
   REGS_reg_33_16_inst : DFF_X1 port map( D => n13269, CK => CLK, Q => n5009, 
                           QN => n53363);
   REGS_reg_33_15_inst : DFF_X1 port map( D => n13268, CK => CLK, Q => n5010, 
                           QN => n53364);
   REGS_reg_33_14_inst : DFF_X1 port map( D => n13267, CK => CLK, Q => n5011, 
                           QN => n53365);
   REGS_reg_33_13_inst : DFF_X1 port map( D => n13266, CK => CLK, Q => n5012, 
                           QN => n53366);
   REGS_reg_33_12_inst : DFF_X1 port map( D => n13265, CK => CLK, Q => n5013, 
                           QN => n53367);
   REGS_reg_33_11_inst : DFF_X1 port map( D => n13264, CK => CLK, Q => n5014, 
                           QN => n53368);
   REGS_reg_33_10_inst : DFF_X1 port map( D => n13263, CK => CLK, Q => n5015, 
                           QN => n53369);
   REGS_reg_33_9_inst : DFF_X1 port map( D => n13262, CK => CLK, Q => n5016, QN
                           => n53370);
   REGS_reg_33_8_inst : DFF_X1 port map( D => n13261, CK => CLK, Q => n5017, QN
                           => n53371);
   REGS_reg_33_7_inst : DFF_X1 port map( D => n13260, CK => CLK, Q => n5018, QN
                           => n53372);
   REGS_reg_33_6_inst : DFF_X1 port map( D => n13259, CK => CLK, Q => n5019, QN
                           => n53373);
   REGS_reg_33_5_inst : DFF_X1 port map( D => n13258, CK => CLK, Q => n5020, QN
                           => n53374);
   REGS_reg_33_4_inst : DFF_X1 port map( D => n13257, CK => CLK, Q => n5021, QN
                           => n53375);
   REGS_reg_33_3_inst : DFF_X1 port map( D => n13256, CK => CLK, Q => n5022, QN
                           => n53376);
   REGS_reg_33_2_inst : DFF_X1 port map( D => n13255, CK => CLK, Q => n5023, QN
                           => n53377);
   REGS_reg_33_1_inst : DFF_X1 port map( D => n13254, CK => CLK, Q => n5024, QN
                           => n53378);
   REGS_reg_33_0_inst : DFF_X1 port map( D => n13253, CK => CLK, Q => n5025, QN
                           => n53379);
   REGS_reg_32_23_inst : DFF_X1 port map( D => n13308, CK => CLK, Q => n5026, 
                           QN => n53380);
   REGS_reg_32_22_inst : DFF_X1 port map( D => n13307, CK => CLK, Q => n5027, 
                           QN => n53381);
   REGS_reg_32_21_inst : DFF_X1 port map( D => n13306, CK => CLK, Q => n5028, 
                           QN => n53382);
   REGS_reg_32_20_inst : DFF_X1 port map( D => n13305, CK => CLK, Q => n5029, 
                           QN => n53383);
   REGS_reg_32_19_inst : DFF_X1 port map( D => n13304, CK => CLK, Q => n5030, 
                           QN => n53384);
   REGS_reg_32_18_inst : DFF_X1 port map( D => n13303, CK => CLK, Q => n5031, 
                           QN => n53385);
   REGS_reg_32_17_inst : DFF_X1 port map( D => n13302, CK => CLK, Q => n5032, 
                           QN => n53386);
   REGS_reg_32_16_inst : DFF_X1 port map( D => n13301, CK => CLK, Q => n5033, 
                           QN => n53387);
   REGS_reg_32_15_inst : DFF_X1 port map( D => n13300, CK => CLK, Q => n5034, 
                           QN => n53388);
   REGS_reg_32_14_inst : DFF_X1 port map( D => n13299, CK => CLK, Q => n5035, 
                           QN => n53389);
   REGS_reg_32_13_inst : DFF_X1 port map( D => n13298, CK => CLK, Q => n5036, 
                           QN => n53390);
   REGS_reg_32_12_inst : DFF_X1 port map( D => n13297, CK => CLK, Q => n5037, 
                           QN => n53391);
   REGS_reg_32_11_inst : DFF_X1 port map( D => n13296, CK => CLK, Q => n5038, 
                           QN => n53392);
   REGS_reg_32_10_inst : DFF_X1 port map( D => n13295, CK => CLK, Q => n5039, 
                           QN => n53393);
   REGS_reg_32_9_inst : DFF_X1 port map( D => n13294, CK => CLK, Q => n5040, QN
                           => n53394);
   REGS_reg_32_8_inst : DFF_X1 port map( D => n13293, CK => CLK, Q => n5041, QN
                           => n53395);
   REGS_reg_32_7_inst : DFF_X1 port map( D => n13292, CK => CLK, Q => n5042, QN
                           => n53396);
   REGS_reg_32_6_inst : DFF_X1 port map( D => n13291, CK => CLK, Q => n5043, QN
                           => n53397);
   REGS_reg_32_5_inst : DFF_X1 port map( D => n13290, CK => CLK, Q => n5044, QN
                           => n53398);
   REGS_reg_32_4_inst : DFF_X1 port map( D => n13289, CK => CLK, Q => n5045, QN
                           => n53399);
   REGS_reg_32_3_inst : DFF_X1 port map( D => n13288, CK => CLK, Q => n5046, QN
                           => n53400);
   REGS_reg_32_2_inst : DFF_X1 port map( D => n13287, CK => CLK, Q => n5047, QN
                           => n53401);
   REGS_reg_32_1_inst : DFF_X1 port map( D => n13286, CK => CLK, Q => n5048, QN
                           => n53402);
   REGS_reg_32_0_inst : DFF_X1 port map( D => n13285, CK => CLK, Q => n5049, QN
                           => n53403);
   REGS_reg_7_23_inst : DFF_X1 port map( D => n14108, CK => CLK, Q => n4432, QN
                           => n53404);
   REGS_reg_7_22_inst : DFF_X1 port map( D => n14107, CK => CLK, Q => n4433, QN
                           => n53405);
   REGS_reg_7_21_inst : DFF_X1 port map( D => n14106, CK => CLK, Q => n4434, QN
                           => n53406);
   REGS_reg_7_20_inst : DFF_X1 port map( D => n14105, CK => CLK, Q => n4435, QN
                           => n53407);
   REGS_reg_7_19_inst : DFF_X1 port map( D => n14104, CK => CLK, Q => n4436, QN
                           => n53408);
   REGS_reg_7_18_inst : DFF_X1 port map( D => n14103, CK => CLK, Q => n4437, QN
                           => n53409);
   REGS_reg_7_17_inst : DFF_X1 port map( D => n14102, CK => CLK, Q => n4438, QN
                           => n53410);
   REGS_reg_7_16_inst : DFF_X1 port map( D => n14101, CK => CLK, Q => n4439, QN
                           => n53411);
   REGS_reg_7_15_inst : DFF_X1 port map( D => n14100, CK => CLK, Q => n4440, QN
                           => n53412);
   REGS_reg_7_14_inst : DFF_X1 port map( D => n14099, CK => CLK, Q => n4441, QN
                           => n53413);
   REGS_reg_7_13_inst : DFF_X1 port map( D => n14098, CK => CLK, Q => n4442, QN
                           => n53414);
   REGS_reg_7_12_inst : DFF_X1 port map( D => n14097, CK => CLK, Q => n4443, QN
                           => n53415);
   REGS_reg_7_11_inst : DFF_X1 port map( D => n14096, CK => CLK, Q => n4444, QN
                           => n53416);
   REGS_reg_7_10_inst : DFF_X1 port map( D => n14095, CK => CLK, Q => n4445, QN
                           => n53417);
   REGS_reg_7_9_inst : DFF_X1 port map( D => n14094, CK => CLK, Q => n4446, QN 
                           => n53418);
   REGS_reg_7_8_inst : DFF_X1 port map( D => n14093, CK => CLK, Q => n4447, QN 
                           => n53419);
   REGS_reg_7_7_inst : DFF_X1 port map( D => n14092, CK => CLK, Q => n4448, QN 
                           => n53420);
   REGS_reg_7_6_inst : DFF_X1 port map( D => n14091, CK => CLK, Q => n4449, QN 
                           => n53421);
   REGS_reg_7_5_inst : DFF_X1 port map( D => n14090, CK => CLK, Q => n4450, QN 
                           => n53422);
   REGS_reg_7_4_inst : DFF_X1 port map( D => n14089, CK => CLK, Q => n4451, QN 
                           => n53423);
   REGS_reg_7_3_inst : DFF_X1 port map( D => n14088, CK => CLK, Q => n4452, QN 
                           => n53424);
   REGS_reg_7_2_inst : DFF_X1 port map( D => n14087, CK => CLK, Q => n4453, QN 
                           => n53425);
   REGS_reg_7_1_inst : DFF_X1 port map( D => n14086, CK => CLK, Q => n4454, QN 
                           => n53426);
   REGS_reg_7_0_inst : DFF_X1 port map( D => n14085, CK => CLK, Q => n4455, QN 
                           => n53427);
   REGS_reg_15_23_inst : DFF_X1 port map( D => n13852, CK => CLK, Q => n4456, 
                           QN => n864);
   REGS_reg_15_22_inst : DFF_X1 port map( D => n13851, CK => CLK, Q => n4457, 
                           QN => n865);
   REGS_reg_15_21_inst : DFF_X1 port map( D => n13850, CK => CLK, Q => n4458, 
                           QN => n866);
   REGS_reg_15_20_inst : DFF_X1 port map( D => n13849, CK => CLK, Q => n4459, 
                           QN => n867);
   REGS_reg_15_19_inst : DFF_X1 port map( D => n13848, CK => CLK, Q => n4460, 
                           QN => n868);
   REGS_reg_15_18_inst : DFF_X1 port map( D => n13847, CK => CLK, Q => n4461, 
                           QN => n869);
   REGS_reg_15_17_inst : DFF_X1 port map( D => n13846, CK => CLK, Q => n4462, 
                           QN => n870);
   REGS_reg_15_16_inst : DFF_X1 port map( D => n13845, CK => CLK, Q => n4463, 
                           QN => n871);
   REGS_reg_15_15_inst : DFF_X1 port map( D => n13844, CK => CLK, Q => n4464, 
                           QN => n872);
   REGS_reg_15_14_inst : DFF_X1 port map( D => n13843, CK => CLK, Q => n4465, 
                           QN => n873);
   REGS_reg_15_13_inst : DFF_X1 port map( D => n13842, CK => CLK, Q => n4466, 
                           QN => n874);
   REGS_reg_15_12_inst : DFF_X1 port map( D => n13841, CK => CLK, Q => n4467, 
                           QN => n875);
   REGS_reg_15_11_inst : DFF_X1 port map( D => n13840, CK => CLK, Q => n4468, 
                           QN => n876);
   REGS_reg_15_10_inst : DFF_X1 port map( D => n13839, CK => CLK, Q => n4469, 
                           QN => n877);
   REGS_reg_15_9_inst : DFF_X1 port map( D => n13838, CK => CLK, Q => n4470, QN
                           => n878);
   REGS_reg_15_8_inst : DFF_X1 port map( D => n13837, CK => CLK, Q => n4471, QN
                           => n879);
   REGS_reg_15_7_inst : DFF_X1 port map( D => n13836, CK => CLK, Q => n4472, QN
                           => n880);
   REGS_reg_15_6_inst : DFF_X1 port map( D => n13835, CK => CLK, Q => n4473, QN
                           => n881);
   REGS_reg_15_5_inst : DFF_X1 port map( D => n13834, CK => CLK, Q => n4474, QN
                           => n882);
   REGS_reg_15_4_inst : DFF_X1 port map( D => n13833, CK => CLK, Q => n4475, QN
                           => n883);
   REGS_reg_15_3_inst : DFF_X1 port map( D => n13832, CK => CLK, Q => n4476, QN
                           => n884);
   REGS_reg_15_2_inst : DFF_X1 port map( D => n13831, CK => CLK, Q => n4477, QN
                           => n885);
   REGS_reg_15_1_inst : DFF_X1 port map( D => n13830, CK => CLK, Q => n4478, QN
                           => n886);
   REGS_reg_15_0_inst : DFF_X1 port map( D => n13829, CK => CLK, Q => n4479, QN
                           => n887);
   REGS_reg_14_23_inst : DFF_X1 port map( D => n13884, CK => CLK, Q => n4480, 
                           QN => n888);
   REGS_reg_14_22_inst : DFF_X1 port map( D => n13883, CK => CLK, Q => n4481, 
                           QN => n889);
   REGS_reg_14_21_inst : DFF_X1 port map( D => n13882, CK => CLK, Q => n4482, 
                           QN => n890);
   REGS_reg_14_20_inst : DFF_X1 port map( D => n13881, CK => CLK, Q => n4483, 
                           QN => n891);
   REGS_reg_14_19_inst : DFF_X1 port map( D => n13880, CK => CLK, Q => n4484, 
                           QN => n892);
   REGS_reg_14_18_inst : DFF_X1 port map( D => n13879, CK => CLK, Q => n4485, 
                           QN => n893);
   REGS_reg_14_17_inst : DFF_X1 port map( D => n13878, CK => CLK, Q => n4486, 
                           QN => n894);
   REGS_reg_14_16_inst : DFF_X1 port map( D => n13877, CK => CLK, Q => n4487, 
                           QN => n895);
   REGS_reg_14_15_inst : DFF_X1 port map( D => n13876, CK => CLK, Q => n4488, 
                           QN => n896);
   REGS_reg_14_14_inst : DFF_X1 port map( D => n13875, CK => CLK, Q => n4489, 
                           QN => n897);
   REGS_reg_14_13_inst : DFF_X1 port map( D => n13874, CK => CLK, Q => n4490, 
                           QN => n898);
   REGS_reg_14_12_inst : DFF_X1 port map( D => n13873, CK => CLK, Q => n4491, 
                           QN => n899);
   REGS_reg_14_11_inst : DFF_X1 port map( D => n13872, CK => CLK, Q => n4492, 
                           QN => n900);
   REGS_reg_14_10_inst : DFF_X1 port map( D => n13871, CK => CLK, Q => n4493, 
                           QN => n901);
   REGS_reg_14_9_inst : DFF_X1 port map( D => n13870, CK => CLK, Q => n4494, QN
                           => n902);
   REGS_reg_14_8_inst : DFF_X1 port map( D => n13869, CK => CLK, Q => n4495, QN
                           => n903);
   REGS_reg_14_7_inst : DFF_X1 port map( D => n13868, CK => CLK, Q => n4496, QN
                           => n904);
   REGS_reg_14_6_inst : DFF_X1 port map( D => n13867, CK => CLK, Q => n4497, QN
                           => n905);
   REGS_reg_14_5_inst : DFF_X1 port map( D => n13866, CK => CLK, Q => n4498, QN
                           => n906);
   REGS_reg_14_4_inst : DFF_X1 port map( D => n13865, CK => CLK, Q => n4499, QN
                           => n907);
   REGS_reg_14_3_inst : DFF_X1 port map( D => n13864, CK => CLK, Q => n4500, QN
                           => n908);
   REGS_reg_14_2_inst : DFF_X1 port map( D => n13863, CK => CLK, Q => n4501, QN
                           => n909);
   REGS_reg_14_1_inst : DFF_X1 port map( D => n13862, CK => CLK, Q => n4502, QN
                           => n910);
   REGS_reg_14_0_inst : DFF_X1 port map( D => n13861, CK => CLK, Q => n4503, QN
                           => n911);
   REGS_reg_11_23_inst : DFF_X1 port map( D => n13980, CK => CLK, Q => n4552, 
                           QN => n912);
   REGS_reg_11_22_inst : DFF_X1 port map( D => n13979, CK => CLK, Q => n4553, 
                           QN => n913);
   REGS_reg_11_21_inst : DFF_X1 port map( D => n13978, CK => CLK, Q => n4554, 
                           QN => n914);
   REGS_reg_11_20_inst : DFF_X1 port map( D => n13977, CK => CLK, Q => n4555, 
                           QN => n915);
   REGS_reg_11_19_inst : DFF_X1 port map( D => n13976, CK => CLK, Q => n4556, 
                           QN => n916);
   REGS_reg_11_18_inst : DFF_X1 port map( D => n13975, CK => CLK, Q => n4557, 
                           QN => n917);
   REGS_reg_11_17_inst : DFF_X1 port map( D => n13974, CK => CLK, Q => n4558, 
                           QN => n918);
   REGS_reg_11_16_inst : DFF_X1 port map( D => n13973, CK => CLK, Q => n4559, 
                           QN => n919);
   REGS_reg_11_15_inst : DFF_X1 port map( D => n13972, CK => CLK, Q => n4560, 
                           QN => n920);
   REGS_reg_11_14_inst : DFF_X1 port map( D => n13971, CK => CLK, Q => n4561, 
                           QN => n921);
   REGS_reg_11_13_inst : DFF_X1 port map( D => n13970, CK => CLK, Q => n4562, 
                           QN => n922);
   REGS_reg_11_12_inst : DFF_X1 port map( D => n13969, CK => CLK, Q => n4563, 
                           QN => n923);
   REGS_reg_11_11_inst : DFF_X1 port map( D => n13968, CK => CLK, Q => n4564, 
                           QN => n924);
   REGS_reg_11_10_inst : DFF_X1 port map( D => n13967, CK => CLK, Q => n4565, 
                           QN => n925);
   REGS_reg_11_9_inst : DFF_X1 port map( D => n13966, CK => CLK, Q => n4566, QN
                           => n926);
   REGS_reg_11_8_inst : DFF_X1 port map( D => n13965, CK => CLK, Q => n4567, QN
                           => n927);
   REGS_reg_11_7_inst : DFF_X1 port map( D => n13964, CK => CLK, Q => n4568, QN
                           => n928);
   REGS_reg_11_6_inst : DFF_X1 port map( D => n13963, CK => CLK, Q => n4569, QN
                           => n929);
   REGS_reg_11_5_inst : DFF_X1 port map( D => n13962, CK => CLK, Q => n4570, QN
                           => n930);
   REGS_reg_11_4_inst : DFF_X1 port map( D => n13961, CK => CLK, Q => n4571, QN
                           => n931);
   REGS_reg_11_3_inst : DFF_X1 port map( D => n13960, CK => CLK, Q => n4572, QN
                           => n932);
   REGS_reg_11_2_inst : DFF_X1 port map( D => n13959, CK => CLK, Q => n4573, QN
                           => n933);
   REGS_reg_11_1_inst : DFF_X1 port map( D => n13958, CK => CLK, Q => n4574, QN
                           => n934);
   REGS_reg_11_0_inst : DFF_X1 port map( D => n13957, CK => CLK, Q => n4575, QN
                           => n935);
   REGS_reg_6_23_inst : DFF_X1 port map( D => n14140, CK => CLK, Q => n4624, QN
                           => n53548);
   REGS_reg_6_22_inst : DFF_X1 port map( D => n14139, CK => CLK, Q => n4625, QN
                           => n53549);
   REGS_reg_6_21_inst : DFF_X1 port map( D => n14138, CK => CLK, Q => n4626, QN
                           => n53550);
   REGS_reg_6_20_inst : DFF_X1 port map( D => n14137, CK => CLK, Q => n4627, QN
                           => n53551);
   REGS_reg_6_19_inst : DFF_X1 port map( D => n14136, CK => CLK, Q => n4628, QN
                           => n53552);
   REGS_reg_6_18_inst : DFF_X1 port map( D => n14135, CK => CLK, Q => n4629, QN
                           => n53553);
   REGS_reg_6_17_inst : DFF_X1 port map( D => n14134, CK => CLK, Q => n4630, QN
                           => n53554);
   REGS_reg_6_16_inst : DFF_X1 port map( D => n14133, CK => CLK, Q => n4631, QN
                           => n53555);
   REGS_reg_6_15_inst : DFF_X1 port map( D => n14132, CK => CLK, Q => n4632, QN
                           => n53556);
   REGS_reg_6_14_inst : DFF_X1 port map( D => n14131, CK => CLK, Q => n4633, QN
                           => n53557);
   REGS_reg_6_13_inst : DFF_X1 port map( D => n14130, CK => CLK, Q => n4634, QN
                           => n53558);
   REGS_reg_6_12_inst : DFF_X1 port map( D => n14129, CK => CLK, Q => n4635, QN
                           => n53559);
   REGS_reg_6_11_inst : DFF_X1 port map( D => n14128, CK => CLK, Q => n4636, QN
                           => n53560);
   REGS_reg_6_10_inst : DFF_X1 port map( D => n14127, CK => CLK, Q => n4637, QN
                           => n53561);
   REGS_reg_6_9_inst : DFF_X1 port map( D => n14126, CK => CLK, Q => n4638, QN 
                           => n53562);
   REGS_reg_6_8_inst : DFF_X1 port map( D => n14125, CK => CLK, Q => n4639, QN 
                           => n53563);
   REGS_reg_6_7_inst : DFF_X1 port map( D => n14124, CK => CLK, Q => n4640, QN 
                           => n53564);
   REGS_reg_6_6_inst : DFF_X1 port map( D => n14123, CK => CLK, Q => n4641, QN 
                           => n53565);
   REGS_reg_6_5_inst : DFF_X1 port map( D => n14122, CK => CLK, Q => n4642, QN 
                           => n53566);
   REGS_reg_6_4_inst : DFF_X1 port map( D => n14121, CK => CLK, Q => n4643, QN 
                           => n53567);
   REGS_reg_6_3_inst : DFF_X1 port map( D => n14120, CK => CLK, Q => n4644, QN 
                           => n53568);
   REGS_reg_6_2_inst : DFF_X1 port map( D => n14119, CK => CLK, Q => n4645, QN 
                           => n53569);
   REGS_reg_6_1_inst : DFF_X1 port map( D => n14118, CK => CLK, Q => n4646, QN 
                           => n53570);
   REGS_reg_6_0_inst : DFF_X1 port map( D => n14117, CK => CLK, Q => n4647, QN 
                           => n53571);
   REGS_reg_3_2_inst : DFF_X1 port map( D => n14215, CK => CLK, Q => n4696, QN 
                           => n53572);
   REGS_reg_3_1_inst : DFF_X1 port map( D => n14214, CK => CLK, Q => n4697, QN 
                           => n53573);
   REGS_reg_3_0_inst : DFF_X1 port map( D => n14213, CK => CLK, Q => n4698, QN 
                           => n53574);
   REGS_reg_2_23_inst : DFF_X1 port map( D => n14268, CK => CLK, Q => n4699, QN
                           => n53575);
   REGS_reg_2_22_inst : DFF_X1 port map( D => n14267, CK => CLK, Q => n4700, QN
                           => n957);
   REGS_reg_2_21_inst : DFF_X1 port map( D => n14266, CK => CLK, Q => n4701, QN
                           => n53576);
   REGS_reg_2_20_inst : DFF_X1 port map( D => n14265, CK => CLK, Q => n4702, QN
                           => n53577);
   REGS_reg_2_19_inst : DFF_X1 port map( D => n14264, CK => CLK, Q => n4703, QN
                           => n53578);
   REGS_reg_2_18_inst : DFF_X1 port map( D => n14263, CK => CLK, Q => n4704, QN
                           => n53579);
   REGS_reg_2_17_inst : DFF_X1 port map( D => n14262, CK => CLK, Q => n4705, QN
                           => n53580);
   REGS_reg_2_16_inst : DFF_X1 port map( D => n14261, CK => CLK, Q => n4706, QN
                           => n53581);
   REGS_reg_2_15_inst : DFF_X1 port map( D => n14260, CK => CLK, Q => n4707, QN
                           => n53582);
   REGS_reg_2_14_inst : DFF_X1 port map( D => n14259, CK => CLK, Q => n4708, QN
                           => n53583);
   REGS_reg_2_13_inst : DFF_X1 port map( D => n14258, CK => CLK, Q => n4709, QN
                           => n958);
   REGS_reg_2_12_inst : DFF_X1 port map( D => n14257, CK => CLK, Q => n4710, QN
                           => n959);
   REGS_reg_2_11_inst : DFF_X1 port map( D => n14256, CK => CLK, Q => n4711, QN
                           => n960);
   REGS_reg_2_10_inst : DFF_X1 port map( D => n14255, CK => CLK, Q => n4712, QN
                           => n961);
   REGS_reg_2_9_inst : DFF_X1 port map( D => n14254, CK => CLK, Q => n4713, QN 
                           => n962);
   REGS_reg_1_23_inst : DFF_X1 port map( D => n14300, CK => CLK, Q => n_2268, 
                           QN => n2213);
   REGS_reg_1_22_inst : DFF_X1 port map( D => n14299, CK => CLK, Q => n_2269, 
                           QN => n2214);
   REGS_reg_1_21_inst : DFF_X1 port map( D => n14298, CK => CLK, Q => n_2270, 
                           QN => n2215);
   REGS_reg_1_20_inst : DFF_X1 port map( D => n14297, CK => CLK, Q => n_2271, 
                           QN => n2216);
   REGS_reg_1_19_inst : DFF_X1 port map( D => n14296, CK => CLK, Q => n_2272, 
                           QN => n2217);
   REGS_reg_1_18_inst : DFF_X1 port map( D => n14295, CK => CLK, Q => n_2273, 
                           QN => n2218);
   REGS_reg_1_17_inst : DFF_X1 port map( D => n14294, CK => CLK, Q => n_2274, 
                           QN => n2219);
   REGS_reg_1_16_inst : DFF_X1 port map( D => n14293, CK => CLK, Q => n_2275, 
                           QN => n2220);
   REGS_reg_1_15_inst : DFF_X1 port map( D => n14292, CK => CLK, Q => n_2276, 
                           QN => n2235);
   REGS_reg_1_14_inst : DFF_X1 port map( D => n14291, CK => CLK, Q => n_2277, 
                           QN => n2236);
   REGS_reg_1_13_inst : DFF_X1 port map( D => n14290, CK => CLK, Q => n_2278, 
                           QN => n2237);
   REGS_reg_1_12_inst : DFF_X1 port map( D => n14289, CK => CLK, Q => n_2279, 
                           QN => n2238);
   REGS_reg_1_11_inst : DFF_X1 port map( D => n14288, CK => CLK, Q => n_2280, 
                           QN => n2075);
   REGS_reg_1_10_inst : DFF_X1 port map( D => n14287, CK => CLK, Q => n_2281, 
                           QN => n2239);
   OUT2_reg_7_inst : DFF_X1 port map( D => n9932, CK => CLK, Q => OUT2(7), QN 
                           => n9339);
   OUT2_reg_6_inst : DFF_X1 port map( D => n9931, CK => CLK, Q => OUT2(6), QN 
                           => n9340);
   OUT2_reg_5_inst : DFF_X1 port map( D => n9930, CK => CLK, Q => OUT2(5), QN 
                           => n9341);
   OUT2_reg_4_inst : DFF_X1 port map( D => n9929, CK => CLK, Q => OUT2(4), QN 
                           => n9342);
   OUT2_reg_3_inst : DFF_X1 port map( D => n9928, CK => CLK, Q => OUT2(3), QN 
                           => n9343);
   OUT2_reg_2_inst : DFF_X1 port map( D => n9927, CK => CLK, Q => OUT2(2), QN 
                           => n9344);
   OUT2_reg_1_inst : DFF_X1 port map( D => n9926, CK => CLK, Q => OUT2(1), QN 
                           => n9345);
   OUT2_reg_0_inst : DFF_X1 port map( D => n9925, CK => CLK, Q => OUT2(0), QN 
                           => n9346);
   OUT2_reg_31_inst : DFF_X1 port map( D => n9956, CK => CLK, Q => OUT2(31), QN
                           => n9315);
   OUT2_reg_30_inst : DFF_X1 port map( D => n9955, CK => CLK, Q => OUT2(30), QN
                           => n9316);
   OUT2_reg_29_inst : DFF_X1 port map( D => n9954, CK => CLK, Q => OUT2(29), QN
                           => n9317);
   OUT2_reg_28_inst : DFF_X1 port map( D => n9953, CK => CLK, Q => OUT2(28), QN
                           => n9318);
   OUT2_reg_27_inst : DFF_X1 port map( D => n9952, CK => CLK, Q => OUT2(27), QN
                           => n9319);
   OUT2_reg_26_inst : DFF_X1 port map( D => n9951, CK => CLK, Q => OUT2(26), QN
                           => n9320);
   OUT2_reg_25_inst : DFF_X1 port map( D => n9950, CK => CLK, Q => OUT2(25), QN
                           => n9321);
   OUT2_reg_24_inst : DFF_X1 port map( D => n9949, CK => CLK, Q => OUT2(24), QN
                           => n9322);
   OUT2_reg_23_inst : DFF_X1 port map( D => n9948, CK => CLK, Q => OUT2(23), QN
                           => n9323);
   OUT2_reg_22_inst : DFF_X1 port map( D => n9947, CK => CLK, Q => OUT2(22), QN
                           => n9324);
   OUT2_reg_21_inst : DFF_X1 port map( D => n9946, CK => CLK, Q => OUT2(21), QN
                           => n9325);
   OUT2_reg_20_inst : DFF_X1 port map( D => n9945, CK => CLK, Q => OUT2(20), QN
                           => n9326);
   OUT2_reg_19_inst : DFF_X1 port map( D => n9944, CK => CLK, Q => OUT2(19), QN
                           => n9327);
   OUT2_reg_18_inst : DFF_X1 port map( D => n9943, CK => CLK, Q => OUT2(18), QN
                           => n9328);
   OUT2_reg_17_inst : DFF_X1 port map( D => n9942, CK => CLK, Q => OUT2(17), QN
                           => n9329);
   OUT2_reg_16_inst : DFF_X1 port map( D => n9941, CK => CLK, Q => OUT2(16), QN
                           => n9330);
   OUT2_reg_15_inst : DFF_X1 port map( D => n9940, CK => CLK, Q => OUT2(15), QN
                           => n9331);
   OUT2_reg_14_inst : DFF_X1 port map( D => n9939, CK => CLK, Q => OUT2(14), QN
                           => n9332);
   OUT2_reg_13_inst : DFF_X1 port map( D => n9938, CK => CLK, Q => OUT2(13), QN
                           => n9333);
   OUT2_reg_12_inst : DFF_X1 port map( D => n9937, CK => CLK, Q => OUT2(12), QN
                           => n9334);
   OUT2_reg_11_inst : DFF_X1 port map( D => n9936, CK => CLK, Q => OUT2(11), QN
                           => n9335);
   OUT2_reg_10_inst : DFF_X1 port map( D => n9935, CK => CLK, Q => OUT2(10), QN
                           => n9336);
   OUT2_reg_9_inst : DFF_X1 port map( D => n9934, CK => CLK, Q => OUT2(9), QN 
                           => n9337);
   OUT2_reg_8_inst : DFF_X1 port map( D => n9933, CK => CLK, Q => OUT2(8), QN 
                           => n9338);
   OUT1_reg_31_inst : DFF_X1 port map( D => n9988, CK => CLK, Q => OUT1(31), QN
                           => n9283);
   OUT1_reg_30_inst : DFF_X1 port map( D => n9987, CK => CLK, Q => OUT1(30), QN
                           => n9284);
   OUT1_reg_29_inst : DFF_X1 port map( D => n9986, CK => CLK, Q => OUT1(29), QN
                           => n9285);
   OUT1_reg_28_inst : DFF_X1 port map( D => n9985, CK => CLK, Q => OUT1(28), QN
                           => n9286);
   OUT1_reg_27_inst : DFF_X1 port map( D => n9984, CK => CLK, Q => OUT1(27), QN
                           => n9287);
   OUT1_reg_26_inst : DFF_X1 port map( D => n9983, CK => CLK, Q => OUT1(26), QN
                           => n9288);
   OUT1_reg_25_inst : DFF_X1 port map( D => n9982, CK => CLK, Q => OUT1(25), QN
                           => n9289);
   OUT1_reg_24_inst : DFF_X1 port map( D => n9981, CK => CLK, Q => OUT1(24), QN
                           => n9290);
   OUT1_reg_23_inst : DFF_X1 port map( D => n9980, CK => CLK, Q => OUT1(23), QN
                           => n9291);
   OUT1_reg_22_inst : DFF_X1 port map( D => n9979, CK => CLK, Q => OUT1(22), QN
                           => n9292);
   OUT1_reg_21_inst : DFF_X1 port map( D => n9978, CK => CLK, Q => OUT1(21), QN
                           => n9293);
   OUT1_reg_20_inst : DFF_X1 port map( D => n9977, CK => CLK, Q => OUT1(20), QN
                           => n9294);
   OUT1_reg_19_inst : DFF_X1 port map( D => n9976, CK => CLK, Q => OUT1(19), QN
                           => n9295);
   OUT1_reg_18_inst : DFF_X1 port map( D => n9975, CK => CLK, Q => OUT1(18), QN
                           => n9296);
   OUT1_reg_17_inst : DFF_X1 port map( D => n9974, CK => CLK, Q => OUT1(17), QN
                           => n9297);
   OUT1_reg_16_inst : DFF_X1 port map( D => n9973, CK => CLK, Q => OUT1(16), QN
                           => n9298);
   OUT1_reg_15_inst : DFF_X1 port map( D => n9972, CK => CLK, Q => OUT1(15), QN
                           => n9299);
   OUT1_reg_14_inst : DFF_X1 port map( D => n9971, CK => CLK, Q => OUT1(14), QN
                           => n9300);
   OUT1_reg_13_inst : DFF_X1 port map( D => n9970, CK => CLK, Q => OUT1(13), QN
                           => n9301);
   OUT1_reg_12_inst : DFF_X1 port map( D => n9969, CK => CLK, Q => OUT1(12), QN
                           => n9302);
   OUT1_reg_11_inst : DFF_X1 port map( D => n9968, CK => CLK, Q => OUT1(11), QN
                           => n9303);
   OUT1_reg_10_inst : DFF_X1 port map( D => n9967, CK => CLK, Q => OUT1(10), QN
                           => n9304);
   OUT1_reg_9_inst : DFF_X1 port map( D => n9966, CK => CLK, Q => OUT1(9), QN 
                           => n9305);
   OUT1_reg_7_inst : DFF_X1 port map( D => n9964, CK => CLK, Q => OUT1(7), QN 
                           => n9307);
   OUT1_reg_8_inst : DFF_X1 port map( D => n9965, CK => CLK, Q => OUT1(8), QN 
                           => n9306);
   OUT1_reg_6_inst : DFF_X1 port map( D => n9963, CK => CLK, Q => OUT1(6), QN 
                           => n9308);
   OUT1_reg_5_inst : DFF_X1 port map( D => n9962, CK => CLK, Q => OUT1(5), QN 
                           => n9309);
   OUT1_reg_4_inst : DFF_X1 port map( D => n9961, CK => CLK, Q => OUT1(4), QN 
                           => n9310);
   OUT1_reg_3_inst : DFF_X1 port map( D => n9960, CK => CLK, Q => OUT1(3), QN 
                           => n9311);
   OUT1_reg_2_inst : DFF_X1 port map( D => n9959, CK => CLK, Q => OUT1(2), QN 
                           => n9312);
   OUT1_reg_1_inst : DFF_X1 port map( D => n9958, CK => CLK, Q => OUT1(1), QN 
                           => n9313);
   U2 : NOR3_X2 port map( A1 => n5360, A2 => n5361, A3 => n5359, ZN => n14983);
   U3 : NOR3_X2 port map( A1 => n5360, A2 => ADDR_RD2(0), A3 => n5359, ZN => 
                           n14984);
   U4 : NOR3_X2 port map( A1 => ADDR_RD2(0), A2 => ADDR_RD2(2), A3 => n5360, ZN
                           => n14979);
   U5 : NOR3_X2 port map( A1 => n5361, A2 => ADDR_RD2(2), A3 => n5360, ZN => 
                           n14978);
   U6 : NOR3_X2 port map( A1 => n5352, A2 => n5353, A3 => n5351, ZN => n7849);
   U7 : AND2_X1 port map( A1 => n7853, A2 => n7850, ZN => n59635);
   U8 : AND2_X1 port map( A1 => n7883, A2 => n7862, ZN => n59636);
   U9 : AND2_X1 port map( A1 => n7883, A2 => n7864, ZN => n59637);
   U10 : AND2_X1 port map( A1 => n7855, A2 => n7864, ZN => n59638);
   U11 : AND2_X1 port map( A1 => n7861, A2 => n7856, ZN => n59639);
   U12 : AND2_X1 port map( A1 => n7857, A2 => n7849, ZN => n59640);
   U13 : AND2_X1 port map( A1 => n7934, A2 => n7849, ZN => n59641);
   U14 : AND2_X1 port map( A1 => n7920, A2 => n7849, ZN => n59642);
   U15 : AND2_X1 port map( A1 => n7920, A2 => n7859, ZN => n59643);
   U16 : AND2_X1 port map( A1 => n7886, A2 => n7852, ZN => n59644);
   U17 : AND2_X1 port map( A1 => n7883, A2 => n7852, ZN => n59645);
   U18 : AND2_X1 port map( A1 => n7853, A2 => n7856, ZN => n59646);
   U19 : AND2_X1 port map( A1 => n7924, A2 => n7852, ZN => n59647);
   U20 : AND2_X1 port map( A1 => n7859, A2 => n7914, ZN => n59648);
   U21 : NAND3_X1 port map( A1 => ADDR_WR(5), A2 => n15126, A3 => ADDR_WR(6), 
                           ZN => n15230);
   U22 : NAND3_X1 port map( A1 => ADDR_WR(5), A2 => n15145, A3 => ADDR_WR(6), 
                           ZN => n15247);
   U23 : NAND3_X1 port map( A1 => n15126, A2 => n5279, A3 => ADDR_WR(6), ZN => 
                           n15188);
   U24 : NAND3_X1 port map( A1 => n15145, A2 => n5279, A3 => ADDR_WR(6), ZN => 
                           n15213);
   U25 : NAND3_X1 port map( A1 => n15126, A2 => n5278, A3 => ADDR_WR(5), ZN => 
                           n15147);
   U26 : NAND3_X1 port map( A1 => n15145, A2 => n5278, A3 => ADDR_WR(5), ZN => 
                           n15164);
   U27 : NAND2_X1 port map( A1 => n15145, A2 => n15127, ZN => n15129);
   U28 : INV_X1 port map( A => n61698, ZN => n61697);
   U29 : INV_X1 port map( A => n59640, ZN => n61733);
   U30 : INV_X1 port map( A => n59641, ZN => n61675);
   U31 : INV_X1 port map( A => n59640, ZN => n61734);
   U32 : INV_X1 port map( A => n59641, ZN => n61676);
   U33 : INV_X1 port map( A => n59642, ZN => n61683);
   U34 : INV_X1 port map( A => n59642, ZN => n61684);
   U35 : BUF_X1 port map( A => n5290, Z => n62179);
   U36 : BUF_X1 port map( A => n5290, Z => n62178);
   U37 : INV_X1 port map( A => n61702, ZN => n61701);
   U38 : INV_X1 port map( A => n61706, ZN => n61705);
   U39 : INV_X1 port map( A => n61724, ZN => n61723);
   U40 : INV_X1 port map( A => n59635, ZN => n61717);
   U41 : INV_X1 port map( A => n61682, ZN => n61681);
   U42 : INV_X1 port map( A => n61690, ZN => n61689);
   U43 : INV_X1 port map( A => n61694, ZN => n61693);
   U44 : INV_X1 port map( A => n61678, ZN => n61677);
   U45 : INV_X1 port map( A => n61710, ZN => n61709);
   U46 : INV_X1 port map( A => n59964, ZN => n59957);
   U47 : INV_X1 port map( A => n59838, ZN => n59831);
   U48 : INV_X1 port map( A => n59829, ZN => n59822);
   U49 : INV_X1 port map( A => n60675, ZN => n60668);
   U50 : INV_X1 port map( A => n60666, ZN => n60659);
   U51 : INV_X1 port map( A => n60657, ZN => n60650);
   U52 : INV_X1 port map( A => n60648, ZN => n60641);
   U53 : INV_X1 port map( A => n60621, ZN => n60614);
   U54 : INV_X1 port map( A => n60612, ZN => n60605);
   U55 : INV_X1 port map( A => n60585, ZN => n60578);
   U56 : INV_X1 port map( A => n60576, ZN => n60569);
   U57 : INV_X1 port map( A => n60549, ZN => n60542);
   U58 : INV_X1 port map( A => n60522, ZN => n60515);
   U59 : INV_X1 port map( A => n60504, ZN => n60497);
   U60 : INV_X1 port map( A => n60495, ZN => n60488);
   U61 : INV_X1 port map( A => n60432, ZN => n60425);
   U62 : INV_X1 port map( A => n60423, ZN => n60416);
   U63 : INV_X1 port map( A => n60927, ZN => n60920);
   U64 : INV_X1 port map( A => n60918, ZN => n60911);
   U65 : INV_X1 port map( A => n60909, ZN => n60902);
   U66 : INV_X1 port map( A => n60891, ZN => n60884);
   U67 : INV_X1 port map( A => n60882, ZN => n60875);
   U68 : INV_X1 port map( A => n60864, ZN => n60857);
   U69 : INV_X1 port map( A => n60855, ZN => n60848);
   U70 : INV_X1 port map( A => n60846, ZN => n60839);
   U71 : INV_X1 port map( A => n60837, ZN => n60830);
   U72 : INV_X1 port map( A => n60828, ZN => n60821);
   U73 : INV_X1 port map( A => n60900, ZN => n60893);
   U74 : INV_X1 port map( A => n60180, ZN => n60173);
   U75 : INV_X1 port map( A => n60819, ZN => n60812);
   U76 : INV_X1 port map( A => n60810, ZN => n60803);
   U77 : INV_X1 port map( A => n60801, ZN => n60794);
   U78 : INV_X1 port map( A => n60720, ZN => n60713);
   U79 : INV_X1 port map( A => n60711, ZN => n60704);
   U80 : INV_X1 port map( A => n60099, ZN => n60092);
   U81 : INV_X1 port map( A => n60090, ZN => n60083);
   U82 : INV_X1 port map( A => n60081, ZN => n60074);
   U83 : INV_X1 port map( A => n60072, ZN => n60065);
   U84 : INV_X1 port map( A => n60063, ZN => n60056);
   U85 : INV_X1 port map( A => n60054, ZN => n60047);
   U86 : INV_X1 port map( A => n60045, ZN => n60038);
   U87 : INV_X1 port map( A => n60036, ZN => n60029);
   U88 : INV_X1 port map( A => n60027, ZN => n60020);
   U89 : INV_X1 port map( A => n60018, ZN => n60011);
   U90 : INV_X1 port map( A => n60009, ZN => n60002);
   U91 : INV_X1 port map( A => n60000, ZN => n59993);
   U92 : INV_X1 port map( A => n59991, ZN => n59984);
   U93 : INV_X1 port map( A => n59982, ZN => n59975);
   U94 : INV_X1 port map( A => n59973, ZN => n59966);
   U95 : INV_X1 port map( A => n59955, ZN => n59948);
   U96 : INV_X1 port map( A => n59946, ZN => n59939);
   U97 : INV_X1 port map( A => n59937, ZN => n59930);
   U98 : INV_X1 port map( A => n59928, ZN => n59921);
   U99 : INV_X1 port map( A => n59919, ZN => n59912);
   U100 : INV_X1 port map( A => n59910, ZN => n59903);
   U101 : INV_X1 port map( A => n59901, ZN => n59894);
   U102 : INV_X1 port map( A => n59892, ZN => n59885);
   U103 : INV_X1 port map( A => n59883, ZN => n59876);
   U104 : INV_X1 port map( A => n59874, ZN => n59867);
   U105 : INV_X1 port map( A => n59865, ZN => n59858);
   U106 : INV_X1 port map( A => n59856, ZN => n59849);
   U107 : INV_X1 port map( A => n59847, ZN => n59840);
   U108 : INV_X1 port map( A => n59820, ZN => n59813);
   U109 : INV_X1 port map( A => n60639, ZN => n60632);
   U110 : INV_X1 port map( A => n60630, ZN => n60623);
   U111 : INV_X1 port map( A => n60603, ZN => n60596);
   U112 : INV_X1 port map( A => n60594, ZN => n60587);
   U113 : INV_X1 port map( A => n60567, ZN => n60560);
   U114 : INV_X1 port map( A => n60558, ZN => n60551);
   U115 : INV_X1 port map( A => n60540, ZN => n60533);
   U116 : INV_X1 port map( A => n60531, ZN => n60524);
   U117 : INV_X1 port map( A => n60513, ZN => n60506);
   U118 : INV_X1 port map( A => n60486, ZN => n60479);
   U119 : INV_X1 port map( A => n60477, ZN => n60470);
   U120 : INV_X1 port map( A => n60468, ZN => n60461);
   U121 : INV_X1 port map( A => n60459, ZN => n60452);
   U122 : INV_X1 port map( A => n60450, ZN => n60443);
   U123 : INV_X1 port map( A => n60441, ZN => n60434);
   U124 : INV_X1 port map( A => n60414, ZN => n60407);
   U125 : INV_X1 port map( A => n60405, ZN => n60398);
   U126 : INV_X1 port map( A => n60396, ZN => n60389);
   U127 : INV_X1 port map( A => n61243, ZN => n61236);
   U128 : INV_X1 port map( A => n60954, ZN => n60947);
   U129 : INV_X1 port map( A => n60945, ZN => n60938);
   U130 : INV_X1 port map( A => n60936, ZN => n60929);
   U131 : INV_X1 port map( A => n60873, ZN => n60866);
   U132 : INV_X1 port map( A => n60387, ZN => n60380);
   U133 : INV_X1 port map( A => n60378, ZN => n60371);
   U134 : INV_X1 port map( A => n60369, ZN => n60362);
   U135 : INV_X1 port map( A => n60360, ZN => n60353);
   U136 : INV_X1 port map( A => n60351, ZN => n60344);
   U137 : INV_X1 port map( A => n60342, ZN => n60335);
   U138 : INV_X1 port map( A => n60333, ZN => n60326);
   U139 : INV_X1 port map( A => n60324, ZN => n60317);
   U140 : INV_X1 port map( A => n60315, ZN => n60308);
   U141 : INV_X1 port map( A => n60306, ZN => n60299);
   U142 : INV_X1 port map( A => n60297, ZN => n60290);
   U143 : INV_X1 port map( A => n60288, ZN => n60281);
   U144 : INV_X1 port map( A => n60279, ZN => n60272);
   U145 : INV_X1 port map( A => n60270, ZN => n60263);
   U146 : INV_X1 port map( A => n60261, ZN => n60254);
   U147 : INV_X1 port map( A => n60252, ZN => n60245);
   U148 : INV_X1 port map( A => n60243, ZN => n60236);
   U149 : INV_X1 port map( A => n60234, ZN => n60227);
   U150 : INV_X1 port map( A => n60225, ZN => n60218);
   U151 : INV_X1 port map( A => n60216, ZN => n60209);
   U152 : INV_X1 port map( A => n60207, ZN => n60200);
   U153 : INV_X1 port map( A => n60198, ZN => n60191);
   U154 : INV_X1 port map( A => n60189, ZN => n60182);
   U155 : INV_X1 port map( A => n60171, ZN => n60164);
   U156 : INV_X1 port map( A => n60162, ZN => n60155);
   U157 : INV_X1 port map( A => n60153, ZN => n60146);
   U158 : INV_X1 port map( A => n60144, ZN => n60137);
   U159 : INV_X1 port map( A => n60135, ZN => n60128);
   U160 : INV_X1 port map( A => n60126, ZN => n60119);
   U161 : INV_X1 port map( A => n60117, ZN => n60110);
   U162 : INV_X1 port map( A => n60108, ZN => n60101);
   U163 : INV_X1 port map( A => n60792, ZN => n60785);
   U164 : INV_X1 port map( A => n60783, ZN => n60776);
   U165 : INV_X1 port map( A => n60774, ZN => n60767);
   U166 : INV_X1 port map( A => n60765, ZN => n60758);
   U167 : INV_X1 port map( A => n60756, ZN => n60749);
   U168 : INV_X1 port map( A => n60747, ZN => n60740);
   U169 : INV_X1 port map( A => n60738, ZN => n60731);
   U170 : INV_X1 port map( A => n60729, ZN => n60722);
   U171 : INV_X1 port map( A => n60702, ZN => n60695);
   U172 : INV_X1 port map( A => n60693, ZN => n60686);
   U173 : INV_X1 port map( A => n60684, ZN => n60677);
   U174 : INV_X1 port map( A => n59645, ZN => n61699);
   U175 : INV_X1 port map( A => n59638, ZN => n61715);
   U176 : INV_X1 port map( A => n59646, ZN => n61725);
   U177 : INV_X1 port map( A => n61722, ZN => n61721);
   U178 : INV_X1 port map( A => n59639, ZN => n61729);
   U179 : INV_X1 port map( A => n59643, ZN => n61687);
   U180 : INV_X1 port map( A => n59645, ZN => n61700);
   U181 : INV_X1 port map( A => n59638, ZN => n61716);
   U182 : INV_X1 port map( A => n59646, ZN => n61726);
   U183 : INV_X1 port map( A => n59639, ZN => n61730);
   U184 : INV_X1 port map( A => n59643, ZN => n61688);
   U185 : INV_X1 port map( A => n61714, ZN => n61713);
   U186 : INV_X1 port map( A => n61720, ZN => n61719);
   U187 : INV_X1 port map( A => n61732, ZN => n61731);
   U188 : INV_X1 port map( A => n61728, ZN => n61727);
   U189 : INV_X1 port map( A => n61686, ZN => n61685);
   U190 : INV_X1 port map( A => n61674, ZN => n61673);
   U191 : INV_X1 port map( A => n59637, ZN => n61703);
   U192 : INV_X1 port map( A => n59636, ZN => n61707);
   U193 : INV_X1 port map( A => n61712, ZN => n61711);
   U194 : INV_X1 port map( A => n59648, ZN => n61691);
   U195 : INV_X1 port map( A => n59644, ZN => n61695);
   U196 : INV_X1 port map( A => n59647, ZN => n61679);
   U197 : INV_X1 port map( A => n59637, ZN => n61704);
   U198 : INV_X1 port map( A => n59636, ZN => n61708);
   U199 : INV_X1 port map( A => n59648, ZN => n61692);
   U200 : INV_X1 port map( A => n59644, ZN => n61696);
   U201 : INV_X1 port map( A => n59647, ZN => n61680);
   U202 : AND2_X1 port map( A1 => n7931, A2 => n7885, ZN => n7896);
   U203 : BUF_X1 port map( A => n5338, Z => n62135);
   U204 : BUF_X1 port map( A => n5338, Z => n62134);
   U205 : BUF_X1 port map( A => n5334, Z => n62139);
   U206 : BUF_X1 port map( A => n5324, Z => n62151);
   U207 : BUF_X1 port map( A => n5334, Z => n62138);
   U208 : BUF_X1 port map( A => n5324, Z => n62150);
   U209 : BUF_X1 port map( A => n5300, Z => n62175);
   U210 : BUF_X1 port map( A => n5300, Z => n62174);
   U211 : BUF_X1 port map( A => n5326, Z => n62147);
   U212 : BUF_X1 port map( A => n5326, Z => n62146);
   U213 : BUF_X1 port map( A => n5321, Z => n62155);
   U214 : BUF_X1 port map( A => n5321, Z => n62154);
   U215 : BUF_X1 port map( A => n5308, Z => n62169);
   U216 : BUF_X1 port map( A => n5308, Z => n62168);
   U217 : BUF_X1 port map( A => n5451, Z => n61873);
   U218 : BUF_X1 port map( A => n5495, Z => n61831);
   U219 : BUF_X1 port map( A => n5451, Z => n61874);
   U220 : BUF_X1 port map( A => n5495, Z => n61832);
   U221 : BUF_X1 port map( A => n5339, Z => n62133);
   U222 : BUF_X1 port map( A => n5339, Z => n62132);
   U223 : BUF_X1 port map( A => n5313, Z => n62165);
   U224 : BUF_X1 port map( A => n5313, Z => n62164);
   U225 : BUF_X1 port map( A => n5322, Z => n62153);
   U226 : BUF_X1 port map( A => n5322, Z => n62152);
   U227 : BUF_X1 port map( A => n5309, Z => n62167);
   U228 : BUF_X1 port map( A => n5335, Z => n62137);
   U229 : BUF_X1 port map( A => n5346, Z => n62127);
   U230 : BUF_X1 port map( A => n5327, Z => n62145);
   U231 : BUF_X1 port map( A => n5309, Z => n62166);
   U232 : BUF_X1 port map( A => n5335, Z => n62136);
   U233 : BUF_X1 port map( A => n5346, Z => n62126);
   U234 : BUF_X1 port map( A => n5327, Z => n62144);
   U235 : BUF_X1 port map( A => n5325, Z => n62149);
   U236 : BUF_X1 port map( A => n5325, Z => n62148);
   U237 : BUF_X1 port map( A => n5414, Z => n61912);
   U238 : BUF_X1 port map( A => n5525, Z => n61789);
   U239 : BUF_X1 port map( A => n5478, Z => n61849);
   U240 : BUF_X1 port map( A => n5548, Z => n61750);
   U241 : BUF_X1 port map( A => n5520, Z => n61801);
   U242 : BUF_X1 port map( A => n5414, Z => n61913);
   U243 : BUF_X1 port map( A => n5525, Z => n61790);
   U244 : BUF_X1 port map( A => n5478, Z => n61850);
   U245 : BUF_X1 port map( A => n5548, Z => n61751);
   U246 : BUF_X1 port map( A => n5520, Z => n61802);
   U247 : INV_X1 port map( A => n59635, ZN => n61718);
   U248 : BUF_X1 port map( A => n5487, Z => n61834);
   U249 : BUF_X1 port map( A => n5487, Z => n61835);
   U250 : BUF_X1 port map( A => n5400, Z => n61937);
   U251 : BUF_X1 port map( A => n5342, Z => n62131);
   U252 : BUF_X1 port map( A => n5342, Z => n62130);
   U253 : BUF_X1 port map( A => n5307, Z => n62171);
   U254 : BUF_X1 port map( A => n5307, Z => n62170);
   U255 : BUF_X1 port map( A => n5316, Z => n62159);
   U256 : BUF_X1 port map( A => n5297, Z => n62177);
   U257 : BUF_X1 port map( A => n5331, Z => n62143);
   U258 : BUF_X1 port map( A => n5316, Z => n62158);
   U259 : BUF_X1 port map( A => n5297, Z => n62176);
   U260 : BUF_X1 port map( A => n5331, Z => n62142);
   U261 : INV_X1 port map( A => n59757, ZN => n59748);
   U262 : BUF_X1 port map( A => n5472, Z => n61861);
   U263 : BUF_X1 port map( A => n8021, Z => n61524);
   U264 : BUF_X1 port map( A => n8021, Z => n61523);
   U265 : BUF_X1 port map( A => n5472, Z => n61862);
   U266 : BUF_X1 port map( A => n5343, Z => n62129);
   U267 : BUF_X1 port map( A => n5343, Z => n62128);
   U268 : BUF_X1 port map( A => n5333, Z => n62140);
   U269 : BUF_X1 port map( A => n5314, Z => n62163);
   U270 : BUF_X1 port map( A => n5314, Z => n62162);
   U271 : BUF_X1 port map( A => n5306, Z => n62173);
   U272 : BUF_X1 port map( A => n5306, Z => n62172);
   U273 : AND2_X1 port map( A1 => n15005, A2 => n15057, ZN => n15068);
   U274 : BUF_X1 port map( A => n5333, Z => n62141);
   U275 : BUF_X1 port map( A => n5284, Z => n62181);
   U276 : BUF_X1 port map( A => n5284, Z => n62180);
   U277 : BUF_X1 port map( A => n5443, Z => n61876);
   U278 : BUF_X1 port map( A => n5400, Z => n61936);
   U279 : BUF_X1 port map( A => n5319, Z => n62157);
   U280 : BUF_X1 port map( A => n5319, Z => n62156);
   U281 : BUF_X1 port map( A => n8062, Z => n61455);
   U282 : BUF_X1 port map( A => n8072, Z => n61431);
   U283 : BUF_X1 port map( A => n8062, Z => n61454);
   U284 : BUF_X1 port map( A => n8072, Z => n61430);
   U285 : BUF_X1 port map( A => n5443, Z => n61877);
   U286 : BUF_X1 port map( A => n8045, Z => n61476);
   U287 : BUF_X1 port map( A => n8134, Z => n61308);
   U288 : BUF_X1 port map( A => n8045, Z => n61475);
   U289 : BUF_X1 port map( A => n8134, Z => n61307);
   U290 : BUF_X1 port map( A => n5451, Z => n61875);
   U291 : BUF_X1 port map( A => n5495, Z => n61833);
   U292 : BUF_X1 port map( A => n5414, Z => n61914);
   U293 : BUF_X1 port map( A => n5520, Z => n61803);
   U294 : BUF_X1 port map( A => n5525, Z => n61791);
   U295 : BUF_X1 port map( A => n5548, Z => n61752);
   U296 : BUF_X1 port map( A => n5478, Z => n61851);
   U297 : BUF_X1 port map( A => n5315, Z => n62161);
   U298 : BUF_X1 port map( A => n5315, Z => n62160);
   U299 : BUF_X1 port map( A => n7974, Z => n61620);
   U300 : BUF_X1 port map( A => n7974, Z => n61619);
   U301 : BUF_X1 port map( A => n8014, Z => n61542);
   U302 : BUF_X1 port map( A => n7989, Z => n61593);
   U303 : BUF_X1 port map( A => n8039, Z => n61491);
   U304 : BUF_X1 port map( A => n7964, Z => n61644);
   U305 : BUF_X1 port map( A => n8113, Z => n61350);
   U306 : BUF_X1 port map( A => n8123, Z => n61326);
   U307 : BUF_X1 port map( A => n8098, Z => n61377);
   U308 : BUF_X1 port map( A => n8088, Z => n61401);
   U309 : BUF_X1 port map( A => n8148, Z => n61275);
   U310 : BUF_X1 port map( A => n8014, Z => n61541);
   U311 : BUF_X1 port map( A => n7989, Z => n61592);
   U312 : BUF_X1 port map( A => n8039, Z => n61490);
   U313 : BUF_X1 port map( A => n7964, Z => n61643);
   U314 : BUF_X1 port map( A => n8113, Z => n61349);
   U315 : BUF_X1 port map( A => n8123, Z => n61325);
   U316 : BUF_X1 port map( A => n8098, Z => n61376);
   U317 : BUF_X1 port map( A => n8088, Z => n61400);
   U318 : BUF_X1 port map( A => n8148, Z => n61274);
   U319 : BUF_X1 port map( A => n8000, Z => n61566);
   U320 : BUF_X1 port map( A => n8000, Z => n61565);
   U321 : BUF_X1 port map( A => n5472, Z => n61863);
   U322 : BUF_X1 port map( A => n8021, Z => n61525);
   U323 : BUF_X1 port map( A => n5487, Z => n61836);
   U324 : BUF_X1 port map( A => n5443, Z => n61878);
   U325 : BUF_X1 port map( A => n8062, Z => n61456);
   U326 : BUF_X1 port map( A => n8072, Z => n61432);
   U327 : BUF_X1 port map( A => n8045, Z => n61477);
   U328 : BUF_X1 port map( A => n8134, Z => n61309);
   U329 : BUF_X1 port map( A => n7974, Z => n61621);
   U330 : BUF_X1 port map( A => n8014, Z => n61543);
   U331 : BUF_X1 port map( A => n7989, Z => n61594);
   U332 : BUF_X1 port map( A => n8039, Z => n61492);
   U333 : BUF_X1 port map( A => n7964, Z => n61645);
   U334 : BUF_X1 port map( A => n8113, Z => n61351);
   U335 : BUF_X1 port map( A => n8123, Z => n61327);
   U336 : BUF_X1 port map( A => n8098, Z => n61378);
   U337 : BUF_X1 port map( A => n8088, Z => n61402);
   U338 : BUF_X1 port map( A => n8148, Z => n61276);
   U339 : BUF_X1 port map( A => n8000, Z => n61567);
   U340 : BUF_X1 port map( A => n5400, Z => n61938);
   U341 : INV_X1 port map( A => n5387, ZN => n5290);
   U342 : INV_X1 port map( A => n59811, ZN => n59804);
   U343 : INV_X1 port map( A => n59802, ZN => n59795);
   U344 : INV_X1 port map( A => n59793, ZN => n59786);
   U345 : INV_X1 port map( A => n59784, ZN => n59777);
   U346 : INV_X1 port map( A => n59775, ZN => n59768);
   U347 : INV_X1 port map( A => n59766, ZN => n59759);
   U348 : INV_X1 port map( A => n62125, ZN => n62118);
   U349 : INV_X1 port map( A => n62125, ZN => n62117);
   U350 : INV_X1 port map( A => n5419, ZN => n5293);
   U351 : INV_X1 port map( A => n5415, ZN => n5289);
   U352 : INV_X1 port map( A => n5416, ZN => n5288);
   U353 : NAND2_X1 port map( A1 => n15284, A2 => n15263, ZN => n15109);
   U354 : NAND2_X1 port map( A1 => n7851, A2 => n7849, ZN => n5387);
   U355 : NAND2_X1 port map( A1 => n15256, A2 => n15263, ZN => n15117);
   U356 : AND2_X1 port map( A1 => n7910, A2 => n7877, ZN => n7914);
   U357 : AND2_X1 port map( A1 => n7889, A2 => n7877, ZN => n7875);
   U358 : AND2_X1 port map( A1 => n7889, A2 => n7885, ZN => n7883);
   U359 : AND2_X1 port map( A1 => n7872, A2 => n7877, ZN => n7853);
   U360 : AND2_X1 port map( A1 => n7873, A2 => n7910, ZN => n7912);
   U361 : AND2_X1 port map( A1 => n7885, A2 => n7910, ZN => n7920);
   U362 : AND2_X1 port map( A1 => n7890, A2 => n7910, ZN => n7886);
   U363 : AND2_X1 port map( A1 => n7889, A2 => n7890, ZN => n7855);
   U364 : AND2_X1 port map( A1 => n15012, A2 => n14993, ZN => n15013);
   U365 : AND2_X1 port map( A1 => n7931, A2 => n7873, ZN => n7848);
   U366 : AND2_X1 port map( A1 => n15036, A2 => n15001, ZN => n15041);
   U367 : AND2_X1 port map( A1 => n15057, A2 => n15001, ZN => n15061);
   U368 : AND2_X1 port map( A1 => n7931, A2 => n7877, ZN => n7934);
   U369 : AND2_X1 port map( A1 => n15012, A2 => n15005, ZN => n15023);
   U370 : BUF_X1 port map( A => n5392, Z => n61949);
   U371 : AND2_X1 port map( A1 => n14993, A2 => n15036, ZN => n15038);
   U372 : BUF_X1 port map( A => n5421, Z => n61906);
   U373 : BUF_X1 port map( A => n5393, Z => n61946);
   U374 : BUF_X1 port map( A => n5526, Z => n61786);
   U375 : BUF_X1 port map( A => n5526, Z => n61787);
   U376 : BUF_X1 port map( A => n5427, Z => n61900);
   U377 : BUF_X1 port map( A => n5432, Z => n61888);
   U378 : BUF_X1 port map( A => n5539, Z => n61771);
   U379 : BUF_X1 port map( A => n5544, Z => n61759);
   U380 : BUF_X1 port map( A => n5511, Z => n61816);
   U381 : BUF_X1 port map( A => n5432, Z => n61889);
   U382 : BUF_X1 port map( A => n5539, Z => n61772);
   U383 : BUF_X1 port map( A => n5544, Z => n61760);
   U384 : BUF_X1 port map( A => n5511, Z => n61817);
   U385 : BUF_X1 port map( A => n5482, Z => n61840);
   U386 : BUF_X1 port map( A => n5482, Z => n61841);
   U387 : BUF_X1 port map( A => n5389, Z => n61954);
   U388 : BUF_X1 port map( A => n5389, Z => n61955);
   U389 : BUF_X1 port map( A => n5438, Z => n61882);
   U390 : BUF_X1 port map( A => n5430, Z => n61894);
   U391 : BUF_X1 port map( A => n5408, Z => n61927);
   U392 : BUF_X1 port map( A => n5413, Z => n61915);
   U393 : BUF_X1 port map( A => n5524, Z => n61792);
   U394 : BUF_X1 port map( A => n5395, Z => n61942);
   U395 : BUF_X1 port map( A => n5477, Z => n61852);
   U396 : BUF_X1 port map( A => n5542, Z => n61765);
   U397 : BUF_X1 port map( A => n5547, Z => n61753);
   U398 : BUF_X1 port map( A => n5514, Z => n61810);
   U399 : BUF_X1 port map( A => n5519, Z => n61804);
   U400 : BUF_X1 port map( A => n5438, Z => n61883);
   U401 : BUF_X1 port map( A => n5430, Z => n61895);
   U402 : BUF_X1 port map( A => n5408, Z => n61928);
   U403 : BUF_X1 port map( A => n5413, Z => n61916);
   U404 : BUF_X1 port map( A => n5524, Z => n61793);
   U405 : BUF_X1 port map( A => n5395, Z => n61943);
   U406 : BUF_X1 port map( A => n5477, Z => n61853);
   U407 : BUF_X1 port map( A => n5542, Z => n61766);
   U408 : BUF_X1 port map( A => n5547, Z => n61754);
   U409 : BUF_X1 port map( A => n5514, Z => n61811);
   U410 : BUF_X1 port map( A => n5519, Z => n61805);
   U411 : BUF_X1 port map( A => n5497, Z => n61825);
   U412 : BUF_X1 port map( A => n5479, Z => n61846);
   U413 : BUF_X1 port map( A => n5474, Z => n61858);
   U414 : BUF_X1 port map( A => n5549, Z => n61747);
   U415 : BUF_X1 port map( A => n5497, Z => n61826);
   U416 : BUF_X1 port map( A => n5479, Z => n61847);
   U417 : BUF_X1 port map( A => n5474, Z => n61859);
   U418 : BUF_X1 port map( A => n5549, Z => n61748);
   U419 : BUF_X1 port map( A => n5553, Z => n61739);
   U420 : BUF_X1 port map( A => n5421, Z => n61907);
   U421 : BUF_X1 port map( A => n5471, Z => n61865);
   U422 : BUF_X1 port map( A => n5427, Z => n61901);
   U423 : BUF_X1 port map( A => n5410, Z => n61922);
   U424 : BUF_X1 port map( A => n5521, Z => n61799);
   U425 : BUF_X1 port map( A => n5439, Z => n61879);
   U426 : BUF_X1 port map( A => n5431, Z => n61891);
   U427 : BUF_X1 port map( A => n5452, Z => n61870);
   U428 : BUF_X1 port map( A => n5409, Z => n61924);
   U429 : BUF_X1 port map( A => n5496, Z => n61828);
   U430 : BUF_X1 port map( A => n5483, Z => n61837);
   U431 : BUF_X1 port map( A => n5543, Z => n61762);
   U432 : BUF_X1 port map( A => n5515, Z => n61807);
   U433 : BUF_X1 port map( A => n5439, Z => n61880);
   U434 : BUF_X1 port map( A => n5431, Z => n61892);
   U435 : BUF_X1 port map( A => n5452, Z => n61871);
   U436 : BUF_X1 port map( A => n5409, Z => n61925);
   U437 : BUF_X1 port map( A => n5496, Z => n61829);
   U438 : BUF_X1 port map( A => n5483, Z => n61838);
   U439 : BUF_X1 port map( A => n5543, Z => n61763);
   U440 : BUF_X1 port map( A => n5515, Z => n61808);
   U441 : AND2_X1 port map( A1 => n15005, A2 => n15036, ZN => n15047);
   U442 : AND2_X1 port map( A1 => n7872, A2 => n7873, ZN => n7857);
   U443 : AND2_X1 port map( A1 => n15057, A2 => n14993, ZN => n15058);
   U444 : AND2_X1 port map( A1 => n7872, A2 => n7885, ZN => n7851);
   U445 : AND2_X1 port map( A1 => n14988, A2 => n15001, ZN => n14992);
   U446 : AND2_X1 port map( A1 => n14988, A2 => n15005, ZN => n15000);
   U447 : AND2_X1 port map( A1 => n14988, A2 => n14993, ZN => n14990);
   U448 : AND2_X1 port map( A1 => n7889, A2 => n7873, ZN => n7870);
   U449 : AND2_X1 port map( A1 => n7931, A2 => n7890, ZN => n7924);
   U450 : BUF_X1 port map( A => n5392, Z => n61948);
   U451 : BUF_X1 port map( A => n5393, Z => n61945);
   U452 : BUF_X1 port map( A => n5553, Z => n61738);
   U453 : BUF_X1 port map( A => n5462, Z => n61867);
   U454 : BUF_X1 port map( A => n5530, Z => n61777);
   U455 : BUF_X1 port map( A => n5462, Z => n61868);
   U456 : BUF_X1 port map( A => n5506, Z => n61819);
   U457 : BUF_X1 port map( A => n5530, Z => n61778);
   U458 : BUF_X1 port map( A => n5411, Z => n61919);
   U459 : BUF_X1 port map( A => n5471, Z => n61864);
   U460 : BUF_X1 port map( A => n5410, Z => n61921);
   U461 : BUF_X1 port map( A => n5521, Z => n61798);
   U462 : BUF_X1 port map( A => n5540, Z => n61769);
   U463 : BUF_X1 port map( A => n5428, Z => n61898);
   U464 : BUF_X1 port map( A => n5554, Z => n61735);
   U465 : BUF_X1 port map( A => n5531, Z => n61774);
   U466 : BUF_X1 port map( A => n5554, Z => n61736);
   U467 : BUF_X1 port map( A => n5531, Z => n61775);
   U468 : BUF_X1 port map( A => n5422, Z => n61904);
   U469 : BUF_X1 port map( A => n5396, Z => n61940);
   U470 : BUF_X1 port map( A => n5506, Z => n61820);
   U471 : BUF_X1 port map( A => n5396, Z => n61939);
   U472 : BUF_X1 port map( A => n5411, Z => n61918);
   U473 : BUF_X1 port map( A => n5418, Z => n61909);
   U474 : BUF_X1 port map( A => n5522, Z => n61795);
   U475 : BUF_X1 port map( A => n5418, Z => n61910);
   U476 : BUF_X1 port map( A => n5522, Z => n61796);
   U477 : BUF_X1 port map( A => n8011, Z => n61548);
   U478 : BUF_X1 port map( A => n8046, Z => n61473);
   U479 : BUF_X1 port map( A => n7956, Z => n61662);
   U480 : BUF_X1 port map( A => n7966, Z => n61638);
   U481 : BUF_X1 port map( A => n8110, Z => n61356);
   U482 : BUF_X1 port map( A => n8120, Z => n61332);
   U483 : BUF_X1 port map( A => n8135, Z => n61305);
   U484 : BUF_X1 port map( A => n8065, Z => n61446);
   U485 : BUF_X1 port map( A => n8011, Z => n61547);
   U486 : BUF_X1 port map( A => n8046, Z => n61472);
   U487 : BUF_X1 port map( A => n7956, Z => n61661);
   U488 : BUF_X1 port map( A => n7966, Z => n61637);
   U489 : BUF_X1 port map( A => n8110, Z => n61355);
   U490 : BUF_X1 port map( A => n8120, Z => n61331);
   U491 : BUF_X1 port map( A => n8135, Z => n61304);
   U492 : BUF_X1 port map( A => n8065, Z => n61445);
   U493 : BUF_X1 port map( A => n8006, Z => n61560);
   U494 : BUF_X1 port map( A => n8016, Z => n61536);
   U495 : BUF_X1 port map( A => n8031, Z => n61509);
   U496 : BUF_X1 port map( A => n8041, Z => n61485);
   U497 : BUF_X1 port map( A => n7961, Z => n61650);
   U498 : BUF_X1 port map( A => n8115, Z => n61344);
   U499 : BUF_X1 port map( A => n8140, Z => n61293);
   U500 : BUF_X1 port map( A => n8150, Z => n61269);
   U501 : BUF_X1 port map( A => n8006, Z => n61559);
   U502 : BUF_X1 port map( A => n8016, Z => n61535);
   U503 : BUF_X1 port map( A => n8031, Z => n61508);
   U504 : BUF_X1 port map( A => n8041, Z => n61484);
   U505 : BUF_X1 port map( A => n7961, Z => n61649);
   U506 : BUF_X1 port map( A => n8115, Z => n61343);
   U507 : BUF_X1 port map( A => n8140, Z => n61292);
   U508 : BUF_X1 port map( A => n8150, Z => n61268);
   U509 : BUF_X1 port map( A => n7996, Z => n61575);
   U510 : BUF_X1 port map( A => n7986, Z => n61599);
   U511 : BUF_X1 port map( A => n7991, Z => n61587);
   U512 : BUF_X1 port map( A => n8036, Z => n61497);
   U513 : BUF_X1 port map( A => n8100, Z => n61371);
   U514 : BUF_X1 port map( A => n8095, Z => n61383);
   U515 : BUF_X1 port map( A => n8145, Z => n61281);
   U516 : BUF_X1 port map( A => n7996, Z => n61574);
   U517 : BUF_X1 port map( A => n7986, Z => n61598);
   U518 : BUF_X1 port map( A => n7991, Z => n61586);
   U519 : BUF_X1 port map( A => n8036, Z => n61496);
   U520 : BUF_X1 port map( A => n8100, Z => n61370);
   U521 : BUF_X1 port map( A => n8095, Z => n61382);
   U522 : BUF_X1 port map( A => n8145, Z => n61280);
   U523 : BUF_X1 port map( A => n8085, Z => n61407);
   U524 : BUF_X1 port map( A => n8085, Z => n61406);
   U525 : BUF_X1 port map( A => n7981, Z => n61611);
   U526 : BUF_X1 port map( A => n8090, Z => n61395);
   U527 : BUF_X1 port map( A => n7981, Z => n61610);
   U528 : BUF_X1 port map( A => n8090, Z => n61394);
   U529 : BUF_X1 port map( A => n5406, Z => n61930);
   U530 : BUF_X1 port map( A => n7971, Z => n61626);
   U531 : BUF_X1 port map( A => n8060, Z => n61458);
   U532 : BUF_X1 port map( A => n7971, Z => n61625);
   U533 : BUF_X1 port map( A => n8060, Z => n61457);
   U534 : BUF_X1 port map( A => n8125, Z => n61320);
   U535 : BUF_X1 port map( A => n8075, Z => n61422);
   U536 : BUF_X1 port map( A => n8070, Z => n61434);
   U537 : BUF_X1 port map( A => n8125, Z => n61319);
   U538 : BUF_X1 port map( A => n8075, Z => n61421);
   U539 : BUF_X1 port map( A => n8070, Z => n61433);
   U540 : BUF_X1 port map( A => n5406, Z => n61931);
   U541 : BUF_X1 port map( A => n5552, Z => n61741);
   U542 : BUF_X1 port map( A => n5529, Z => n61780);
   U543 : BUF_X1 port map( A => n5529, Z => n61781);
   U544 : AND2_X1 port map( A1 => n14987, A2 => n15036, ZN => n15026);
   U545 : BUF_X1 port map( A => n5422, Z => n61903);
   U546 : BUF_X1 port map( A => n5552, Z => n61742);
   U547 : BUF_X1 port map( A => n8077, Z => n61419);
   U548 : BUF_X1 port map( A => n8077, Z => n61418);
   U549 : BUF_X1 port map( A => n8023, Z => n61521);
   U550 : BUF_X1 port map( A => n7998, Z => n61572);
   U551 : BUF_X1 port map( A => n8048, Z => n61470);
   U552 : BUF_X1 port map( A => n7973, Z => n61623);
   U553 : BUF_X1 port map( A => n8127, Z => n61317);
   U554 : BUF_X1 port map( A => n8102, Z => n61368);
   U555 : BUF_X1 port map( A => n8152, Z => n61266);
   U556 : BUF_X1 port map( A => n8023, Z => n61520);
   U557 : BUF_X1 port map( A => n7998, Z => n61571);
   U558 : BUF_X1 port map( A => n8048, Z => n61469);
   U559 : BUF_X1 port map( A => n7973, Z => n61622);
   U560 : BUF_X1 port map( A => n8127, Z => n61316);
   U561 : BUF_X1 port map( A => n8102, Z => n61367);
   U562 : BUF_X1 port map( A => n8152, Z => n61265);
   U563 : BUF_X1 port map( A => n5540, Z => n61768);
   U564 : BUF_X1 port map( A => n5428, Z => n61897);
   U565 : BUF_X1 port map( A => n8008, Z => n61557);
   U566 : BUF_X1 port map( A => n8013, Z => n61545);
   U567 : BUF_X1 port map( A => n8018, Z => n61533);
   U568 : BUF_X1 port map( A => n7983, Z => n61608);
   U569 : BUF_X1 port map( A => n7988, Z => n61596);
   U570 : BUF_X1 port map( A => n7993, Z => n61584);
   U571 : BUF_X1 port map( A => n8033, Z => n61506);
   U572 : BUF_X1 port map( A => n8038, Z => n61494);
   U573 : BUF_X1 port map( A => n8043, Z => n61482);
   U574 : BUF_X1 port map( A => n7958, Z => n61659);
   U575 : BUF_X1 port map( A => n7963, Z => n61647);
   U576 : BUF_X1 port map( A => n7968, Z => n61635);
   U577 : BUF_X1 port map( A => n8112, Z => n61353);
   U578 : BUF_X1 port map( A => n8117, Z => n61341);
   U579 : BUF_X1 port map( A => n8122, Z => n61329);
   U580 : BUF_X1 port map( A => n8097, Z => n61380);
   U581 : BUF_X1 port map( A => n8087, Z => n61404);
   U582 : BUF_X1 port map( A => n8092, Z => n61392);
   U583 : BUF_X1 port map( A => n8137, Z => n61302);
   U584 : BUF_X1 port map( A => n8142, Z => n61290);
   U585 : BUF_X1 port map( A => n8147, Z => n61278);
   U586 : BUF_X1 port map( A => n8067, Z => n61443);
   U587 : BUF_X1 port map( A => n8008, Z => n61556);
   U588 : BUF_X1 port map( A => n8013, Z => n61544);
   U589 : BUF_X1 port map( A => n8018, Z => n61532);
   U590 : BUF_X1 port map( A => n7983, Z => n61607);
   U591 : BUF_X1 port map( A => n7988, Z => n61595);
   U592 : BUF_X1 port map( A => n7993, Z => n61583);
   U593 : BUF_X1 port map( A => n8033, Z => n61505);
   U594 : BUF_X1 port map( A => n8038, Z => n61493);
   U595 : BUF_X1 port map( A => n8043, Z => n61481);
   U596 : BUF_X1 port map( A => n7958, Z => n61658);
   U597 : BUF_X1 port map( A => n7963, Z => n61646);
   U598 : BUF_X1 port map( A => n7968, Z => n61634);
   U599 : BUF_X1 port map( A => n8112, Z => n61352);
   U600 : BUF_X1 port map( A => n8117, Z => n61340);
   U601 : BUF_X1 port map( A => n8122, Z => n61328);
   U602 : BUF_X1 port map( A => n8097, Z => n61379);
   U603 : BUF_X1 port map( A => n8087, Z => n61403);
   U604 : BUF_X1 port map( A => n8092, Z => n61391);
   U605 : BUF_X1 port map( A => n8137, Z => n61301);
   U606 : BUF_X1 port map( A => n8142, Z => n61289);
   U607 : BUF_X1 port map( A => n8147, Z => n61277);
   U608 : BUF_X1 port map( A => n8067, Z => n61442);
   U609 : BUF_X1 port map( A => n5405, Z => n61933);
   U610 : BUF_X1 port map( A => n5405, Z => n61934);
   U611 : BUF_X1 port map( A => n7970, Z => n61629);
   U612 : BUF_X1 port map( A => n8059, Z => n61461);
   U613 : BUF_X1 port map( A => n8069, Z => n61437);
   U614 : BUF_X1 port map( A => n7970, Z => n61628);
   U615 : BUF_X1 port map( A => n8059, Z => n61460);
   U616 : BUF_X1 port map( A => n8069, Z => n61436);
   U617 : BUF_X1 port map( A => n8020, Z => n61527);
   U618 : BUF_X1 port map( A => n7980, Z => n61614);
   U619 : BUF_X1 port map( A => n8124, Z => n61323);
   U620 : BUF_X1 port map( A => n8089, Z => n61398);
   U621 : BUF_X1 port map( A => n8020, Z => n61526);
   U622 : BUF_X1 port map( A => n7980, Z => n61613);
   U623 : BUF_X1 port map( A => n8124, Z => n61322);
   U624 : BUF_X1 port map( A => n8089, Z => n61397);
   U625 : BUF_X1 port map( A => n8074, Z => n61425);
   U626 : BUF_X1 port map( A => n8074, Z => n61424);
   U627 : BUF_X1 port map( A => n8010, Z => n61551);
   U628 : BUF_X1 port map( A => n7990, Z => n61590);
   U629 : BUF_X1 port map( A => n8035, Z => n61500);
   U630 : BUF_X1 port map( A => n7955, Z => n61665);
   U631 : BUF_X1 port map( A => n7965, Z => n61641);
   U632 : BUF_X1 port map( A => n8109, Z => n61359);
   U633 : BUF_X1 port map( A => n8119, Z => n61335);
   U634 : BUF_X1 port map( A => n8099, Z => n61374);
   U635 : BUF_X1 port map( A => n8144, Z => n61284);
   U636 : BUF_X1 port map( A => n8064, Z => n61449);
   U637 : BUF_X1 port map( A => n8010, Z => n61550);
   U638 : BUF_X1 port map( A => n7990, Z => n61589);
   U639 : BUF_X1 port map( A => n8035, Z => n61499);
   U640 : BUF_X1 port map( A => n7955, Z => n61664);
   U641 : BUF_X1 port map( A => n7965, Z => n61640);
   U642 : BUF_X1 port map( A => n8109, Z => n61358);
   U643 : BUF_X1 port map( A => n8119, Z => n61334);
   U644 : BUF_X1 port map( A => n8099, Z => n61373);
   U645 : BUF_X1 port map( A => n8144, Z => n61283);
   U646 : BUF_X1 port map( A => n8064, Z => n61448);
   U647 : BUF_X1 port map( A => n8005, Z => n61563);
   U648 : BUF_X1 port map( A => n8015, Z => n61539);
   U649 : BUF_X1 port map( A => n7995, Z => n61578);
   U650 : BUF_X1 port map( A => n7985, Z => n61602);
   U651 : BUF_X1 port map( A => n7960, Z => n61653);
   U652 : BUF_X1 port map( A => n8114, Z => n61347);
   U653 : BUF_X1 port map( A => n8094, Z => n61386);
   U654 : BUF_X1 port map( A => n8005, Z => n61562);
   U655 : BUF_X1 port map( A => n8015, Z => n61538);
   U656 : BUF_X1 port map( A => n7995, Z => n61577);
   U657 : BUF_X1 port map( A => n7985, Z => n61601);
   U658 : BUF_X1 port map( A => n7960, Z => n61652);
   U659 : BUF_X1 port map( A => n8114, Z => n61346);
   U660 : BUF_X1 port map( A => n8094, Z => n61385);
   U661 : BUF_X1 port map( A => n5526, Z => n61788);
   U662 : BUF_X1 port map( A => n8030, Z => n61512);
   U663 : BUF_X1 port map( A => n8040, Z => n61488);
   U664 : BUF_X1 port map( A => n8084, Z => n61410);
   U665 : BUF_X1 port map( A => n8139, Z => n61296);
   U666 : BUF_X1 port map( A => n8149, Z => n61272);
   U667 : BUF_X1 port map( A => n8030, Z => n61511);
   U668 : BUF_X1 port map( A => n8040, Z => n61487);
   U669 : BUF_X1 port map( A => n8084, Z => n61409);
   U670 : BUF_X1 port map( A => n8139, Z => n61295);
   U671 : BUF_X1 port map( A => n8149, Z => n61271);
   U672 : BUF_X1 port map( A => n5432, Z => n61890);
   U673 : BUF_X1 port map( A => n5511, Z => n61818);
   U674 : BUF_X1 port map( A => n5544, Z => n61761);
   U675 : BUF_X1 port map( A => n5482, Z => n61842);
   U676 : BUF_X1 port map( A => n5389, Z => n61956);
   U677 : BUF_X1 port map( A => n5549, Z => n61749);
   U678 : BUF_X1 port map( A => n5408, Z => n61929);
   U679 : BUF_X1 port map( A => n5413, Z => n61917);
   U680 : BUF_X1 port map( A => n5438, Z => n61884);
   U681 : BUF_X1 port map( A => n5430, Z => n61896);
   U682 : BUF_X1 port map( A => n5395, Z => n61944);
   U683 : BUF_X1 port map( A => n5514, Z => n61812);
   U684 : BUF_X1 port map( A => n5519, Z => n61806);
   U685 : BUF_X1 port map( A => n5524, Z => n61794);
   U686 : BUF_X1 port map( A => n5542, Z => n61767);
   U687 : BUF_X1 port map( A => n5547, Z => n61755);
   U688 : BUF_X1 port map( A => n5477, Z => n61854);
   U689 : BUF_X1 port map( A => n5497, Z => n61827);
   U690 : BUF_X1 port map( A => n5474, Z => n61860);
   U691 : BUF_X1 port map( A => n5479, Z => n61848);
   U692 : BUF_X1 port map( A => n5409, Z => n61926);
   U693 : BUF_X1 port map( A => n5452, Z => n61872);
   U694 : BUF_X1 port map( A => n5439, Z => n61881);
   U695 : BUF_X1 port map( A => n5431, Z => n61893);
   U696 : BUF_X1 port map( A => n5515, Z => n61809);
   U697 : BUF_X1 port map( A => n5543, Z => n61764);
   U698 : BUF_X1 port map( A => n5496, Z => n61830);
   U699 : BUF_X1 port map( A => n5483, Z => n61839);
   U700 : NOR2_X1 port map( A1 => n5350, A2 => n5349, ZN => n7885);
   U701 : NOR2_X1 port map( A1 => n5358, A2 => n5357, ZN => n15005);
   U702 : NOR2_X1 port map( A1 => n5356, A2 => n5355, ZN => n15057);
   U703 : BUF_X1 port map( A => n8024, Z => n61518);
   U704 : BUF_X1 port map( A => n7999, Z => n61569);
   U705 : BUF_X1 port map( A => n8049, Z => n61467);
   U706 : BUF_X1 port map( A => n8128, Z => n61314);
   U707 : BUF_X1 port map( A => n8103, Z => n61365);
   U708 : BUF_X1 port map( A => n8153, Z => n61263);
   U709 : BUF_X1 port map( A => n8078, Z => n61416);
   U710 : BUF_X1 port map( A => n8024, Z => n61517);
   U711 : BUF_X1 port map( A => n7999, Z => n61568);
   U712 : BUF_X1 port map( A => n8049, Z => n61466);
   U713 : BUF_X1 port map( A => n8128, Z => n61313);
   U714 : BUF_X1 port map( A => n8103, Z => n61364);
   U715 : BUF_X1 port map( A => n8153, Z => n61262);
   U716 : BUF_X1 port map( A => n8078, Z => n61415);
   U717 : NOR2_X1 port map( A1 => n5348, A2 => n5347, ZN => n7931);
   U718 : BUF_X1 port map( A => n5433, Z => n61885);
   U719 : BUF_X1 port map( A => n5475, Z => n61855);
   U720 : BUF_X1 port map( A => n5512, Z => n61813);
   U721 : BUF_X1 port map( A => n5433, Z => n61886);
   U722 : BUF_X1 port map( A => n5475, Z => n61856);
   U723 : BUF_X1 port map( A => n5512, Z => n61814);
   U724 : BUF_X1 port map( A => n5390, Z => n61951);
   U725 : BUF_X1 port map( A => n5550, Z => n61744);
   U726 : BUF_X1 port map( A => n5390, Z => n61952);
   U727 : BUF_X1 port map( A => n5550, Z => n61745);
   U728 : BUF_X1 port map( A => n5545, Z => n61756);
   U729 : BUF_X1 port map( A => n5545, Z => n61757);
   U730 : BUF_X1 port map( A => n5480, Z => n61843);
   U731 : BUF_X1 port map( A => n5480, Z => n61844);
   U732 : BUF_X1 port map( A => n5498, Z => n61822);
   U733 : BUF_X1 port map( A => n5498, Z => n61823);
   U734 : BUF_X1 port map( A => n5527, Z => n61783);
   U735 : BUF_X1 port map( A => n5527, Z => n61784);
   U736 : BUF_X1 port map( A => n8009, Z => n61554);
   U737 : BUF_X1 port map( A => n8019, Z => n61530);
   U738 : BUF_X1 port map( A => n7984, Z => n61605);
   U739 : BUF_X1 port map( A => n7994, Z => n61581);
   U740 : BUF_X1 port map( A => n8034, Z => n61503);
   U741 : BUF_X1 port map( A => n8044, Z => n61479);
   U742 : BUF_X1 port map( A => n7959, Z => n61656);
   U743 : BUF_X1 port map( A => n7969, Z => n61632);
   U744 : BUF_X1 port map( A => n8118, Z => n61338);
   U745 : BUF_X1 port map( A => n8093, Z => n61389);
   U746 : BUF_X1 port map( A => n8138, Z => n61299);
   U747 : BUF_X1 port map( A => n8143, Z => n61287);
   U748 : BUF_X1 port map( A => n8063, Z => n61452);
   U749 : BUF_X1 port map( A => n8068, Z => n61440);
   U750 : BUF_X1 port map( A => n8073, Z => n61428);
   U751 : BUF_X1 port map( A => n8009, Z => n61553);
   U752 : BUF_X1 port map( A => n8019, Z => n61529);
   U753 : BUF_X1 port map( A => n7984, Z => n61604);
   U754 : BUF_X1 port map( A => n7994, Z => n61580);
   U755 : BUF_X1 port map( A => n8034, Z => n61502);
   U756 : BUF_X1 port map( A => n8044, Z => n61478);
   U757 : BUF_X1 port map( A => n7959, Z => n61655);
   U758 : BUF_X1 port map( A => n7969, Z => n61631);
   U759 : BUF_X1 port map( A => n8118, Z => n61337);
   U760 : BUF_X1 port map( A => n8093, Z => n61388);
   U761 : BUF_X1 port map( A => n8138, Z => n61298);
   U762 : BUF_X1 port map( A => n8143, Z => n61286);
   U763 : BUF_X1 port map( A => n8063, Z => n61451);
   U764 : BUF_X1 port map( A => n8068, Z => n61439);
   U765 : BUF_X1 port map( A => n8073, Z => n61427);
   U766 : AND2_X1 port map( A1 => n15057, A2 => n14987, ZN => n15050);
   U767 : AND2_X1 port map( A1 => n15012, A2 => n14987, ZN => n15004);
   U768 : AND2_X1 port map( A1 => n15012, A2 => n15001, ZN => n15016);
   U769 : BUF_X1 port map( A => n5531, Z => n61776);
   U770 : BUF_X1 port map( A => n5539, Z => n61773);
   U771 : BUF_X1 port map( A => n8025, Z => n61515);
   U772 : BUF_X1 port map( A => n8050, Z => n61464);
   U773 : BUF_X1 port map( A => n7975, Z => n61617);
   U774 : BUF_X1 port map( A => n8129, Z => n61311);
   U775 : BUF_X1 port map( A => n8104, Z => n61362);
   U776 : BUF_X1 port map( A => n8154, Z => n61260);
   U777 : BUF_X1 port map( A => n8079, Z => n61413);
   U778 : BUF_X1 port map( A => n8025, Z => n61514);
   U779 : BUF_X1 port map( A => n8050, Z => n61463);
   U780 : BUF_X1 port map( A => n7975, Z => n61616);
   U781 : BUF_X1 port map( A => n8129, Z => n61310);
   U782 : BUF_X1 port map( A => n8104, Z => n61361);
   U783 : BUF_X1 port map( A => n8154, Z => n61259);
   U784 : BUF_X1 port map( A => n8079, Z => n61412);
   U785 : BUF_X1 port map( A => n8011, Z => n61549);
   U786 : BUF_X1 port map( A => n8046, Z => n61474);
   U787 : BUF_X1 port map( A => n7956, Z => n61663);
   U788 : BUF_X1 port map( A => n7966, Z => n61639);
   U789 : BUF_X1 port map( A => n8110, Z => n61357);
   U790 : BUF_X1 port map( A => n8120, Z => n61333);
   U791 : BUF_X1 port map( A => n8135, Z => n61306);
   U792 : BUF_X1 port map( A => n8065, Z => n61447);
   U793 : BUF_X1 port map( A => n8006, Z => n61561);
   U794 : BUF_X1 port map( A => n8016, Z => n61537);
   U795 : BUF_X1 port map( A => n8031, Z => n61510);
   U796 : BUF_X1 port map( A => n8041, Z => n61486);
   U797 : BUF_X1 port map( A => n7961, Z => n61651);
   U798 : BUF_X1 port map( A => n8115, Z => n61345);
   U799 : BUF_X1 port map( A => n8140, Z => n61294);
   U800 : BUF_X1 port map( A => n8150, Z => n61270);
   U801 : BUF_X1 port map( A => n7996, Z => n61576);
   U802 : BUF_X1 port map( A => n7986, Z => n61600);
   U803 : BUF_X1 port map( A => n7991, Z => n61588);
   U804 : BUF_X1 port map( A => n8036, Z => n61498);
   U805 : BUF_X1 port map( A => n8100, Z => n61372);
   U806 : BUF_X1 port map( A => n8095, Z => n61384);
   U807 : BUF_X1 port map( A => n8145, Z => n61282);
   U808 : BUF_X1 port map( A => n8085, Z => n61408);
   U809 : BUF_X1 port map( A => n7981, Z => n61612);
   U810 : BUF_X1 port map( A => n8090, Z => n61396);
   U811 : BUF_X1 port map( A => n5406, Z => n61932);
   U812 : BUF_X1 port map( A => n7971, Z => n61627);
   U813 : BUF_X1 port map( A => n8060, Z => n61459);
   U814 : BUF_X1 port map( A => n8125, Z => n61321);
   U815 : BUF_X1 port map( A => n8075, Z => n61423);
   U816 : BUF_X1 port map( A => n8070, Z => n61435);
   U817 : BUF_X1 port map( A => n5462, Z => n61869);
   U818 : BUF_X1 port map( A => n8077, Z => n61420);
   U819 : BUF_X1 port map( A => n5529, Z => n61782);
   U820 : BUF_X1 port map( A => n5552, Z => n61743);
   U821 : BUF_X1 port map( A => n8023, Z => n61522);
   U822 : BUF_X1 port map( A => n7998, Z => n61573);
   U823 : BUF_X1 port map( A => n8048, Z => n61471);
   U824 : BUF_X1 port map( A => n7973, Z => n61624);
   U825 : BUF_X1 port map( A => n8127, Z => n61318);
   U826 : BUF_X1 port map( A => n8102, Z => n61369);
   U827 : BUF_X1 port map( A => n8152, Z => n61267);
   U828 : BUF_X1 port map( A => n8008, Z => n61558);
   U829 : BUF_X1 port map( A => n8013, Z => n61546);
   U830 : BUF_X1 port map( A => n8018, Z => n61534);
   U831 : BUF_X1 port map( A => n7983, Z => n61609);
   U832 : BUF_X1 port map( A => n7988, Z => n61597);
   U833 : BUF_X1 port map( A => n7993, Z => n61585);
   U834 : BUF_X1 port map( A => n8033, Z => n61507);
   U835 : BUF_X1 port map( A => n8038, Z => n61495);
   U836 : BUF_X1 port map( A => n8043, Z => n61483);
   U837 : BUF_X1 port map( A => n7958, Z => n61660);
   U838 : BUF_X1 port map( A => n7963, Z => n61648);
   U839 : BUF_X1 port map( A => n7968, Z => n61636);
   U840 : BUF_X1 port map( A => n8112, Z => n61354);
   U841 : BUF_X1 port map( A => n8117, Z => n61342);
   U842 : BUF_X1 port map( A => n8122, Z => n61330);
   U843 : BUF_X1 port map( A => n8097, Z => n61381);
   U844 : BUF_X1 port map( A => n8087, Z => n61405);
   U845 : BUF_X1 port map( A => n8092, Z => n61393);
   U846 : BUF_X1 port map( A => n8137, Z => n61303);
   U847 : BUF_X1 port map( A => n8142, Z => n61291);
   U848 : BUF_X1 port map( A => n8147, Z => n61279);
   U849 : BUF_X1 port map( A => n8067, Z => n61444);
   U850 : BUF_X1 port map( A => n5418, Z => n61911);
   U851 : BUF_X1 port map( A => n5405, Z => n61935);
   U852 : BUF_X1 port map( A => n7970, Z => n61630);
   U853 : BUF_X1 port map( A => n8059, Z => n61462);
   U854 : BUF_X1 port map( A => n8069, Z => n61438);
   U855 : BUF_X1 port map( A => n8020, Z => n61528);
   U856 : BUF_X1 port map( A => n7980, Z => n61615);
   U857 : BUF_X1 port map( A => n8124, Z => n61324);
   U858 : BUF_X1 port map( A => n8089, Z => n61399);
   U859 : BUF_X1 port map( A => n8074, Z => n61426);
   U860 : BUF_X1 port map( A => n8010, Z => n61552);
   U861 : BUF_X1 port map( A => n7990, Z => n61591);
   U862 : BUF_X1 port map( A => n8035, Z => n61501);
   U863 : BUF_X1 port map( A => n7955, Z => n61666);
   U864 : BUF_X1 port map( A => n7965, Z => n61642);
   U865 : BUF_X1 port map( A => n8109, Z => n61360);
   U866 : BUF_X1 port map( A => n8119, Z => n61336);
   U867 : BUF_X1 port map( A => n8099, Z => n61375);
   U868 : BUF_X1 port map( A => n8144, Z => n61285);
   U869 : BUF_X1 port map( A => n8064, Z => n61450);
   U870 : BUF_X1 port map( A => n8005, Z => n61564);
   U871 : BUF_X1 port map( A => n8015, Z => n61540);
   U872 : BUF_X1 port map( A => n7995, Z => n61579);
   U873 : BUF_X1 port map( A => n7985, Z => n61603);
   U874 : BUF_X1 port map( A => n7960, Z => n61654);
   U875 : BUF_X1 port map( A => n8114, Z => n61348);
   U876 : BUF_X1 port map( A => n8094, Z => n61387);
   U877 : BUF_X1 port map( A => n8030, Z => n61513);
   U878 : BUF_X1 port map( A => n8040, Z => n61489);
   U879 : BUF_X1 port map( A => n8084, Z => n61411);
   U880 : BUF_X1 port map( A => n8139, Z => n61297);
   U881 : BUF_X1 port map( A => n8149, Z => n61273);
   U882 : BUF_X1 port map( A => n5554, Z => n61737);
   U883 : BUF_X1 port map( A => n5530, Z => n61779);
   U884 : BUF_X1 port map( A => n5506, Z => n61821);
   U885 : BUF_X1 port map( A => n8024, Z => n61519);
   U886 : BUF_X1 port map( A => n7999, Z => n61570);
   U887 : BUF_X1 port map( A => n8049, Z => n61468);
   U888 : BUF_X1 port map( A => n8128, Z => n61315);
   U889 : BUF_X1 port map( A => n8103, Z => n61366);
   U890 : BUF_X1 port map( A => n8153, Z => n61264);
   U891 : BUF_X1 port map( A => n8078, Z => n61417);
   U892 : BUF_X1 port map( A => n5433, Z => n61887);
   U893 : BUF_X1 port map( A => n5512, Z => n61815);
   U894 : BUF_X1 port map( A => n5475, Z => n61857);
   U895 : BUF_X1 port map( A => n5390, Z => n61953);
   U896 : BUF_X1 port map( A => n5522, Z => n61797);
   U897 : BUF_X1 port map( A => n5550, Z => n61746);
   U898 : BUF_X1 port map( A => n5545, Z => n61758);
   U899 : BUF_X1 port map( A => n5480, Z => n61845);
   U900 : BUF_X1 port map( A => n5498, Z => n61824);
   U901 : BUF_X1 port map( A => n5527, Z => n61785);
   U902 : BUF_X1 port map( A => n8009, Z => n61555);
   U903 : BUF_X1 port map( A => n8019, Z => n61531);
   U904 : BUF_X1 port map( A => n7984, Z => n61606);
   U905 : BUF_X1 port map( A => n7994, Z => n61582);
   U906 : BUF_X1 port map( A => n8034, Z => n61504);
   U907 : BUF_X1 port map( A => n8044, Z => n61480);
   U908 : BUF_X1 port map( A => n7959, Z => n61657);
   U909 : BUF_X1 port map( A => n7969, Z => n61633);
   U910 : BUF_X1 port map( A => n8118, Z => n61339);
   U911 : BUF_X1 port map( A => n8093, Z => n61390);
   U912 : BUF_X1 port map( A => n8138, Z => n61300);
   U913 : BUF_X1 port map( A => n8143, Z => n61288);
   U914 : BUF_X1 port map( A => n8063, Z => n61453);
   U915 : BUF_X1 port map( A => n8068, Z => n61441);
   U916 : BUF_X1 port map( A => n8073, Z => n61429);
   U917 : BUF_X1 port map( A => n8025, Z => n61516);
   U918 : BUF_X1 port map( A => n8050, Z => n61465);
   U919 : BUF_X1 port map( A => n7975, Z => n61618);
   U920 : BUF_X1 port map( A => n8129, Z => n61312);
   U921 : BUF_X1 port map( A => n8104, Z => n61363);
   U922 : BUF_X1 port map( A => n8154, Z => n61261);
   U923 : BUF_X1 port map( A => n8079, Z => n61414);
   U924 : NAND2_X1 port map( A1 => n7875, A2 => n7849, ZN => n6062);
   U925 : NAND2_X1 port map( A1 => n7883, A2 => n7849, ZN => n5472);
   U926 : BUF_X1 port map( A => n5471, Z => n61866);
   U927 : BUF_X1 port map( A => n5427, Z => n61902);
   U928 : BUF_X1 port map( A => n5392, Z => n61950);
   U929 : BUF_X1 port map( A => n5410, Z => n61923);
   U930 : BUF_X1 port map( A => n5521, Z => n61800);
   U931 : NAND2_X1 port map( A1 => n15013, A2 => n14983, ZN => n8021);
   U932 : NAND2_X1 port map( A1 => n15023, A2 => n14983, ZN => n8045);
   U933 : NAND2_X1 port map( A1 => n15061, A2 => n14983, ZN => n8134);
   U934 : BUF_X1 port map( A => n5553, Z => n61740);
   U935 : BUF_X1 port map( A => n5411, Z => n61920);
   U936 : BUF_X1 port map( A => n5540, Z => n61770);
   U937 : BUF_X1 port map( A => n5428, Z => n61899);
   U938 : BUF_X1 port map( A => n5393, Z => n61947);
   U939 : BUF_X1 port map( A => n5422, Z => n61905);
   U940 : BUF_X1 port map( A => n5396, Z => n61941);
   U941 : INV_X1 port map( A => n5484, ZN => n5342);
   U942 : INV_X1 port map( A => n5493, ZN => n5339);
   U943 : INV_X1 port map( A => n5492, ZN => n5338);
   U944 : INV_X1 port map( A => n5485, ZN => n5343);
   U945 : BUF_X1 port map( A => n5421, Z => n61908);
   U946 : INV_X1 port map( A => n5500, ZN => n5334);
   U947 : INV_X1 port map( A => n5456, ZN => n5307);
   U948 : INV_X1 port map( A => n5536, ZN => n5324);
   U949 : BUF_X1 port map( A => n5416, Z => n59737);
   U950 : INV_X1 port map( A => n5397, ZN => n5297);
   U951 : INV_X1 port map( A => n5386, ZN => n5319);
   U952 : INV_X1 port map( A => n5435, ZN => n5316);
   U953 : INV_X1 port map( A => n5503, ZN => n5331);
   U954 : INV_X1 port map( A => n5440, ZN => n5313);
   U955 : INV_X1 port map( A => n5459, ZN => n5300);
   U956 : INV_X1 port map( A => n5516, ZN => n5326);
   U957 : INV_X1 port map( A => n5448, ZN => n5321);
   U958 : INV_X1 port map( A => n5460, ZN => n5346);
   U959 : INV_X1 port map( A => n5441, ZN => n5315);
   U960 : INV_X1 port map( A => n5449, ZN => n5322);
   U961 : INV_X1 port map( A => n5501, ZN => n5335);
   U962 : INV_X1 port map( A => n5517, ZN => n5327);
   U963 : INV_X1 port map( A => n5454, ZN => n5309);
   U964 : INV_X1 port map( A => n5504, ZN => n5333);
   U965 : INV_X1 port map( A => n5453, ZN => n5308);
   U966 : INV_X1 port map( A => n5436, ZN => n5314);
   U967 : INV_X1 port map( A => n5457, ZN => n5306);
   U968 : INV_X1 port map( A => n5537, ZN => n5325);
   U969 : INV_X1 port map( A => n5398, ZN => n5284);
   U970 : BUF_X1 port map( A => n59965, Z => n59958);
   U971 : BUF_X1 port map( A => n59965, Z => n59959);
   U972 : BUF_X1 port map( A => n59965, Z => n59960);
   U973 : BUF_X1 port map( A => n59965, Z => n59961);
   U974 : BUF_X1 port map( A => n59839, Z => n59832);
   U975 : BUF_X1 port map( A => n59839, Z => n59833);
   U976 : BUF_X1 port map( A => n59839, Z => n59834);
   U977 : BUF_X1 port map( A => n59839, Z => n59835);
   U978 : BUF_X1 port map( A => n59830, Z => n59823);
   U979 : BUF_X1 port map( A => n59830, Z => n59824);
   U980 : BUF_X1 port map( A => n59830, Z => n59825);
   U981 : BUF_X1 port map( A => n59830, Z => n59826);
   U982 : BUF_X1 port map( A => n60676, Z => n60669);
   U983 : BUF_X1 port map( A => n60676, Z => n60670);
   U984 : BUF_X1 port map( A => n60676, Z => n60671);
   U985 : BUF_X1 port map( A => n60676, Z => n60672);
   U986 : BUF_X1 port map( A => n60667, Z => n60660);
   U987 : BUF_X1 port map( A => n60667, Z => n60661);
   U988 : BUF_X1 port map( A => n60667, Z => n60662);
   U989 : BUF_X1 port map( A => n60667, Z => n60663);
   U990 : BUF_X1 port map( A => n60658, Z => n60651);
   U991 : BUF_X1 port map( A => n60658, Z => n60652);
   U992 : BUF_X1 port map( A => n60658, Z => n60653);
   U993 : BUF_X1 port map( A => n60658, Z => n60654);
   U994 : BUF_X1 port map( A => n60649, Z => n60642);
   U995 : BUF_X1 port map( A => n60649, Z => n60643);
   U996 : BUF_X1 port map( A => n60649, Z => n60644);
   U997 : BUF_X1 port map( A => n60649, Z => n60645);
   U998 : BUF_X1 port map( A => n60622, Z => n60615);
   U999 : BUF_X1 port map( A => n60622, Z => n60616);
   U1000 : BUF_X1 port map( A => n60622, Z => n60617);
   U1001 : BUF_X1 port map( A => n60622, Z => n60618);
   U1002 : BUF_X1 port map( A => n60613, Z => n60606);
   U1003 : BUF_X1 port map( A => n60613, Z => n60607);
   U1004 : BUF_X1 port map( A => n60613, Z => n60608);
   U1005 : BUF_X1 port map( A => n60613, Z => n60609);
   U1006 : BUF_X1 port map( A => n60586, Z => n60579);
   U1007 : BUF_X1 port map( A => n60586, Z => n60580);
   U1008 : BUF_X1 port map( A => n60586, Z => n60581);
   U1009 : BUF_X1 port map( A => n60586, Z => n60582);
   U1010 : BUF_X1 port map( A => n60577, Z => n60570);
   U1011 : BUF_X1 port map( A => n60577, Z => n60571);
   U1012 : BUF_X1 port map( A => n60577, Z => n60572);
   U1013 : BUF_X1 port map( A => n60577, Z => n60573);
   U1014 : BUF_X1 port map( A => n60568, Z => n60563);
   U1015 : BUF_X1 port map( A => n60568, Z => n60564);
   U1016 : BUF_X1 port map( A => n60550, Z => n60543);
   U1017 : BUF_X1 port map( A => n60550, Z => n60544);
   U1018 : BUF_X1 port map( A => n60550, Z => n60545);
   U1019 : BUF_X1 port map( A => n60550, Z => n60546);
   U1020 : BUF_X1 port map( A => n60541, Z => n60537);
   U1021 : BUF_X1 port map( A => n60532, Z => n60527);
   U1022 : BUF_X1 port map( A => n60532, Z => n60528);
   U1023 : BUF_X1 port map( A => n60523, Z => n60516);
   U1024 : BUF_X1 port map( A => n60523, Z => n60517);
   U1025 : BUF_X1 port map( A => n60523, Z => n60518);
   U1026 : BUF_X1 port map( A => n60523, Z => n60519);
   U1027 : BUF_X1 port map( A => n60505, Z => n60498);
   U1028 : BUF_X1 port map( A => n60505, Z => n60499);
   U1029 : BUF_X1 port map( A => n60505, Z => n60500);
   U1030 : BUF_X1 port map( A => n60505, Z => n60501);
   U1031 : BUF_X1 port map( A => n60496, Z => n60489);
   U1032 : BUF_X1 port map( A => n60496, Z => n60490);
   U1033 : BUF_X1 port map( A => n60496, Z => n60491);
   U1034 : BUF_X1 port map( A => n60496, Z => n60492);
   U1035 : BUF_X1 port map( A => n60433, Z => n60426);
   U1036 : BUF_X1 port map( A => n60433, Z => n60427);
   U1037 : BUF_X1 port map( A => n60433, Z => n60428);
   U1038 : BUF_X1 port map( A => n60433, Z => n60429);
   U1039 : BUF_X1 port map( A => n60424, Z => n60417);
   U1040 : BUF_X1 port map( A => n60424, Z => n60418);
   U1041 : BUF_X1 port map( A => n60424, Z => n60419);
   U1042 : BUF_X1 port map( A => n60424, Z => n60420);
   U1043 : BUF_X1 port map( A => n60946, Z => n60941);
   U1044 : BUF_X1 port map( A => n60946, Z => n60942);
   U1045 : BUF_X1 port map( A => n60928, Z => n60921);
   U1046 : BUF_X1 port map( A => n60928, Z => n60922);
   U1047 : BUF_X1 port map( A => n60928, Z => n60923);
   U1048 : BUF_X1 port map( A => n60928, Z => n60924);
   U1049 : BUF_X1 port map( A => n60919, Z => n60912);
   U1050 : BUF_X1 port map( A => n60919, Z => n60913);
   U1051 : BUF_X1 port map( A => n60919, Z => n60914);
   U1052 : BUF_X1 port map( A => n60919, Z => n60915);
   U1053 : BUF_X1 port map( A => n60910, Z => n60903);
   U1054 : BUF_X1 port map( A => n60910, Z => n60904);
   U1055 : BUF_X1 port map( A => n60910, Z => n60905);
   U1056 : BUF_X1 port map( A => n60910, Z => n60906);
   U1057 : BUF_X1 port map( A => n60892, Z => n60885);
   U1058 : BUF_X1 port map( A => n60892, Z => n60886);
   U1059 : BUF_X1 port map( A => n60892, Z => n60887);
   U1060 : BUF_X1 port map( A => n60892, Z => n60888);
   U1061 : BUF_X1 port map( A => n60883, Z => n60876);
   U1062 : BUF_X1 port map( A => n60883, Z => n60877);
   U1063 : BUF_X1 port map( A => n60883, Z => n60878);
   U1064 : BUF_X1 port map( A => n60883, Z => n60879);
   U1065 : BUF_X1 port map( A => n60865, Z => n60858);
   U1066 : BUF_X1 port map( A => n60865, Z => n60859);
   U1067 : BUF_X1 port map( A => n60865, Z => n60860);
   U1068 : BUF_X1 port map( A => n60865, Z => n60861);
   U1069 : BUF_X1 port map( A => n60856, Z => n60849);
   U1070 : BUF_X1 port map( A => n60856, Z => n60850);
   U1071 : BUF_X1 port map( A => n60856, Z => n60851);
   U1072 : BUF_X1 port map( A => n60856, Z => n60852);
   U1073 : BUF_X1 port map( A => n60847, Z => n60840);
   U1074 : BUF_X1 port map( A => n60847, Z => n60841);
   U1075 : BUF_X1 port map( A => n60847, Z => n60842);
   U1076 : BUF_X1 port map( A => n60847, Z => n60843);
   U1077 : BUF_X1 port map( A => n60838, Z => n60831);
   U1078 : BUF_X1 port map( A => n60838, Z => n60832);
   U1079 : BUF_X1 port map( A => n60838, Z => n60833);
   U1080 : BUF_X1 port map( A => n60838, Z => n60834);
   U1081 : BUF_X1 port map( A => n60829, Z => n60822);
   U1082 : BUF_X1 port map( A => n60829, Z => n60823);
   U1083 : BUF_X1 port map( A => n60829, Z => n60824);
   U1084 : BUF_X1 port map( A => n60829, Z => n60825);
   U1085 : BUF_X1 port map( A => n60901, Z => n60894);
   U1086 : BUF_X1 port map( A => n60901, Z => n60895);
   U1087 : BUF_X1 port map( A => n60901, Z => n60896);
   U1088 : BUF_X1 port map( A => n60901, Z => n60897);
   U1089 : BUF_X1 port map( A => n60181, Z => n60174);
   U1090 : BUF_X1 port map( A => n60181, Z => n60175);
   U1091 : BUF_X1 port map( A => n60181, Z => n60176);
   U1092 : BUF_X1 port map( A => n60181, Z => n60177);
   U1093 : BUF_X1 port map( A => n60109, Z => n60102);
   U1094 : BUF_X1 port map( A => n60820, Z => n60813);
   U1095 : BUF_X1 port map( A => n60820, Z => n60814);
   U1096 : BUF_X1 port map( A => n60820, Z => n60815);
   U1097 : BUF_X1 port map( A => n60820, Z => n60816);
   U1098 : BUF_X1 port map( A => n60811, Z => n60804);
   U1099 : BUF_X1 port map( A => n60811, Z => n60805);
   U1100 : BUF_X1 port map( A => n60811, Z => n60806);
   U1101 : BUF_X1 port map( A => n60811, Z => n60807);
   U1102 : BUF_X1 port map( A => n60802, Z => n60795);
   U1103 : BUF_X1 port map( A => n60802, Z => n60796);
   U1104 : BUF_X1 port map( A => n60802, Z => n60797);
   U1105 : BUF_X1 port map( A => n60802, Z => n60798);
   U1106 : BUF_X1 port map( A => n60721, Z => n60715);
   U1107 : BUF_X1 port map( A => n60721, Z => n60716);
   U1108 : BUF_X1 port map( A => n60721, Z => n60717);
   U1109 : BUF_X1 port map( A => n60712, Z => n60705);
   U1110 : BUF_X1 port map( A => n60712, Z => n60706);
   U1111 : BUF_X1 port map( A => n60712, Z => n60707);
   U1112 : BUF_X1 port map( A => n60712, Z => n60708);
   U1113 : BUF_X1 port map( A => n59938, Z => n59936);
   U1114 : BUF_X1 port map( A => n59929, Z => n59927);
   U1115 : BUF_X1 port map( A => n59866, Z => n59864);
   U1116 : BUF_X1 port map( A => n59839, Z => n59836);
   U1117 : BUF_X1 port map( A => n59839, Z => n59837);
   U1118 : BUF_X1 port map( A => n59830, Z => n59828);
   U1119 : BUF_X1 port map( A => n60658, Z => n60655);
   U1120 : BUF_X1 port map( A => n60658, Z => n60656);
   U1121 : BUF_X1 port map( A => n60649, Z => n60646);
   U1122 : BUF_X1 port map( A => n60649, Z => n60647);
   U1123 : BUF_X1 port map( A => n60622, Z => n60619);
   U1124 : BUF_X1 port map( A => n60622, Z => n60620);
   U1125 : BUF_X1 port map( A => n60613, Z => n60610);
   U1126 : BUF_X1 port map( A => n60613, Z => n60611);
   U1127 : BUF_X1 port map( A => n60586, Z => n60583);
   U1128 : BUF_X1 port map( A => n60586, Z => n60584);
   U1129 : BUF_X1 port map( A => n60577, Z => n60574);
   U1130 : BUF_X1 port map( A => n60577, Z => n60575);
   U1131 : BUF_X1 port map( A => n60550, Z => n60547);
   U1132 : BUF_X1 port map( A => n60550, Z => n60548);
   U1133 : BUF_X1 port map( A => n60541, Z => n60538);
   U1134 : BUF_X1 port map( A => n60541, Z => n60539);
   U1135 : BUF_X1 port map( A => n60487, Z => n60485);
   U1136 : BUF_X1 port map( A => n60469, Z => n60467);
   U1137 : BUF_X1 port map( A => n60460, Z => n60458);
   U1138 : BUF_X1 port map( A => n60415, Z => n60413);
   U1139 : BUF_X1 port map( A => n60406, Z => n60404);
   U1140 : BUF_X1 port map( A => n60946, Z => n60943);
   U1141 : BUF_X1 port map( A => n60946, Z => n60944);
   U1142 : BUF_X1 port map( A => n60937, Z => n60935);
   U1143 : BUF_X1 port map( A => n60928, Z => n60925);
   U1144 : BUF_X1 port map( A => n60928, Z => n60926);
   U1145 : BUF_X1 port map( A => n60919, Z => n60916);
   U1146 : BUF_X1 port map( A => n60919, Z => n60917);
   U1147 : BUF_X1 port map( A => n60892, Z => n60889);
   U1148 : BUF_X1 port map( A => n60892, Z => n60890);
   U1149 : BUF_X1 port map( A => n60883, Z => n60880);
   U1150 : BUF_X1 port map( A => n60883, Z => n60881);
   U1151 : BUF_X1 port map( A => n60856, Z => n60853);
   U1152 : BUF_X1 port map( A => n60856, Z => n60854);
   U1153 : BUF_X1 port map( A => n60847, Z => n60844);
   U1154 : BUF_X1 port map( A => n60847, Z => n60845);
   U1155 : BUF_X1 port map( A => n60838, Z => n60835);
   U1156 : BUF_X1 port map( A => n60838, Z => n60836);
   U1157 : BUF_X1 port map( A => n60829, Z => n60826);
   U1158 : BUF_X1 port map( A => n60829, Z => n60827);
   U1159 : BUF_X1 port map( A => n60379, Z => n60377);
   U1160 : BUF_X1 port map( A => n60370, Z => n60368);
   U1161 : BUF_X1 port map( A => n60361, Z => n60359);
   U1162 : BUF_X1 port map( A => n60352, Z => n60350);
   U1163 : BUF_X1 port map( A => n60343, Z => n60341);
   U1164 : BUF_X1 port map( A => n60280, Z => n60278);
   U1165 : BUF_X1 port map( A => n60271, Z => n60269);
   U1166 : BUF_X1 port map( A => n60226, Z => n60224);
   U1167 : BUF_X1 port map( A => n60217, Z => n60215);
   U1168 : BUF_X1 port map( A => n60163, Z => n60161);
   U1169 : BUF_X1 port map( A => n60154, Z => n60152);
   U1170 : BUF_X1 port map( A => n60811, Z => n60808);
   U1171 : BUF_X1 port map( A => n60811, Z => n60809);
   U1172 : BUF_X1 port map( A => n60802, Z => n60799);
   U1173 : BUF_X1 port map( A => n60802, Z => n60800);
   U1174 : BUF_X1 port map( A => n60721, Z => n60718);
   U1175 : BUF_X1 port map( A => n60721, Z => n60719);
   U1176 : BUF_X1 port map( A => n60712, Z => n60709);
   U1177 : BUF_X1 port map( A => n60712, Z => n60710);
   U1178 : BUF_X1 port map( A => n60685, Z => n60683);
   U1179 : BUF_X1 port map( A => n60100, Z => n60093);
   U1180 : BUF_X1 port map( A => n60100, Z => n60094);
   U1181 : BUF_X1 port map( A => n60100, Z => n60095);
   U1182 : BUF_X1 port map( A => n60100, Z => n60096);
   U1183 : BUF_X1 port map( A => n60091, Z => n60084);
   U1184 : BUF_X1 port map( A => n60091, Z => n60085);
   U1185 : BUF_X1 port map( A => n60091, Z => n60086);
   U1186 : BUF_X1 port map( A => n60091, Z => n60087);
   U1187 : BUF_X1 port map( A => n60082, Z => n60075);
   U1188 : BUF_X1 port map( A => n60082, Z => n60076);
   U1189 : BUF_X1 port map( A => n60082, Z => n60077);
   U1190 : BUF_X1 port map( A => n60082, Z => n60078);
   U1191 : BUF_X1 port map( A => n60073, Z => n60066);
   U1192 : BUF_X1 port map( A => n60073, Z => n60067);
   U1193 : BUF_X1 port map( A => n60073, Z => n60068);
   U1194 : BUF_X1 port map( A => n60073, Z => n60069);
   U1195 : BUF_X1 port map( A => n60064, Z => n60057);
   U1196 : BUF_X1 port map( A => n60064, Z => n60058);
   U1197 : BUF_X1 port map( A => n60064, Z => n60059);
   U1198 : BUF_X1 port map( A => n60064, Z => n60060);
   U1199 : BUF_X1 port map( A => n60055, Z => n60048);
   U1200 : BUF_X1 port map( A => n60055, Z => n60049);
   U1201 : BUF_X1 port map( A => n60055, Z => n60050);
   U1202 : BUF_X1 port map( A => n60055, Z => n60051);
   U1203 : BUF_X1 port map( A => n60046, Z => n60039);
   U1204 : BUF_X1 port map( A => n60046, Z => n60040);
   U1205 : BUF_X1 port map( A => n60046, Z => n60041);
   U1206 : BUF_X1 port map( A => n60046, Z => n60042);
   U1207 : BUF_X1 port map( A => n60037, Z => n60030);
   U1208 : BUF_X1 port map( A => n60037, Z => n60031);
   U1209 : BUF_X1 port map( A => n60037, Z => n60032);
   U1210 : BUF_X1 port map( A => n60037, Z => n60033);
   U1211 : BUF_X1 port map( A => n60028, Z => n60021);
   U1212 : BUF_X1 port map( A => n60028, Z => n60022);
   U1213 : BUF_X1 port map( A => n60028, Z => n60023);
   U1214 : BUF_X1 port map( A => n60028, Z => n60024);
   U1215 : BUF_X1 port map( A => n60019, Z => n60012);
   U1216 : BUF_X1 port map( A => n60019, Z => n60013);
   U1217 : BUF_X1 port map( A => n60019, Z => n60014);
   U1218 : BUF_X1 port map( A => n60019, Z => n60015);
   U1219 : BUF_X1 port map( A => n60010, Z => n60003);
   U1220 : BUF_X1 port map( A => n60010, Z => n60004);
   U1221 : BUF_X1 port map( A => n60010, Z => n60005);
   U1222 : BUF_X1 port map( A => n60010, Z => n60006);
   U1223 : BUF_X1 port map( A => n60001, Z => n59994);
   U1224 : BUF_X1 port map( A => n60001, Z => n59995);
   U1225 : BUF_X1 port map( A => n60001, Z => n59996);
   U1226 : BUF_X1 port map( A => n60001, Z => n59997);
   U1227 : BUF_X1 port map( A => n59992, Z => n59985);
   U1228 : BUF_X1 port map( A => n59992, Z => n59986);
   U1229 : BUF_X1 port map( A => n59992, Z => n59987);
   U1230 : BUF_X1 port map( A => n59992, Z => n59988);
   U1231 : BUF_X1 port map( A => n59983, Z => n59976);
   U1232 : BUF_X1 port map( A => n59983, Z => n59977);
   U1233 : BUF_X1 port map( A => n59983, Z => n59978);
   U1234 : BUF_X1 port map( A => n59983, Z => n59979);
   U1235 : BUF_X1 port map( A => n59974, Z => n59967);
   U1236 : BUF_X1 port map( A => n59974, Z => n59968);
   U1237 : BUF_X1 port map( A => n59974, Z => n59969);
   U1238 : BUF_X1 port map( A => n59974, Z => n59970);
   U1239 : BUF_X1 port map( A => n59956, Z => n59949);
   U1240 : BUF_X1 port map( A => n59956, Z => n59950);
   U1241 : BUF_X1 port map( A => n59956, Z => n59951);
   U1242 : BUF_X1 port map( A => n59956, Z => n59952);
   U1243 : BUF_X1 port map( A => n59947, Z => n59940);
   U1244 : BUF_X1 port map( A => n59947, Z => n59941);
   U1245 : BUF_X1 port map( A => n59947, Z => n59942);
   U1246 : BUF_X1 port map( A => n59947, Z => n59943);
   U1247 : BUF_X1 port map( A => n59938, Z => n59931);
   U1248 : BUF_X1 port map( A => n59938, Z => n59932);
   U1249 : BUF_X1 port map( A => n59938, Z => n59933);
   U1250 : BUF_X1 port map( A => n59938, Z => n59934);
   U1251 : BUF_X1 port map( A => n59929, Z => n59922);
   U1252 : BUF_X1 port map( A => n59929, Z => n59923);
   U1253 : BUF_X1 port map( A => n59929, Z => n59924);
   U1254 : BUF_X1 port map( A => n59929, Z => n59925);
   U1255 : BUF_X1 port map( A => n59929, Z => n59926);
   U1256 : BUF_X1 port map( A => n59920, Z => n59913);
   U1257 : BUF_X1 port map( A => n59920, Z => n59914);
   U1258 : BUF_X1 port map( A => n59920, Z => n59915);
   U1259 : BUF_X1 port map( A => n59920, Z => n59916);
   U1260 : BUF_X1 port map( A => n59911, Z => n59904);
   U1261 : BUF_X1 port map( A => n59911, Z => n59905);
   U1262 : BUF_X1 port map( A => n59911, Z => n59906);
   U1263 : BUF_X1 port map( A => n59911, Z => n59907);
   U1264 : BUF_X1 port map( A => n59902, Z => n59895);
   U1265 : BUF_X1 port map( A => n59902, Z => n59896);
   U1266 : BUF_X1 port map( A => n59902, Z => n59897);
   U1267 : BUF_X1 port map( A => n59902, Z => n59898);
   U1268 : BUF_X1 port map( A => n59893, Z => n59886);
   U1269 : BUF_X1 port map( A => n59893, Z => n59887);
   U1270 : BUF_X1 port map( A => n59893, Z => n59888);
   U1271 : BUF_X1 port map( A => n59893, Z => n59889);
   U1272 : BUF_X1 port map( A => n59884, Z => n59877);
   U1273 : BUF_X1 port map( A => n59884, Z => n59878);
   U1274 : BUF_X1 port map( A => n59884, Z => n59879);
   U1275 : BUF_X1 port map( A => n59884, Z => n59880);
   U1276 : BUF_X1 port map( A => n59875, Z => n59868);
   U1277 : BUF_X1 port map( A => n59875, Z => n59869);
   U1278 : BUF_X1 port map( A => n59875, Z => n59870);
   U1279 : BUF_X1 port map( A => n59875, Z => n59871);
   U1280 : BUF_X1 port map( A => n59866, Z => n59859);
   U1281 : BUF_X1 port map( A => n59866, Z => n59860);
   U1282 : BUF_X1 port map( A => n59866, Z => n59861);
   U1283 : BUF_X1 port map( A => n59866, Z => n59862);
   U1284 : BUF_X1 port map( A => n59866, Z => n59863);
   U1285 : BUF_X1 port map( A => n59857, Z => n59850);
   U1286 : BUF_X1 port map( A => n59857, Z => n59851);
   U1287 : BUF_X1 port map( A => n59857, Z => n59852);
   U1288 : BUF_X1 port map( A => n59857, Z => n59853);
   U1289 : BUF_X1 port map( A => n59848, Z => n59841);
   U1290 : BUF_X1 port map( A => n59848, Z => n59842);
   U1291 : BUF_X1 port map( A => n59848, Z => n59843);
   U1292 : BUF_X1 port map( A => n59848, Z => n59844);
   U1293 : BUF_X1 port map( A => n59830, Z => n59827);
   U1294 : BUF_X1 port map( A => n59821, Z => n59814);
   U1295 : BUF_X1 port map( A => n59821, Z => n59815);
   U1296 : BUF_X1 port map( A => n59821, Z => n59816);
   U1297 : BUF_X1 port map( A => n59821, Z => n59817);
   U1298 : BUF_X1 port map( A => n60640, Z => n60633);
   U1299 : BUF_X1 port map( A => n60640, Z => n60634);
   U1300 : BUF_X1 port map( A => n60640, Z => n60635);
   U1301 : BUF_X1 port map( A => n60640, Z => n60636);
   U1302 : BUF_X1 port map( A => n60631, Z => n60624);
   U1303 : BUF_X1 port map( A => n60631, Z => n60625);
   U1304 : BUF_X1 port map( A => n60631, Z => n60626);
   U1305 : BUF_X1 port map( A => n60631, Z => n60627);
   U1306 : BUF_X1 port map( A => n60604, Z => n60597);
   U1307 : BUF_X1 port map( A => n60604, Z => n60598);
   U1308 : BUF_X1 port map( A => n60604, Z => n60599);
   U1309 : BUF_X1 port map( A => n60604, Z => n60600);
   U1310 : BUF_X1 port map( A => n60595, Z => n60588);
   U1311 : BUF_X1 port map( A => n60595, Z => n60589);
   U1312 : BUF_X1 port map( A => n60595, Z => n60590);
   U1313 : BUF_X1 port map( A => n60595, Z => n60591);
   U1314 : BUF_X1 port map( A => n60568, Z => n60561);
   U1315 : BUF_X1 port map( A => n60568, Z => n60562);
   U1316 : BUF_X1 port map( A => n60559, Z => n60552);
   U1317 : BUF_X1 port map( A => n60559, Z => n60553);
   U1318 : BUF_X1 port map( A => n60559, Z => n60554);
   U1319 : BUF_X1 port map( A => n60559, Z => n60555);
   U1320 : BUF_X1 port map( A => n60559, Z => n60556);
   U1321 : BUF_X1 port map( A => n60541, Z => n60534);
   U1322 : BUF_X1 port map( A => n60541, Z => n60535);
   U1323 : BUF_X1 port map( A => n60541, Z => n60536);
   U1324 : BUF_X1 port map( A => n60532, Z => n60525);
   U1325 : BUF_X1 port map( A => n60532, Z => n60526);
   U1326 : BUF_X1 port map( A => n60514, Z => n60507);
   U1327 : BUF_X1 port map( A => n60514, Z => n60508);
   U1328 : BUF_X1 port map( A => n60514, Z => n60509);
   U1329 : BUF_X1 port map( A => n60514, Z => n60510);
   U1330 : BUF_X1 port map( A => n60487, Z => n60480);
   U1331 : BUF_X1 port map( A => n60487, Z => n60481);
   U1332 : BUF_X1 port map( A => n60487, Z => n60482);
   U1333 : BUF_X1 port map( A => n60487, Z => n60483);
   U1334 : BUF_X1 port map( A => n60487, Z => n60484);
   U1335 : BUF_X1 port map( A => n60478, Z => n60471);
   U1336 : BUF_X1 port map( A => n60478, Z => n60472);
   U1337 : BUF_X1 port map( A => n60478, Z => n60473);
   U1338 : BUF_X1 port map( A => n60478, Z => n60474);
   U1339 : BUF_X1 port map( A => n60469, Z => n60462);
   U1340 : BUF_X1 port map( A => n60469, Z => n60463);
   U1341 : BUF_X1 port map( A => n60469, Z => n60464);
   U1342 : BUF_X1 port map( A => n60469, Z => n60465);
   U1343 : BUF_X1 port map( A => n60469, Z => n60466);
   U1344 : BUF_X1 port map( A => n60460, Z => n60453);
   U1345 : BUF_X1 port map( A => n60460, Z => n60454);
   U1346 : BUF_X1 port map( A => n60460, Z => n60455);
   U1347 : BUF_X1 port map( A => n60460, Z => n60456);
   U1348 : BUF_X1 port map( A => n60460, Z => n60457);
   U1349 : BUF_X1 port map( A => n60451, Z => n60444);
   U1350 : BUF_X1 port map( A => n60451, Z => n60445);
   U1351 : BUF_X1 port map( A => n60451, Z => n60446);
   U1352 : BUF_X1 port map( A => n60451, Z => n60447);
   U1353 : BUF_X1 port map( A => n60442, Z => n60435);
   U1354 : BUF_X1 port map( A => n60442, Z => n60436);
   U1355 : BUF_X1 port map( A => n60442, Z => n60437);
   U1356 : BUF_X1 port map( A => n60442, Z => n60438);
   U1357 : BUF_X1 port map( A => n60415, Z => n60408);
   U1358 : BUF_X1 port map( A => n60415, Z => n60409);
   U1359 : BUF_X1 port map( A => n60415, Z => n60410);
   U1360 : BUF_X1 port map( A => n60415, Z => n60411);
   U1361 : BUF_X1 port map( A => n60415, Z => n60412);
   U1362 : BUF_X1 port map( A => n60406, Z => n60399);
   U1363 : BUF_X1 port map( A => n60406, Z => n60400);
   U1364 : BUF_X1 port map( A => n60406, Z => n60401);
   U1365 : BUF_X1 port map( A => n60406, Z => n60402);
   U1366 : BUF_X1 port map( A => n60406, Z => n60403);
   U1367 : BUF_X1 port map( A => n60397, Z => n60390);
   U1368 : BUF_X1 port map( A => n60397, Z => n60391);
   U1369 : BUF_X1 port map( A => n60397, Z => n60392);
   U1370 : BUF_X1 port map( A => n60397, Z => n60393);
   U1371 : BUF_X1 port map( A => n61244, Z => n61237);
   U1372 : BUF_X1 port map( A => n61244, Z => n61238);
   U1373 : BUF_X1 port map( A => n61244, Z => n61239);
   U1374 : BUF_X1 port map( A => n61244, Z => n61240);
   U1375 : BUF_X1 port map( A => n60955, Z => n60948);
   U1376 : BUF_X1 port map( A => n60955, Z => n60949);
   U1377 : BUF_X1 port map( A => n60955, Z => n60950);
   U1378 : BUF_X1 port map( A => n60955, Z => n60951);
   U1379 : BUF_X1 port map( A => n60946, Z => n60939);
   U1380 : BUF_X1 port map( A => n60946, Z => n60940);
   U1381 : BUF_X1 port map( A => n60937, Z => n60930);
   U1382 : BUF_X1 port map( A => n60937, Z => n60931);
   U1383 : BUF_X1 port map( A => n60937, Z => n60932);
   U1384 : BUF_X1 port map( A => n60937, Z => n60933);
   U1385 : BUF_X1 port map( A => n60937, Z => n60934);
   U1386 : BUF_X1 port map( A => n60874, Z => n60867);
   U1387 : BUF_X1 port map( A => n60874, Z => n60868);
   U1388 : BUF_X1 port map( A => n60874, Z => n60869);
   U1389 : BUF_X1 port map( A => n60874, Z => n60870);
   U1390 : BUF_X1 port map( A => n60388, Z => n60381);
   U1391 : BUF_X1 port map( A => n60388, Z => n60382);
   U1392 : BUF_X1 port map( A => n60388, Z => n60383);
   U1393 : BUF_X1 port map( A => n60388, Z => n60384);
   U1394 : BUF_X1 port map( A => n60379, Z => n60372);
   U1395 : BUF_X1 port map( A => n60379, Z => n60373);
   U1396 : BUF_X1 port map( A => n60379, Z => n60374);
   U1397 : BUF_X1 port map( A => n60379, Z => n60375);
   U1398 : BUF_X1 port map( A => n60379, Z => n60376);
   U1399 : BUF_X1 port map( A => n60370, Z => n60363);
   U1400 : BUF_X1 port map( A => n60370, Z => n60364);
   U1401 : BUF_X1 port map( A => n60370, Z => n60365);
   U1402 : BUF_X1 port map( A => n60370, Z => n60366);
   U1403 : BUF_X1 port map( A => n60370, Z => n60367);
   U1404 : BUF_X1 port map( A => n60361, Z => n60354);
   U1405 : BUF_X1 port map( A => n60361, Z => n60355);
   U1406 : BUF_X1 port map( A => n60361, Z => n60356);
   U1407 : BUF_X1 port map( A => n60361, Z => n60357);
   U1408 : BUF_X1 port map( A => n60361, Z => n60358);
   U1409 : BUF_X1 port map( A => n60352, Z => n60345);
   U1410 : BUF_X1 port map( A => n60352, Z => n60346);
   U1411 : BUF_X1 port map( A => n60352, Z => n60347);
   U1412 : BUF_X1 port map( A => n60352, Z => n60348);
   U1413 : BUF_X1 port map( A => n60352, Z => n60349);
   U1414 : BUF_X1 port map( A => n60343, Z => n60336);
   U1415 : BUF_X1 port map( A => n60343, Z => n60337);
   U1416 : BUF_X1 port map( A => n60343, Z => n60338);
   U1417 : BUF_X1 port map( A => n60343, Z => n60339);
   U1418 : BUF_X1 port map( A => n60343, Z => n60340);
   U1419 : BUF_X1 port map( A => n60334, Z => n60327);
   U1420 : BUF_X1 port map( A => n60334, Z => n60328);
   U1421 : BUF_X1 port map( A => n60334, Z => n60329);
   U1422 : BUF_X1 port map( A => n60334, Z => n60330);
   U1423 : BUF_X1 port map( A => n60325, Z => n60318);
   U1424 : BUF_X1 port map( A => n60325, Z => n60319);
   U1425 : BUF_X1 port map( A => n60325, Z => n60320);
   U1426 : BUF_X1 port map( A => n60325, Z => n60321);
   U1427 : BUF_X1 port map( A => n60316, Z => n60309);
   U1428 : BUF_X1 port map( A => n60316, Z => n60310);
   U1429 : BUF_X1 port map( A => n60316, Z => n60311);
   U1430 : BUF_X1 port map( A => n60316, Z => n60312);
   U1431 : BUF_X1 port map( A => n60307, Z => n60300);
   U1432 : BUF_X1 port map( A => n60307, Z => n60301);
   U1433 : BUF_X1 port map( A => n60307, Z => n60302);
   U1434 : BUF_X1 port map( A => n60307, Z => n60303);
   U1435 : BUF_X1 port map( A => n60298, Z => n60291);
   U1436 : BUF_X1 port map( A => n60298, Z => n60292);
   U1437 : BUF_X1 port map( A => n60298, Z => n60293);
   U1438 : BUF_X1 port map( A => n60298, Z => n60294);
   U1439 : BUF_X1 port map( A => n60289, Z => n60282);
   U1440 : BUF_X1 port map( A => n60289, Z => n60283);
   U1441 : BUF_X1 port map( A => n60289, Z => n60284);
   U1442 : BUF_X1 port map( A => n60289, Z => n60285);
   U1443 : BUF_X1 port map( A => n60280, Z => n60273);
   U1444 : BUF_X1 port map( A => n60280, Z => n60274);
   U1445 : BUF_X1 port map( A => n60280, Z => n60275);
   U1446 : BUF_X1 port map( A => n60280, Z => n60276);
   U1447 : BUF_X1 port map( A => n60280, Z => n60277);
   U1448 : BUF_X1 port map( A => n60271, Z => n60264);
   U1449 : BUF_X1 port map( A => n60271, Z => n60265);
   U1450 : BUF_X1 port map( A => n60271, Z => n60266);
   U1451 : BUF_X1 port map( A => n60271, Z => n60267);
   U1452 : BUF_X1 port map( A => n60271, Z => n60268);
   U1453 : BUF_X1 port map( A => n60262, Z => n60255);
   U1454 : BUF_X1 port map( A => n60262, Z => n60256);
   U1455 : BUF_X1 port map( A => n60262, Z => n60257);
   U1456 : BUF_X1 port map( A => n60262, Z => n60258);
   U1457 : BUF_X1 port map( A => n60253, Z => n60246);
   U1458 : BUF_X1 port map( A => n60253, Z => n60247);
   U1459 : BUF_X1 port map( A => n60253, Z => n60248);
   U1460 : BUF_X1 port map( A => n60253, Z => n60249);
   U1461 : BUF_X1 port map( A => n60244, Z => n60237);
   U1462 : BUF_X1 port map( A => n60244, Z => n60238);
   U1463 : BUF_X1 port map( A => n60244, Z => n60239);
   U1464 : BUF_X1 port map( A => n60244, Z => n60240);
   U1465 : BUF_X1 port map( A => n60235, Z => n60228);
   U1466 : BUF_X1 port map( A => n60235, Z => n60229);
   U1467 : BUF_X1 port map( A => n60235, Z => n60230);
   U1468 : BUF_X1 port map( A => n60235, Z => n60231);
   U1469 : BUF_X1 port map( A => n60226, Z => n60219);
   U1470 : BUF_X1 port map( A => n60226, Z => n60220);
   U1471 : BUF_X1 port map( A => n60226, Z => n60221);
   U1472 : BUF_X1 port map( A => n60226, Z => n60222);
   U1473 : BUF_X1 port map( A => n60226, Z => n60223);
   U1474 : BUF_X1 port map( A => n60217, Z => n60210);
   U1475 : BUF_X1 port map( A => n60217, Z => n60211);
   U1476 : BUF_X1 port map( A => n60217, Z => n60212);
   U1477 : BUF_X1 port map( A => n60217, Z => n60213);
   U1478 : BUF_X1 port map( A => n60217, Z => n60214);
   U1479 : BUF_X1 port map( A => n60208, Z => n60201);
   U1480 : BUF_X1 port map( A => n60208, Z => n60202);
   U1481 : BUF_X1 port map( A => n60208, Z => n60203);
   U1482 : BUF_X1 port map( A => n60208, Z => n60204);
   U1483 : BUF_X1 port map( A => n60199, Z => n60192);
   U1484 : BUF_X1 port map( A => n60199, Z => n60193);
   U1485 : BUF_X1 port map( A => n60199, Z => n60194);
   U1486 : BUF_X1 port map( A => n60199, Z => n60195);
   U1487 : BUF_X1 port map( A => n60190, Z => n60183);
   U1488 : BUF_X1 port map( A => n60190, Z => n60184);
   U1489 : BUF_X1 port map( A => n60190, Z => n60185);
   U1490 : BUF_X1 port map( A => n60190, Z => n60186);
   U1491 : BUF_X1 port map( A => n60172, Z => n60165);
   U1492 : BUF_X1 port map( A => n60172, Z => n60166);
   U1493 : BUF_X1 port map( A => n60172, Z => n60167);
   U1494 : BUF_X1 port map( A => n60172, Z => n60168);
   U1495 : BUF_X1 port map( A => n60163, Z => n60156);
   U1496 : BUF_X1 port map( A => n60163, Z => n60157);
   U1497 : BUF_X1 port map( A => n60163, Z => n60158);
   U1498 : BUF_X1 port map( A => n60163, Z => n60159);
   U1499 : BUF_X1 port map( A => n60163, Z => n60160);
   U1500 : BUF_X1 port map( A => n60154, Z => n60147);
   U1501 : BUF_X1 port map( A => n60154, Z => n60148);
   U1502 : BUF_X1 port map( A => n60154, Z => n60149);
   U1503 : BUF_X1 port map( A => n60154, Z => n60150);
   U1504 : BUF_X1 port map( A => n60154, Z => n60151);
   U1505 : BUF_X1 port map( A => n60145, Z => n60138);
   U1506 : BUF_X1 port map( A => n60145, Z => n60139);
   U1507 : BUF_X1 port map( A => n60145, Z => n60140);
   U1508 : BUF_X1 port map( A => n60145, Z => n60141);
   U1509 : BUF_X1 port map( A => n60136, Z => n60129);
   U1510 : BUF_X1 port map( A => n60136, Z => n60130);
   U1511 : BUF_X1 port map( A => n60136, Z => n60131);
   U1512 : BUF_X1 port map( A => n60136, Z => n60132);
   U1513 : BUF_X1 port map( A => n60127, Z => n60120);
   U1514 : BUF_X1 port map( A => n60127, Z => n60121);
   U1515 : BUF_X1 port map( A => n60127, Z => n60122);
   U1516 : BUF_X1 port map( A => n60127, Z => n60123);
   U1517 : BUF_X1 port map( A => n60118, Z => n60111);
   U1518 : BUF_X1 port map( A => n60118, Z => n60112);
   U1519 : BUF_X1 port map( A => n60118, Z => n60113);
   U1520 : BUF_X1 port map( A => n60118, Z => n60114);
   U1521 : BUF_X1 port map( A => n60109, Z => n60103);
   U1522 : BUF_X1 port map( A => n60109, Z => n60104);
   U1523 : BUF_X1 port map( A => n60109, Z => n60105);
   U1524 : BUF_X1 port map( A => n60793, Z => n60786);
   U1525 : BUF_X1 port map( A => n60793, Z => n60787);
   U1526 : BUF_X1 port map( A => n60793, Z => n60788);
   U1527 : BUF_X1 port map( A => n60793, Z => n60789);
   U1528 : BUF_X1 port map( A => n60784, Z => n60777);
   U1529 : BUF_X1 port map( A => n60784, Z => n60778);
   U1530 : BUF_X1 port map( A => n60784, Z => n60779);
   U1531 : BUF_X1 port map( A => n60784, Z => n60780);
   U1532 : BUF_X1 port map( A => n60775, Z => n60768);
   U1533 : BUF_X1 port map( A => n60775, Z => n60769);
   U1534 : BUF_X1 port map( A => n60775, Z => n60770);
   U1535 : BUF_X1 port map( A => n60775, Z => n60771);
   U1536 : BUF_X1 port map( A => n60766, Z => n60759);
   U1537 : BUF_X1 port map( A => n60766, Z => n60760);
   U1538 : BUF_X1 port map( A => n60766, Z => n60761);
   U1539 : BUF_X1 port map( A => n60766, Z => n60762);
   U1540 : BUF_X1 port map( A => n60757, Z => n60750);
   U1541 : BUF_X1 port map( A => n60757, Z => n60751);
   U1542 : BUF_X1 port map( A => n60757, Z => n60752);
   U1543 : BUF_X1 port map( A => n60757, Z => n60753);
   U1544 : BUF_X1 port map( A => n60748, Z => n60741);
   U1545 : BUF_X1 port map( A => n60748, Z => n60742);
   U1546 : BUF_X1 port map( A => n60748, Z => n60743);
   U1547 : BUF_X1 port map( A => n60748, Z => n60744);
   U1548 : BUF_X1 port map( A => n60739, Z => n60732);
   U1549 : BUF_X1 port map( A => n60739, Z => n60733);
   U1550 : BUF_X1 port map( A => n60739, Z => n60734);
   U1551 : BUF_X1 port map( A => n60739, Z => n60735);
   U1552 : BUF_X1 port map( A => n60730, Z => n60723);
   U1553 : BUF_X1 port map( A => n60730, Z => n60724);
   U1554 : BUF_X1 port map( A => n60730, Z => n60725);
   U1555 : BUF_X1 port map( A => n60730, Z => n60726);
   U1556 : BUF_X1 port map( A => n60721, Z => n60714);
   U1557 : BUF_X1 port map( A => n60703, Z => n60696);
   U1558 : BUF_X1 port map( A => n60703, Z => n60697);
   U1559 : BUF_X1 port map( A => n60703, Z => n60698);
   U1560 : BUF_X1 port map( A => n60703, Z => n60699);
   U1561 : BUF_X1 port map( A => n60694, Z => n60687);
   U1562 : BUF_X1 port map( A => n60694, Z => n60688);
   U1563 : BUF_X1 port map( A => n60694, Z => n60689);
   U1564 : BUF_X1 port map( A => n60694, Z => n60690);
   U1565 : BUF_X1 port map( A => n60685, Z => n60678);
   U1566 : BUF_X1 port map( A => n60685, Z => n60679);
   U1567 : BUF_X1 port map( A => n60685, Z => n60680);
   U1568 : BUF_X1 port map( A => n60685, Z => n60681);
   U1569 : BUF_X1 port map( A => n60685, Z => n60682);
   U1570 : BUF_X1 port map( A => n60100, Z => n60097);
   U1571 : BUF_X1 port map( A => n60100, Z => n60098);
   U1572 : BUF_X1 port map( A => n60091, Z => n60088);
   U1573 : BUF_X1 port map( A => n60091, Z => n60089);
   U1574 : BUF_X1 port map( A => n60082, Z => n60079);
   U1575 : BUF_X1 port map( A => n60082, Z => n60080);
   U1576 : BUF_X1 port map( A => n60073, Z => n60070);
   U1577 : BUF_X1 port map( A => n60073, Z => n60071);
   U1578 : BUF_X1 port map( A => n60064, Z => n60061);
   U1579 : BUF_X1 port map( A => n60064, Z => n60062);
   U1580 : BUF_X1 port map( A => n60055, Z => n60052);
   U1581 : BUF_X1 port map( A => n60055, Z => n60053);
   U1582 : BUF_X1 port map( A => n60046, Z => n60043);
   U1583 : BUF_X1 port map( A => n60046, Z => n60044);
   U1584 : BUF_X1 port map( A => n60037, Z => n60034);
   U1585 : BUF_X1 port map( A => n60037, Z => n60035);
   U1586 : BUF_X1 port map( A => n60028, Z => n60025);
   U1587 : BUF_X1 port map( A => n60028, Z => n60026);
   U1588 : BUF_X1 port map( A => n60019, Z => n60016);
   U1589 : BUF_X1 port map( A => n60019, Z => n60017);
   U1590 : BUF_X1 port map( A => n60010, Z => n60007);
   U1591 : BUF_X1 port map( A => n60010, Z => n60008);
   U1592 : BUF_X1 port map( A => n60001, Z => n59998);
   U1593 : BUF_X1 port map( A => n60001, Z => n59999);
   U1594 : BUF_X1 port map( A => n59992, Z => n59989);
   U1595 : BUF_X1 port map( A => n59992, Z => n59990);
   U1596 : BUF_X1 port map( A => n59983, Z => n59980);
   U1597 : BUF_X1 port map( A => n59983, Z => n59981);
   U1598 : BUF_X1 port map( A => n59974, Z => n59971);
   U1599 : BUF_X1 port map( A => n59974, Z => n59972);
   U1600 : BUF_X1 port map( A => n59965, Z => n59962);
   U1601 : BUF_X1 port map( A => n59965, Z => n59963);
   U1602 : BUF_X1 port map( A => n59956, Z => n59953);
   U1603 : BUF_X1 port map( A => n59956, Z => n59954);
   U1604 : BUF_X1 port map( A => n59947, Z => n59944);
   U1605 : BUF_X1 port map( A => n59947, Z => n59945);
   U1606 : BUF_X1 port map( A => n59938, Z => n59935);
   U1607 : BUF_X1 port map( A => n59920, Z => n59917);
   U1608 : BUF_X1 port map( A => n59920, Z => n59918);
   U1609 : BUF_X1 port map( A => n59911, Z => n59908);
   U1610 : BUF_X1 port map( A => n59911, Z => n59909);
   U1611 : BUF_X1 port map( A => n59902, Z => n59899);
   U1612 : BUF_X1 port map( A => n59902, Z => n59900);
   U1613 : BUF_X1 port map( A => n59893, Z => n59890);
   U1614 : BUF_X1 port map( A => n59893, Z => n59891);
   U1615 : BUF_X1 port map( A => n59884, Z => n59881);
   U1616 : BUF_X1 port map( A => n59884, Z => n59882);
   U1617 : BUF_X1 port map( A => n59875, Z => n59872);
   U1618 : BUF_X1 port map( A => n59875, Z => n59873);
   U1619 : BUF_X1 port map( A => n59857, Z => n59854);
   U1620 : BUF_X1 port map( A => n59857, Z => n59855);
   U1621 : BUF_X1 port map( A => n59848, Z => n59845);
   U1622 : BUF_X1 port map( A => n59848, Z => n59846);
   U1623 : BUF_X1 port map( A => n59821, Z => n59818);
   U1624 : BUF_X1 port map( A => n59821, Z => n59819);
   U1625 : BUF_X1 port map( A => n60676, Z => n60673);
   U1626 : BUF_X1 port map( A => n60676, Z => n60674);
   U1627 : BUF_X1 port map( A => n60667, Z => n60664);
   U1628 : BUF_X1 port map( A => n60667, Z => n60665);
   U1629 : BUF_X1 port map( A => n60640, Z => n60637);
   U1630 : BUF_X1 port map( A => n60640, Z => n60638);
   U1631 : BUF_X1 port map( A => n60631, Z => n60628);
   U1632 : BUF_X1 port map( A => n60631, Z => n60629);
   U1633 : BUF_X1 port map( A => n60604, Z => n60601);
   U1634 : BUF_X1 port map( A => n60604, Z => n60602);
   U1635 : BUF_X1 port map( A => n60595, Z => n60592);
   U1636 : BUF_X1 port map( A => n60595, Z => n60593);
   U1637 : BUF_X1 port map( A => n60568, Z => n60565);
   U1638 : BUF_X1 port map( A => n60568, Z => n60566);
   U1639 : BUF_X1 port map( A => n60559, Z => n60557);
   U1640 : BUF_X1 port map( A => n60532, Z => n60529);
   U1641 : BUF_X1 port map( A => n60532, Z => n60530);
   U1642 : BUF_X1 port map( A => n60523, Z => n60520);
   U1643 : BUF_X1 port map( A => n60523, Z => n60521);
   U1644 : BUF_X1 port map( A => n60514, Z => n60511);
   U1645 : BUF_X1 port map( A => n60514, Z => n60512);
   U1646 : BUF_X1 port map( A => n60505, Z => n60502);
   U1647 : BUF_X1 port map( A => n60505, Z => n60503);
   U1648 : BUF_X1 port map( A => n60496, Z => n60493);
   U1649 : BUF_X1 port map( A => n60496, Z => n60494);
   U1650 : BUF_X1 port map( A => n60478, Z => n60475);
   U1651 : BUF_X1 port map( A => n60478, Z => n60476);
   U1652 : BUF_X1 port map( A => n60451, Z => n60448);
   U1653 : BUF_X1 port map( A => n60451, Z => n60449);
   U1654 : BUF_X1 port map( A => n60442, Z => n60439);
   U1655 : BUF_X1 port map( A => n60442, Z => n60440);
   U1656 : BUF_X1 port map( A => n60433, Z => n60430);
   U1657 : BUF_X1 port map( A => n60433, Z => n60431);
   U1658 : BUF_X1 port map( A => n60424, Z => n60421);
   U1659 : BUF_X1 port map( A => n60424, Z => n60422);
   U1660 : BUF_X1 port map( A => n60397, Z => n60394);
   U1661 : BUF_X1 port map( A => n60397, Z => n60395);
   U1662 : BUF_X1 port map( A => n61244, Z => n61241);
   U1663 : BUF_X1 port map( A => n61244, Z => n61242);
   U1664 : BUF_X1 port map( A => n60955, Z => n60952);
   U1665 : BUF_X1 port map( A => n60955, Z => n60953);
   U1666 : BUF_X1 port map( A => n60910, Z => n60907);
   U1667 : BUF_X1 port map( A => n60910, Z => n60908);
   U1668 : BUF_X1 port map( A => n60874, Z => n60871);
   U1669 : BUF_X1 port map( A => n60874, Z => n60872);
   U1670 : BUF_X1 port map( A => n60865, Z => n60862);
   U1671 : BUF_X1 port map( A => n60865, Z => n60863);
   U1672 : BUF_X1 port map( A => n60901, Z => n60898);
   U1673 : BUF_X1 port map( A => n60901, Z => n60899);
   U1674 : BUF_X1 port map( A => n60388, Z => n60385);
   U1675 : BUF_X1 port map( A => n60388, Z => n60386);
   U1676 : BUF_X1 port map( A => n60334, Z => n60331);
   U1677 : BUF_X1 port map( A => n60334, Z => n60332);
   U1678 : BUF_X1 port map( A => n60325, Z => n60322);
   U1679 : BUF_X1 port map( A => n60325, Z => n60323);
   U1680 : BUF_X1 port map( A => n60316, Z => n60313);
   U1681 : BUF_X1 port map( A => n60316, Z => n60314);
   U1682 : BUF_X1 port map( A => n60307, Z => n60304);
   U1683 : BUF_X1 port map( A => n60307, Z => n60305);
   U1684 : BUF_X1 port map( A => n60298, Z => n60295);
   U1685 : BUF_X1 port map( A => n60298, Z => n60296);
   U1686 : BUF_X1 port map( A => n60289, Z => n60286);
   U1687 : BUF_X1 port map( A => n60289, Z => n60287);
   U1688 : BUF_X1 port map( A => n60262, Z => n60259);
   U1689 : BUF_X1 port map( A => n60262, Z => n60260);
   U1690 : BUF_X1 port map( A => n60253, Z => n60250);
   U1691 : BUF_X1 port map( A => n60253, Z => n60251);
   U1692 : BUF_X1 port map( A => n60244, Z => n60241);
   U1693 : BUF_X1 port map( A => n60244, Z => n60242);
   U1694 : BUF_X1 port map( A => n60235, Z => n60232);
   U1695 : BUF_X1 port map( A => n60235, Z => n60233);
   U1696 : BUF_X1 port map( A => n60208, Z => n60205);
   U1697 : BUF_X1 port map( A => n60208, Z => n60206);
   U1698 : BUF_X1 port map( A => n60199, Z => n60196);
   U1699 : BUF_X1 port map( A => n60199, Z => n60197);
   U1700 : BUF_X1 port map( A => n60190, Z => n60187);
   U1701 : BUF_X1 port map( A => n60190, Z => n60188);
   U1702 : BUF_X1 port map( A => n60181, Z => n60178);
   U1703 : BUF_X1 port map( A => n60181, Z => n60179);
   U1704 : BUF_X1 port map( A => n60172, Z => n60169);
   U1705 : BUF_X1 port map( A => n60172, Z => n60170);
   U1706 : BUF_X1 port map( A => n60145, Z => n60142);
   U1707 : BUF_X1 port map( A => n60145, Z => n60143);
   U1708 : BUF_X1 port map( A => n60136, Z => n60133);
   U1709 : BUF_X1 port map( A => n60136, Z => n60134);
   U1710 : BUF_X1 port map( A => n60127, Z => n60124);
   U1711 : BUF_X1 port map( A => n60127, Z => n60125);
   U1712 : BUF_X1 port map( A => n60118, Z => n60115);
   U1713 : BUF_X1 port map( A => n60118, Z => n60116);
   U1714 : BUF_X1 port map( A => n60109, Z => n60106);
   U1715 : BUF_X1 port map( A => n60109, Z => n60107);
   U1716 : BUF_X1 port map( A => n60820, Z => n60817);
   U1717 : BUF_X1 port map( A => n60820, Z => n60818);
   U1718 : BUF_X1 port map( A => n60793, Z => n60790);
   U1719 : BUF_X1 port map( A => n60793, Z => n60791);
   U1720 : BUF_X1 port map( A => n60784, Z => n60781);
   U1721 : BUF_X1 port map( A => n60784, Z => n60782);
   U1722 : BUF_X1 port map( A => n60775, Z => n60772);
   U1723 : BUF_X1 port map( A => n60775, Z => n60773);
   U1724 : BUF_X1 port map( A => n60766, Z => n60763);
   U1725 : BUF_X1 port map( A => n60766, Z => n60764);
   U1726 : BUF_X1 port map( A => n60757, Z => n60754);
   U1727 : BUF_X1 port map( A => n60757, Z => n60755);
   U1728 : BUF_X1 port map( A => n60748, Z => n60745);
   U1729 : BUF_X1 port map( A => n60748, Z => n60746);
   U1730 : BUF_X1 port map( A => n60739, Z => n60736);
   U1731 : BUF_X1 port map( A => n60739, Z => n60737);
   U1732 : BUF_X1 port map( A => n60730, Z => n60727);
   U1733 : BUF_X1 port map( A => n60730, Z => n60728);
   U1734 : BUF_X1 port map( A => n60703, Z => n60700);
   U1735 : BUF_X1 port map( A => n60703, Z => n60701);
   U1736 : BUF_X1 port map( A => n60694, Z => n60691);
   U1737 : BUF_X1 port map( A => n60694, Z => n60692);
   U1738 : BUF_X1 port map( A => n5416, Z => n59738);
   U1739 : BUF_X1 port map( A => n5416, Z => n59739);
   U1740 : AND2_X1 port map( A1 => n7849, A2 => n7914, ZN => n5495);
   U1741 : AND2_X1 port map( A1 => n14983, A2 => n15041, ZN => n8088);
   U1742 : BUF_X1 port map( A => n59839, Z => n59838);
   U1743 : BUF_X1 port map( A => n60658, Z => n60657);
   U1744 : BUF_X1 port map( A => n60649, Z => n60648);
   U1745 : BUF_X1 port map( A => n60622, Z => n60621);
   U1746 : BUF_X1 port map( A => n60613, Z => n60612);
   U1747 : BUF_X1 port map( A => n60586, Z => n60585);
   U1748 : BUF_X1 port map( A => n60577, Z => n60576);
   U1749 : BUF_X1 port map( A => n60550, Z => n60549);
   U1750 : BUF_X1 port map( A => n60928, Z => n60927);
   U1751 : BUF_X1 port map( A => n60919, Z => n60918);
   U1752 : BUF_X1 port map( A => n59830, Z => n59829);
   U1753 : BUF_X1 port map( A => n60541, Z => n60540);
   U1754 : BUF_X1 port map( A => n60487, Z => n60486);
   U1755 : BUF_X1 port map( A => n60469, Z => n60468);
   U1756 : BUF_X1 port map( A => n60460, Z => n60459);
   U1757 : BUF_X1 port map( A => n60415, Z => n60414);
   U1758 : BUF_X1 port map( A => n60406, Z => n60405);
   U1759 : BUF_X1 port map( A => n59992, Z => n59991);
   U1760 : BUF_X1 port map( A => n59983, Z => n59982);
   U1761 : BUF_X1 port map( A => n59974, Z => n59973);
   U1762 : BUF_X1 port map( A => n59965, Z => n59964);
   U1763 : BUF_X1 port map( A => n59956, Z => n59955);
   U1764 : BUF_X1 port map( A => n59947, Z => n59946);
   U1765 : BUF_X1 port map( A => n59938, Z => n59937);
   U1766 : BUF_X1 port map( A => n59920, Z => n59919);
   U1767 : BUF_X1 port map( A => n59911, Z => n59910);
   U1768 : BUF_X1 port map( A => n59902, Z => n59901);
   U1769 : BUF_X1 port map( A => n59893, Z => n59892);
   U1770 : BUF_X1 port map( A => n59884, Z => n59883);
   U1771 : BUF_X1 port map( A => n59875, Z => n59874);
   U1772 : BUF_X1 port map( A => n59857, Z => n59856);
   U1773 : BUF_X1 port map( A => n59848, Z => n59847);
   U1774 : BUF_X1 port map( A => n59821, Z => n59820);
   U1775 : BUF_X1 port map( A => n60676, Z => n60675);
   U1776 : BUF_X1 port map( A => n60667, Z => n60666);
   U1777 : BUF_X1 port map( A => n60640, Z => n60639);
   U1778 : BUF_X1 port map( A => n60631, Z => n60630);
   U1779 : BUF_X1 port map( A => n60604, Z => n60603);
   U1780 : BUF_X1 port map( A => n60595, Z => n60594);
   U1781 : BUF_X1 port map( A => n60568, Z => n60567);
   U1782 : BUF_X1 port map( A => n60559, Z => n60558);
   U1783 : BUF_X1 port map( A => n60532, Z => n60531);
   U1784 : BUF_X1 port map( A => n60523, Z => n60522);
   U1785 : BUF_X1 port map( A => n60514, Z => n60513);
   U1786 : BUF_X1 port map( A => n60505, Z => n60504);
   U1787 : BUF_X1 port map( A => n60496, Z => n60495);
   U1788 : BUF_X1 port map( A => n60478, Z => n60477);
   U1789 : BUF_X1 port map( A => n60451, Z => n60450);
   U1790 : BUF_X1 port map( A => n60442, Z => n60441);
   U1791 : BUF_X1 port map( A => n60433, Z => n60432);
   U1792 : BUF_X1 port map( A => n60424, Z => n60423);
   U1793 : BUF_X1 port map( A => n60397, Z => n60396);
   U1794 : BUF_X1 port map( A => n60127, Z => n60126);
   U1795 : BUF_X1 port map( A => n60118, Z => n60117);
   U1796 : BUF_X1 port map( A => n60109, Z => n60108);
   U1797 : BUF_X1 port map( A => n60892, Z => n60891);
   U1798 : BUF_X1 port map( A => n60883, Z => n60882);
   U1799 : BUF_X1 port map( A => n60856, Z => n60855);
   U1800 : BUF_X1 port map( A => n60847, Z => n60846);
   U1801 : BUF_X1 port map( A => n60838, Z => n60837);
   U1802 : BUF_X1 port map( A => n60829, Z => n60828);
   U1803 : BUF_X1 port map( A => n60811, Z => n60810);
   U1804 : BUF_X1 port map( A => n60802, Z => n60801);
   U1805 : BUF_X1 port map( A => n60712, Z => n60711);
   U1806 : BUF_X1 port map( A => n59929, Z => n59928);
   U1807 : BUF_X1 port map( A => n59866, Z => n59865);
   U1808 : BUF_X1 port map( A => n60946, Z => n60945);
   U1809 : BUF_X1 port map( A => n60937, Z => n60936);
   U1810 : BUF_X1 port map( A => n60379, Z => n60378);
   U1811 : BUF_X1 port map( A => n60370, Z => n60369);
   U1812 : BUF_X1 port map( A => n60361, Z => n60360);
   U1813 : BUF_X1 port map( A => n60352, Z => n60351);
   U1814 : BUF_X1 port map( A => n60343, Z => n60342);
   U1815 : BUF_X1 port map( A => n60280, Z => n60279);
   U1816 : BUF_X1 port map( A => n60271, Z => n60270);
   U1817 : BUF_X1 port map( A => n60226, Z => n60225);
   U1818 : BUF_X1 port map( A => n60217, Z => n60216);
   U1819 : BUF_X1 port map( A => n60163, Z => n60162);
   U1820 : BUF_X1 port map( A => n60154, Z => n60153);
   U1821 : BUF_X1 port map( A => n60721, Z => n60720);
   U1822 : BUF_X1 port map( A => n60685, Z => n60684);
   U1823 : BUF_X1 port map( A => n60100, Z => n60099);
   U1824 : BUF_X1 port map( A => n60091, Z => n60090);
   U1825 : BUF_X1 port map( A => n60082, Z => n60081);
   U1826 : BUF_X1 port map( A => n60073, Z => n60072);
   U1827 : BUF_X1 port map( A => n60064, Z => n60063);
   U1828 : BUF_X1 port map( A => n60055, Z => n60054);
   U1829 : BUF_X1 port map( A => n60046, Z => n60045);
   U1830 : BUF_X1 port map( A => n60037, Z => n60036);
   U1831 : BUF_X1 port map( A => n60028, Z => n60027);
   U1832 : BUF_X1 port map( A => n60019, Z => n60018);
   U1833 : BUF_X1 port map( A => n60010, Z => n60009);
   U1834 : BUF_X1 port map( A => n60001, Z => n60000);
   U1835 : BUF_X1 port map( A => n61244, Z => n61243);
   U1836 : BUF_X1 port map( A => n60955, Z => n60954);
   U1837 : BUF_X1 port map( A => n60910, Z => n60909);
   U1838 : BUF_X1 port map( A => n60325, Z => n60324);
   U1839 : BUF_X1 port map( A => n60316, Z => n60315);
   U1840 : BUF_X1 port map( A => n60307, Z => n60306);
   U1841 : BUF_X1 port map( A => n60298, Z => n60297);
   U1842 : BUF_X1 port map( A => n60289, Z => n60288);
   U1843 : BUF_X1 port map( A => n60262, Z => n60261);
   U1844 : BUF_X1 port map( A => n60253, Z => n60252);
   U1845 : BUF_X1 port map( A => n60244, Z => n60243);
   U1846 : BUF_X1 port map( A => n60235, Z => n60234);
   U1847 : BUF_X1 port map( A => n60208, Z => n60207);
   U1848 : BUF_X1 port map( A => n60199, Z => n60198);
   U1849 : BUF_X1 port map( A => n60190, Z => n60189);
   U1850 : BUF_X1 port map( A => n60181, Z => n60180);
   U1851 : BUF_X1 port map( A => n60172, Z => n60171);
   U1852 : BUF_X1 port map( A => n60145, Z => n60144);
   U1853 : BUF_X1 port map( A => n60136, Z => n60135);
   U1854 : BUF_X1 port map( A => n60874, Z => n60873);
   U1855 : BUF_X1 port map( A => n60865, Z => n60864);
   U1856 : BUF_X1 port map( A => n60901, Z => n60900);
   U1857 : BUF_X1 port map( A => n60388, Z => n60387);
   U1858 : BUF_X1 port map( A => n60334, Z => n60333);
   U1859 : BUF_X1 port map( A => n60820, Z => n60819);
   U1860 : BUF_X1 port map( A => n60793, Z => n60792);
   U1861 : BUF_X1 port map( A => n60784, Z => n60783);
   U1862 : BUF_X1 port map( A => n60775, Z => n60774);
   U1863 : BUF_X1 port map( A => n60766, Z => n60765);
   U1864 : BUF_X1 port map( A => n60757, Z => n60756);
   U1865 : BUF_X1 port map( A => n60748, Z => n60747);
   U1866 : BUF_X1 port map( A => n60739, Z => n60738);
   U1867 : BUF_X1 port map( A => n60730, Z => n60729);
   U1868 : BUF_X1 port map( A => n60703, Z => n60702);
   U1869 : BUF_X1 port map( A => n60694, Z => n60693);
   U1870 : AND2_X1 port map( A1 => n7870, A2 => n7849, ZN => n5451);
   U1871 : AND2_X1 port map( A1 => n7855, A2 => n7849, ZN => n5443);
   U1872 : AND2_X1 port map( A1 => n7853, A2 => n7849, ZN => n5414);
   U1873 : AND2_X1 port map( A1 => n7861, A2 => n7849, ZN => n5400);
   U1874 : AND2_X1 port map( A1 => n7848, A2 => n7849, ZN => n5525);
   U1875 : AND2_X1 port map( A1 => n7912, A2 => n7849, ZN => n5487);
   U1876 : AND2_X1 port map( A1 => n7886, A2 => n7849, ZN => n5478);
   U1877 : AND2_X1 port map( A1 => n7896, A2 => n7849, ZN => n5548);
   U1878 : AND2_X1 port map( A1 => n7924, A2 => n7849, ZN => n5520);
   U1879 : AND2_X1 port map( A1 => n15004, A2 => n14983, ZN => n8014);
   U1880 : AND2_X1 port map( A1 => n15000, A2 => n14983, ZN => n8000);
   U1881 : AND2_X1 port map( A1 => n14992, A2 => n14983, ZN => n7989);
   U1882 : AND2_X1 port map( A1 => n15016, A2 => n14983, ZN => n8039);
   U1883 : AND2_X1 port map( A1 => n14990, A2 => n14983, ZN => n7974);
   U1884 : AND2_X1 port map( A1 => n14977, A2 => n14983, ZN => n7964);
   U1885 : AND2_X1 port map( A1 => n15050, A2 => n14983, ZN => n8113);
   U1886 : AND2_X1 port map( A1 => n15058, A2 => n14983, ZN => n8123);
   U1887 : AND2_X1 port map( A1 => n15047, A2 => n14983, ZN => n8098);
   U1888 : AND2_X1 port map( A1 => n15068, A2 => n14983, ZN => n8148);
   U1889 : AND2_X1 port map( A1 => n15026, A2 => n14983, ZN => n8062);
   U1890 : AND2_X1 port map( A1 => n15038, A2 => n14983, ZN => n8072);
   U1891 : BUF_X1 port map( A => n5419, Z => n59740);
   U1892 : BUF_X1 port map( A => n5419, Z => n59741);
   U1893 : BUF_X1 port map( A => n5415, Z => n59744);
   U1894 : BUF_X1 port map( A => n5415, Z => n59745);
   U1895 : BUF_X1 port map( A => n59758, Z => n59757);
   U1896 : BUF_X1 port map( A => n59758, Z => n59749);
   U1897 : BUF_X1 port map( A => n59758, Z => n59750);
   U1898 : BUF_X1 port map( A => n59758, Z => n59751);
   U1899 : BUF_X1 port map( A => n59758, Z => n59752);
   U1900 : BUF_X1 port map( A => n59758, Z => n59753);
   U1901 : BUF_X1 port map( A => n59758, Z => n59754);
   U1902 : BUF_X1 port map( A => n59749, Z => n59755);
   U1903 : BUF_X1 port map( A => n59750, Z => n59756);
   U1904 : BUF_X1 port map( A => n5419, Z => n59742);
   U1905 : BUF_X1 port map( A => n5419, Z => n59743);
   U1906 : BUF_X1 port map( A => n5415, Z => n59746);
   U1907 : BUF_X1 port map( A => n5415, Z => n59747);
   U1908 : NAND2_X1 port map( A1 => n7862, A2 => n7914, ZN => n5484);
   U1909 : NAND2_X1 port map( A1 => n7852, A2 => n7914, ZN => n5493);
   U1910 : NAND2_X1 port map( A1 => n7860, A2 => n7914, ZN => n5492);
   U1911 : NAND2_X1 port map( A1 => n7850, A2 => n7912, ZN => n5485);
   U1912 : NAND2_X1 port map( A1 => n7920, A2 => n7862, ZN => n5500);
   U1913 : NAND2_X1 port map( A1 => n7875, A2 => n7852, ZN => n5456);
   U1914 : NAND2_X1 port map( A1 => n7934, A2 => n7852, ZN => n5536);
   U1915 : NAND2_X1 port map( A1 => n7857, A2 => n7856, ZN => n5397);
   U1916 : NAND2_X1 port map( A1 => n7855, A2 => n7856, ZN => n5386);
   U1917 : NAND2_X1 port map( A1 => n7855, A2 => n7860, ZN => n5435);
   U1918 : NAND2_X1 port map( A1 => n7924, A2 => n7860, ZN => n5503);
   U1919 : NAND2_X1 port map( A1 => n7870, A2 => n7864, ZN => n5440);
   U1920 : NAND2_X1 port map( A1 => n7883, A2 => n7859, ZN => n5459);
   U1921 : NAND2_X1 port map( A1 => n7848, A2 => n7859, ZN => n5516);
   U1922 : NOR2_X1 port map( A1 => ADDR_WR(6), A2 => ADDR_WR(5), ZN => n15127);
   U1923 : NAND2_X1 port map( A1 => n7896, A2 => n7850, ZN => n5449);
   U1924 : NAND2_X1 port map( A1 => n7855, A2 => n7850, ZN => n5441);
   U1925 : NAND2_X1 port map( A1 => n7886, A2 => n7859, ZN => n5460);
   U1926 : NAND2_X1 port map( A1 => n7896, A2 => n7864, ZN => n5448);
   U1927 : NOR2_X1 port map( A1 => n5282, A2 => n5283, ZN => n15263);
   U1928 : NAND2_X1 port map( A1 => n7848, A2 => n7860, ZN => n5517);
   U1929 : NAND2_X1 port map( A1 => n7920, A2 => n7860, ZN => n5501);
   U1930 : NAND2_X1 port map( A1 => n7875, A2 => n7850, ZN => n5453);
   U1931 : NAND2_X1 port map( A1 => n15261, A2 => n15284, ZN => n15107);
   U1932 : NAND2_X1 port map( A1 => n15259, A2 => n15279, ZN => n15097);
   U1933 : NAND2_X1 port map( A1 => n15261, A2 => n15279, ZN => n15099);
   U1934 : NAND2_X1 port map( A1 => n15279, A2 => n15263, ZN => n15101);
   U1935 : NAND2_X1 port map( A1 => n15257, A2 => n15284, ZN => n15103);
   U1936 : NAND2_X1 port map( A1 => n15259, A2 => n15284, ZN => n15105);
   U1937 : NAND2_X1 port map( A1 => n15279, A2 => n15257, ZN => n15095);
   U1938 : NAND2_X1 port map( A1 => n7875, A2 => n7864, ZN => n5454);
   U1939 : NAND2_X1 port map( A1 => n7920, A2 => n7864, ZN => n5504);
   U1940 : NOR2_X1 port map( A1 => n5281, A2 => ADDR_WR(3), ZN => n15284);
   U1941 : NAND2_X1 port map( A1 => n7855, A2 => n7859, ZN => n5436);
   U1942 : NAND2_X1 port map( A1 => n7875, A2 => n7859, ZN => n5457);
   U1943 : NAND2_X1 port map( A1 => n7934, A2 => n7850, ZN => n5537);
   U1944 : NAND2_X1 port map( A1 => n7861, A2 => n7850, ZN => n5398);
   U1945 : NAND2_X1 port map( A1 => n15265, A2 => n15263, ZN => n15125);
   U1946 : NAND2_X1 port map( A1 => n15256, A2 => n15259, ZN => n15113);
   U1947 : NAND2_X1 port map( A1 => n15265, A2 => n15259, ZN => n15121);
   U1948 : NAND2_X1 port map( A1 => n15265, A2 => n15257, ZN => n15119);
   U1949 : NAND2_X1 port map( A1 => n15256, A2 => n15257, ZN => n15111);
   U1950 : NAND2_X1 port map( A1 => n15256, A2 => n15261, ZN => n15115);
   U1951 : NAND2_X1 port map( A1 => n15265, A2 => n15261, ZN => n15123);
   U1952 : AND3_X1 port map( A1 => n7890, A2 => n5287, A3 => n7872, ZN => n7861
                           );
   U1953 : INV_X1 port map( A => ADDR_RD1(7), ZN => n5287);
   U1954 : NAND2_X1 port map( A1 => n7862, A2 => n7912, ZN => n5474);
   U1955 : NAND2_X1 port map( A1 => n7851, A2 => n7862, ZN => n5415);
   U1956 : NAND2_X1 port map( A1 => n7852, A2 => n7912, ZN => n5480);
   U1957 : NAND2_X1 port map( A1 => n14981, A2 => n15041, ZN => n8075);
   U1958 : NAND2_X1 port map( A1 => n7853, A2 => n7864, ZN => n5419);
   U1959 : NAND2_X1 port map( A1 => n7864, A2 => n7914, ZN => n5497);
   U1960 : NAND2_X1 port map( A1 => n7864, A2 => n7912, ZN => n5479);
   U1961 : NAND2_X1 port map( A1 => n14986, A2 => n15041, ZN => n8084);
   U1962 : NAND2_X1 port map( A1 => n14986, A2 => n15038, ZN => n8070);
   U1963 : NAND2_X1 port map( A1 => n7850, A2 => n7914, ZN => n5498);
   U1964 : NAND2_X1 port map( A1 => n14980, A2 => n15041, ZN => n8074);
   U1965 : AND3_X1 port map( A1 => n14987, A2 => n5354, A3 => n14988, ZN => 
                           n14977);
   U1966 : INV_X1 port map( A => ADDR_RD2(7), ZN => n5354);
   U1967 : NAND2_X1 port map( A1 => n7851, A2 => n7860, ZN => n5416);
   U1968 : NAND2_X1 port map( A1 => n14984, A2 => n15041, ZN => n8085);
   U1969 : NAND2_X1 port map( A1 => n7857, A2 => n7862, ZN => n6025);
   U1970 : NAND2_X1 port map( A1 => n7853, A2 => n7862, ZN => n6033);
   U1971 : NAND2_X1 port map( A1 => n7861, A2 => n7862, ZN => n6021);
   U1972 : NAND2_X1 port map( A1 => n7924, A2 => n7862, ZN => n6092);
   U1973 : NAND2_X1 port map( A1 => n7855, A2 => n7852, ZN => n6044);
   U1974 : NAND2_X1 port map( A1 => n7870, A2 => n7852, ZN => n6048);
   U1975 : NAND2_X1 port map( A1 => n7920, A2 => n7852, ZN => n6086);
   U1976 : NOR2_X1 port map( A1 => n5349, A2 => ADDR_RD1(3), ZN => n7877);
   U1977 : NOR2_X1 port map( A1 => n5357, A2 => ADDR_RD2(3), ZN => n15001);
   U1978 : NAND2_X1 port map( A1 => n7924, A2 => n7856, ZN => n6089);
   U1979 : NAND2_X1 port map( A1 => n7914, A2 => n7856, ZN => n6078);
   U1980 : NAND2_X1 port map( A1 => n7896, A2 => n7856, ZN => n6107);
   U1981 : NAND2_X1 port map( A1 => n7870, A2 => n7862, ZN => n5432);
   U1982 : NAND2_X1 port map( A1 => n7886, A2 => n7862, ZN => n5428);
   U1983 : NAND2_X1 port map( A1 => n7875, A2 => n7862, ZN => n5410);
   U1984 : NAND2_X1 port map( A1 => n7896, A2 => n7862, ZN => n5539);
   U1985 : NAND2_X1 port map( A1 => ADDR_RD1(7), A2 => n7862, ZN => n5544);
   U1986 : NAND2_X1 port map( A1 => n7934, A2 => n7862, ZN => n5527);
   U1987 : NAND2_X1 port map( A1 => n7848, A2 => n7862, ZN => n5511);
   U1988 : NOR2_X1 port map( A1 => n5358, A2 => ADDR_RD2(4), ZN => n14993);
   U1989 : NOR2_X1 port map( A1 => n5350, A2 => ADDR_RD1(4), ZN => n7873);
   U1990 : NOR2_X1 port map( A1 => n5347, A2 => ADDR_RD1(5), ZN => n7910);
   U1991 : NOR2_X1 port map( A1 => n5355, A2 => ADDR_RD2(5), ZN => n15036);
   U1992 : NAND2_X1 port map( A1 => n7883, A2 => n7860, ZN => n6056);
   U1993 : NAND2_X1 port map( A1 => n7875, A2 => n7860, ZN => n6047);
   U1994 : NAND2_X1 port map( A1 => n7853, A2 => n7860, ZN => n6034);
   U1995 : NOR2_X1 port map( A1 => ADDR_RD2(3), A2 => ADDR_RD2(4), ZN => n14987
                           );
   U1996 : NOR2_X1 port map( A1 => ADDR_RD1(3), A2 => ADDR_RD1(4), ZN => n7890)
                           ;
   U1997 : NAND2_X1 port map( A1 => n7853, A2 => n7852, ZN => n5405);
   U1998 : NAND2_X1 port map( A1 => n7861, A2 => n7852, ZN => n5390);
   U1999 : NAND2_X1 port map( A1 => n7851, A2 => n7852, ZN => n5418);
   U2000 : NAND2_X1 port map( A1 => ADDR_RD1(7), A2 => n7852, ZN => n5550);
   U2001 : NAND2_X1 port map( A1 => n7848, A2 => n7852, ZN => n5522);
   U2002 : NOR2_X1 port map( A1 => ADDR_RD1(5), A2 => ADDR_RD1(6), ZN => n7872)
                           ;
   U2003 : NOR2_X1 port map( A1 => ADDR_RD2(5), A2 => ADDR_RD2(6), ZN => n14988
                           );
   U2004 : NOR2_X1 port map( A1 => n5348, A2 => ADDR_RD1(6), ZN => n7889);
   U2005 : NOR2_X1 port map( A1 => n5356, A2 => ADDR_RD2(6), ZN => n15012);
   U2006 : NAND2_X1 port map( A1 => n7886, A2 => n7864, ZN => n6073);
   U2007 : INV_X1 port map( A => ADDR_WR(6), ZN => n5278);
   U2008 : NAND2_X1 port map( A1 => n7870, A2 => n7856, ZN => n5433);
   U2009 : NAND2_X1 port map( A1 => n7875, A2 => n7856, ZN => n5411);
   U2010 : NAND2_X1 port map( A1 => n7886, A2 => n7856, ZN => n5471);
   U2011 : NAND2_X1 port map( A1 => n7912, A2 => n7856, ZN => n5475);
   U2012 : NAND2_X1 port map( A1 => n7934, A2 => n7856, ZN => n5526);
   U2013 : NAND2_X1 port map( A1 => n7848, A2 => n7856, ZN => n5512);
   U2014 : NAND2_X1 port map( A1 => n15013, A2 => n14981, ZN => n8010);
   U2015 : NAND2_X1 port map( A1 => n14992, A2 => n14981, ZN => n7981);
   U2016 : NAND2_X1 port map( A1 => n15000, A2 => n14981, ZN => n7990);
   U2017 : NAND2_X1 port map( A1 => n15023, A2 => n14981, ZN => n8035);
   U2018 : NAND2_X1 port map( A1 => n14977, A2 => n14981, ZN => n7955);
   U2019 : NAND2_X1 port map( A1 => n14990, A2 => n14981, ZN => n7965);
   U2020 : NAND2_X1 port map( A1 => n15058, A2 => n14981, ZN => n8109);
   U2021 : NAND2_X1 port map( A1 => n15061, A2 => n14981, ZN => n8119);
   U2022 : NAND2_X1 port map( A1 => n15050, A2 => n14981, ZN => n8099);
   U2023 : NAND2_X1 port map( A1 => n15047, A2 => n14981, ZN => n8090);
   U2024 : NAND2_X1 port map( A1 => ADDR_RD2(7), A2 => n14981, ZN => n8144);
   U2025 : NAND2_X1 port map( A1 => n15038, A2 => n14981, ZN => n8064);
   U2026 : NAND2_X1 port map( A1 => n7886, A2 => n7860, ZN => n5427);
   U2027 : NAND2_X1 port map( A1 => n7861, A2 => n7860, ZN => n5392);
   U2028 : NAND2_X1 port map( A1 => n7896, A2 => n7860, ZN => n5540);
   U2029 : NAND2_X1 port map( A1 => ADDR_RD1(7), A2 => n7860, ZN => n5545);
   U2030 : NAND2_X1 port map( A1 => n7883, A2 => n7850, ZN => n6059);
   U2031 : NAND2_X1 port map( A1 => n7857, A2 => n7850, ZN => n6018);
   U2032 : INV_X1 port map( A => ADDR_WR(5), ZN => n5279);
   U2033 : NAND2_X1 port map( A1 => n7861, A2 => n7864, ZN => n5389);
   U2034 : NAND2_X1 port map( A1 => n7848, A2 => n7864, ZN => n5521);
   U2035 : NAND2_X1 port map( A1 => n15004, A2 => n14985, ZN => n8006);
   U2036 : NAND2_X1 port map( A1 => n15013, A2 => n14985, ZN => n8016);
   U2037 : NAND2_X1 port map( A1 => n15016, A2 => n14985, ZN => n8031);
   U2038 : NAND2_X1 port map( A1 => n15023, A2 => n14985, ZN => n8041);
   U2039 : NAND2_X1 port map( A1 => n14990, A2 => n14985, ZN => n7970);
   U2040 : NAND2_X1 port map( A1 => n14977, A2 => n14985, ZN => n7961);
   U2041 : NAND2_X1 port map( A1 => n15058, A2 => n14985, ZN => n8115);
   U2042 : NAND2_X1 port map( A1 => n15068, A2 => n14985, ZN => n8140);
   U2043 : NAND2_X1 port map( A1 => ADDR_RD2(7), A2 => n14985, ZN => n8150);
   U2044 : NAND2_X1 port map( A1 => n15026, A2 => n14985, ZN => n8059);
   U2045 : NAND2_X1 port map( A1 => n15038, A2 => n14985, ZN => n8069);
   U2046 : NAND2_X1 port map( A1 => n15004, A2 => n14986, ZN => n8005);
   U2047 : NAND2_X1 port map( A1 => n15013, A2 => n14986, ZN => n8015);
   U2048 : NAND2_X1 port map( A1 => n15000, A2 => n14986, ZN => n7995);
   U2049 : NAND2_X1 port map( A1 => n14992, A2 => n14986, ZN => n7985);
   U2050 : NAND2_X1 port map( A1 => n14990, A2 => n14986, ZN => n7971);
   U2051 : NAND2_X1 port map( A1 => n14977, A2 => n14986, ZN => n7960);
   U2052 : NAND2_X1 port map( A1 => n15058, A2 => n14986, ZN => n8114);
   U2053 : NAND2_X1 port map( A1 => n15047, A2 => n14986, ZN => n8094);
   U2054 : NAND2_X1 port map( A1 => n15026, A2 => n14986, ZN => n8060);
   U2055 : NAND2_X1 port map( A1 => n7861, A2 => n7859, ZN => n5393);
   U2056 : NAND2_X1 port map( A1 => n7853, A2 => n7859, ZN => n5406);
   U2057 : NAND2_X1 port map( A1 => ADDR_RD1(7), A2 => n7859, ZN => n5549);
   U2058 : NAND2_X1 port map( A1 => n15013, A2 => n14980, ZN => n8011);
   U2059 : NAND2_X1 port map( A1 => n15026, A2 => n14980, ZN => n8046);
   U2060 : NAND2_X1 port map( A1 => n14977, A2 => n14980, ZN => n7956);
   U2061 : NAND2_X1 port map( A1 => n14990, A2 => n14980, ZN => n7966);
   U2062 : NAND2_X1 port map( A1 => n15058, A2 => n14980, ZN => n8110);
   U2063 : NAND2_X1 port map( A1 => n15061, A2 => n14980, ZN => n8120);
   U2064 : NAND2_X1 port map( A1 => n15068, A2 => n14980, ZN => n8135);
   U2065 : NAND2_X1 port map( A1 => n15038, A2 => n14980, ZN => n8065);
   U2066 : NAND2_X1 port map( A1 => n14992, A2 => n14979, ZN => n7980);
   U2067 : NAND2_X1 port map( A1 => n15000, A2 => n14979, ZN => n7991);
   U2068 : NAND2_X1 port map( A1 => n15023, A2 => n14979, ZN => n8036);
   U2069 : NAND2_X1 port map( A1 => n15061, A2 => n14979, ZN => n8124);
   U2070 : NAND2_X1 port map( A1 => n15050, A2 => n14979, ZN => n8100);
   U2071 : NAND2_X1 port map( A1 => n15047, A2 => n14979, ZN => n8089);
   U2072 : NAND2_X1 port map( A1 => ADDR_RD2(7), A2 => n14979, ZN => n8145);
   U2073 : NAND2_X1 port map( A1 => n15016, A2 => n14978, ZN => n8030);
   U2074 : NAND2_X1 port map( A1 => n15023, A2 => n14978, ZN => n8040);
   U2075 : NAND2_X1 port map( A1 => n15061, A2 => n14978, ZN => n8125);
   U2076 : NAND2_X1 port map( A1 => n15068, A2 => n14978, ZN => n8139);
   U2077 : NAND2_X1 port map( A1 => ADDR_RD2(7), A2 => n14978, ZN => n8149);
   U2078 : NAND2_X1 port map( A1 => n15013, A2 => n14984, ZN => n8020);
   U2079 : NAND2_X1 port map( A1 => n15000, A2 => n14984, ZN => n7996);
   U2080 : NAND2_X1 port map( A1 => n14992, A2 => n14984, ZN => n7986);
   U2081 : NAND2_X1 port map( A1 => n15047, A2 => n14984, ZN => n8095);
   U2082 : AND2_X1 port map( A1 => ADDR_WR(3), A2 => n5281, ZN => n15256);
   U2083 : BUF_X1 port map( A => n5362, Z => n62120);
   U2084 : BUF_X1 port map( A => n5362, Z => n62119);
   U2085 : BUF_X1 port map( A => n5362, Z => n62122);
   U2086 : BUF_X1 port map( A => n5362, Z => n62121);
   U2087 : BUF_X1 port map( A => n5362, Z => n62124);
   U2088 : BUF_X1 port map( A => n5362, Z => n62123);
   U2089 : AND2_X1 port map( A1 => n7860, A2 => n7912, ZN => n5482);
   U2090 : AND2_X1 port map( A1 => n14985, A2 => n15041, ZN => n8077);
   U2091 : BUF_X1 port map( A => n59812, Z => n59810);
   U2092 : BUF_X1 port map( A => n59812, Z => n59805);
   U2093 : BUF_X1 port map( A => n59812, Z => n59806);
   U2094 : BUF_X1 port map( A => n59812, Z => n59807);
   U2095 : BUF_X1 port map( A => n59812, Z => n59808);
   U2096 : BUF_X1 port map( A => n59812, Z => n59809);
   U2097 : BUF_X1 port map( A => n59803, Z => n59796);
   U2098 : BUF_X1 port map( A => n59803, Z => n59797);
   U2099 : BUF_X1 port map( A => n59803, Z => n59798);
   U2100 : BUF_X1 port map( A => n59803, Z => n59799);
   U2101 : BUF_X1 port map( A => n59794, Z => n59787);
   U2102 : BUF_X1 port map( A => n59794, Z => n59788);
   U2103 : BUF_X1 port map( A => n59794, Z => n59789);
   U2104 : BUF_X1 port map( A => n59794, Z => n59790);
   U2105 : BUF_X1 port map( A => n59785, Z => n59781);
   U2106 : BUF_X1 port map( A => n59776, Z => n59769);
   U2107 : BUF_X1 port map( A => n59776, Z => n59770);
   U2108 : BUF_X1 port map( A => n59785, Z => n59778);
   U2109 : BUF_X1 port map( A => n59785, Z => n59779);
   U2110 : BUF_X1 port map( A => n59785, Z => n59780);
   U2111 : BUF_X1 port map( A => n59776, Z => n59771);
   U2112 : BUF_X1 port map( A => n59776, Z => n59772);
   U2113 : BUF_X1 port map( A => n59767, Z => n59760);
   U2114 : BUF_X1 port map( A => n59767, Z => n59761);
   U2115 : BUF_X1 port map( A => n59767, Z => n59762);
   U2116 : BUF_X1 port map( A => n59767, Z => n59763);
   U2117 : BUF_X1 port map( A => n59767, Z => n59764);
   U2118 : BUF_X1 port map( A => n59803, Z => n59800);
   U2119 : BUF_X1 port map( A => n59803, Z => n59801);
   U2120 : BUF_X1 port map( A => n59794, Z => n59791);
   U2121 : BUF_X1 port map( A => n59794, Z => n59792);
   U2122 : BUF_X1 port map( A => n59785, Z => n59782);
   U2123 : BUF_X1 port map( A => n59785, Z => n59783);
   U2124 : BUF_X1 port map( A => n59776, Z => n59773);
   U2125 : BUF_X1 port map( A => n59776, Z => n59774);
   U2126 : BUF_X1 port map( A => n59767, Z => n59765);
   U2127 : BUF_X1 port map( A => n5362, Z => n62125);
   U2128 : AND2_X1 port map( A1 => n14979, A2 => n15041, ZN => n8079);
   U2129 : AND2_X1 port map( A1 => n7855, A2 => n7862, ZN => n5422);
   U2130 : AND2_X1 port map( A1 => n7857, A2 => n7852, ZN => n5409);
   U2131 : AND2_X1 port map( A1 => n7896, A2 => n7852, ZN => n5542);
   U2132 : AND2_X1 port map( A1 => n14984, A2 => n15038, ZN => n8073);
   U2133 : AND2_X1 port map( A1 => n7883, A2 => n7856, ZN => n5462);
   U2134 : AND2_X1 port map( A1 => n7851, A2 => n7856, ZN => n5413);
   U2135 : AND2_X1 port map( A1 => n7920, A2 => n7856, ZN => n5496);
   U2136 : AND2_X1 port map( A1 => ADDR_RD1(7), A2 => n7856, ZN => n5547);
   U2137 : AND2_X1 port map( A1 => n15016, A2 => n14981, ZN => n8024);
   U2138 : AND2_X1 port map( A1 => n15004, A2 => n14981, ZN => n7998);
   U2139 : AND2_X1 port map( A1 => n15026, A2 => n14981, ZN => n8050);
   U2140 : AND2_X1 port map( A1 => n15068, A2 => n14981, ZN => n8138);
   U2141 : AND2_X1 port map( A1 => n7870, A2 => n7860, ZN => n5438);
   U2142 : AND2_X1 port map( A1 => n7857, A2 => n7860, ZN => n5395);
   U2143 : AND2_X1 port map( A1 => n7934, A2 => n7860, ZN => n5530);
   U2144 : AND2_X1 port map( A1 => n7851, A2 => n7864, ZN => n5431);
   U2145 : AND2_X1 port map( A1 => n7857, A2 => n7864, ZN => n5408);
   U2146 : AND2_X1 port map( A1 => ADDR_RD1(7), A2 => n7864, ZN => n5554);
   U2147 : AND2_X1 port map( A1 => n7934, A2 => n7864, ZN => n5531);
   U2148 : AND2_X1 port map( A1 => n7924, A2 => n7864, ZN => n5514);
   U2149 : AND2_X1 port map( A1 => n14992, A2 => n14985, ZN => n7984);
   U2150 : AND2_X1 port map( A1 => n15000, A2 => n14985, ZN => n7993);
   U2151 : AND2_X1 port map( A1 => n15061, A2 => n14985, ZN => n8129);
   U2152 : AND2_X1 port map( A1 => n15050, A2 => n14985, ZN => n8103);
   U2153 : AND2_X1 port map( A1 => n15047, A2 => n14985, ZN => n8093);
   U2154 : AND2_X1 port map( A1 => n15016, A2 => n14986, ZN => n8034);
   U2155 : AND2_X1 port map( A1 => n15023, A2 => n14986, ZN => n8044);
   U2156 : AND2_X1 port map( A1 => n15061, A2 => n14986, ZN => n8128);
   U2157 : AND2_X1 port map( A1 => n15050, A2 => n14986, ZN => n8102);
   U2158 : AND2_X1 port map( A1 => n15068, A2 => n14986, ZN => n8143);
   U2159 : AND2_X1 port map( A1 => ADDR_RD2(7), A2 => n14986, ZN => n8154);
   U2160 : AND2_X1 port map( A1 => n7851, A2 => n7859, ZN => n5421);
   U2161 : AND2_X1 port map( A1 => n7870, A2 => n7859, ZN => n5439);
   U2162 : AND2_X1 port map( A1 => n7857, A2 => n7859, ZN => n5396);
   U2163 : AND2_X1 port map( A1 => n7912, A2 => n7859, ZN => n5483);
   U2164 : AND2_X1 port map( A1 => n7896, A2 => n7859, ZN => n5543);
   U2165 : AND2_X1 port map( A1 => n7934, A2 => n7859, ZN => n5529);
   U2166 : AND2_X1 port map( A1 => n7924, A2 => n7859, ZN => n5515);
   U2167 : AND2_X1 port map( A1 => n7851, A2 => n7850, ZN => n5430);
   U2168 : AND2_X1 port map( A1 => n7870, A2 => n7850, ZN => n5452);
   U2169 : AND2_X1 port map( A1 => n7848, A2 => n7850, ZN => n5524);
   U2170 : AND2_X1 port map( A1 => n7920, A2 => n7850, ZN => n5506);
   U2171 : AND2_X1 port map( A1 => n7886, A2 => n7850, ZN => n5477);
   U2172 : AND2_X1 port map( A1 => ADDR_RD1(7), A2 => n7850, ZN => n5553);
   U2173 : AND2_X1 port map( A1 => n7924, A2 => n7850, ZN => n5519);
   U2174 : BUF_X1 port map( A => n59812, Z => n59811);
   U2175 : BUF_X1 port map( A => n59803, Z => n59802);
   U2176 : BUF_X1 port map( A => n59794, Z => n59793);
   U2177 : BUF_X1 port map( A => n59785, Z => n59784);
   U2178 : BUF_X1 port map( A => n59776, Z => n59775);
   U2179 : BUF_X1 port map( A => n59767, Z => n59766);
   U2180 : AND2_X1 port map( A1 => n15016, A2 => n14980, ZN => n8025);
   U2181 : AND2_X1 port map( A1 => n15004, A2 => n14980, ZN => n7999);
   U2182 : AND2_X1 port map( A1 => n15000, A2 => n14980, ZN => n7988);
   U2183 : AND2_X1 port map( A1 => n15023, A2 => n14980, ZN => n8038);
   U2184 : AND2_X1 port map( A1 => n14992, A2 => n14980, ZN => n7973);
   U2185 : AND2_X1 port map( A1 => n15050, A2 => n14980, ZN => n8097);
   U2186 : AND2_X1 port map( A1 => n15047, A2 => n14980, ZN => n8087);
   U2187 : AND2_X1 port map( A1 => ADDR_RD2(7), A2 => n14980, ZN => n8147);
   U2188 : AND2_X1 port map( A1 => n15016, A2 => n14979, ZN => n8023);
   U2189 : AND2_X1 port map( A1 => n15004, A2 => n14979, ZN => n8008);
   U2190 : AND2_X1 port map( A1 => n15013, A2 => n14979, ZN => n8018);
   U2191 : AND2_X1 port map( A1 => n15026, A2 => n14979, ZN => n8049);
   U2192 : AND2_X1 port map( A1 => n14977, A2 => n14979, ZN => n7958);
   U2193 : AND2_X1 port map( A1 => n14990, A2 => n14979, ZN => n7968);
   U2194 : AND2_X1 port map( A1 => n15058, A2 => n14979, ZN => n8117);
   U2195 : AND2_X1 port map( A1 => n15068, A2 => n14979, ZN => n8137);
   U2196 : AND2_X1 port map( A1 => n15038, A2 => n14979, ZN => n8067);
   U2197 : AND2_X1 port map( A1 => ADDR_RD1(7), A2 => n7849, ZN => n5552);
   U2198 : AND2_X1 port map( A1 => n15004, A2 => n14978, ZN => n8009);
   U2199 : AND2_X1 port map( A1 => n15013, A2 => n14978, ZN => n8019);
   U2200 : AND2_X1 port map( A1 => n14992, A2 => n14978, ZN => n7983);
   U2201 : AND2_X1 port map( A1 => n15000, A2 => n14978, ZN => n7994);
   U2202 : AND2_X1 port map( A1 => n15026, A2 => n14978, ZN => n8048);
   U2203 : AND2_X1 port map( A1 => n14977, A2 => n14978, ZN => n7959);
   U2204 : AND2_X1 port map( A1 => n14990, A2 => n14978, ZN => n7969);
   U2205 : AND2_X1 port map( A1 => n15058, A2 => n14978, ZN => n8118);
   U2206 : AND2_X1 port map( A1 => n15050, A2 => n14978, ZN => n8104);
   U2207 : AND2_X1 port map( A1 => n15047, A2 => n14978, ZN => n8092);
   U2208 : AND2_X1 port map( A1 => n15041, A2 => n14978, ZN => n8078);
   U2209 : AND2_X1 port map( A1 => n15038, A2 => n14978, ZN => n8068);
   U2210 : AND2_X1 port map( A1 => n15004, A2 => n14984, ZN => n8013);
   U2211 : AND2_X1 port map( A1 => n15016, A2 => n14984, ZN => n8033);
   U2212 : AND2_X1 port map( A1 => n15023, A2 => n14984, ZN => n8043);
   U2213 : AND2_X1 port map( A1 => n14990, A2 => n14984, ZN => n7975);
   U2214 : AND2_X1 port map( A1 => n14977, A2 => n14984, ZN => n7963);
   U2215 : AND2_X1 port map( A1 => n15061, A2 => n14984, ZN => n8127);
   U2216 : AND2_X1 port map( A1 => n15050, A2 => n14984, ZN => n8112);
   U2217 : AND2_X1 port map( A1 => n15058, A2 => n14984, ZN => n8122);
   U2218 : AND2_X1 port map( A1 => n15068, A2 => n14984, ZN => n8142);
   U2219 : AND2_X1 port map( A1 => ADDR_RD2(7), A2 => n14984, ZN => n8153);
   U2220 : AND2_X1 port map( A1 => n15026, A2 => n14984, ZN => n8063);
   U2221 : AND2_X1 port map( A1 => ADDR_RD2(7), A2 => n14983, ZN => n8152);
   U2222 : INV_X1 port map( A => ADDR_RD1(6), ZN => n5347);
   U2223 : INV_X1 port map( A => ADDR_RD2(6), ZN => n5355);
   U2224 : INV_X1 port map( A => ADDR_RD1(5), ZN => n5348);
   U2225 : INV_X1 port map( A => ADDR_RD2(5), ZN => n5356);
   U2226 : INV_X1 port map( A => ADDR_RD2(4), ZN => n5357);
   U2227 : INV_X1 port map( A => ADDR_RD1(4), ZN => n5349);
   U2228 : INV_X1 port map( A => ADDR_WR(4), ZN => n5280);
   U2229 : INV_X1 port map( A => ADDR_RD2(3), ZN => n5358);
   U2230 : INV_X1 port map( A => ADDR_RD1(3), ZN => n5350);
   U2231 : INV_X1 port map( A => n15266, ZN => n59839);
   U2232 : OAI21_X1 port map( B1 => n15121, B2 => n15247, A => n62197, ZN => 
                           n15266);
   U2233 : INV_X1 port map( A => n15250, ZN => n59929);
   U2234 : OAI21_X1 port map( B1 => n15101, B2 => n15247, A => n62196, ZN => 
                           n15250);
   U2235 : INV_X1 port map( A => n15260, ZN => n59866);
   U2236 : OAI21_X1 port map( B1 => n15115, B2 => n15247, A => n62197, ZN => 
                           n15260);
   U2237 : INV_X1 port map( A => n15267, ZN => n59830);
   U2238 : OAI21_X1 port map( B1 => n15123, B2 => n15247, A => n62197, ZN => 
                           n15267);
   U2239 : INV_X1 port map( A => n15229, ZN => n60100);
   U2240 : OAI21_X1 port map( B1 => n15095, B2 => n15230, A => n62195, ZN => 
                           n15229);
   U2241 : INV_X1 port map( A => n15231, ZN => n60091);
   U2242 : OAI21_X1 port map( B1 => n15097, B2 => n15230, A => n62195, ZN => 
                           n15231);
   U2243 : INV_X1 port map( A => n15232, ZN => n60082);
   U2244 : OAI21_X1 port map( B1 => n15099, B2 => n15230, A => n62195, ZN => 
                           n15232);
   U2245 : INV_X1 port map( A => n15233, ZN => n60073);
   U2246 : OAI21_X1 port map( B1 => n15101, B2 => n15230, A => n62195, ZN => 
                           n15233);
   U2247 : INV_X1 port map( A => n15234, ZN => n60064);
   U2248 : OAI21_X1 port map( B1 => n15103, B2 => n15230, A => n62195, ZN => 
                           n15234);
   U2249 : INV_X1 port map( A => n15235, ZN => n60055);
   U2250 : OAI21_X1 port map( B1 => n15105, B2 => n15230, A => n62195, ZN => 
                           n15235);
   U2251 : INV_X1 port map( A => n15236, ZN => n60046);
   U2252 : OAI21_X1 port map( B1 => n15107, B2 => n15230, A => n62195, ZN => 
                           n15236);
   U2253 : INV_X1 port map( A => n15237, ZN => n60037);
   U2254 : OAI21_X1 port map( B1 => n15109, B2 => n15230, A => n62195, ZN => 
                           n15237);
   U2255 : INV_X1 port map( A => n15238, ZN => n60028);
   U2256 : OAI21_X1 port map( B1 => n15111, B2 => n15230, A => n62195, ZN => 
                           n15238);
   U2257 : INV_X1 port map( A => n15239, ZN => n60019);
   U2258 : OAI21_X1 port map( B1 => n15113, B2 => n15230, A => n62195, ZN => 
                           n15239);
   U2259 : INV_X1 port map( A => n15240, ZN => n60010);
   U2260 : OAI21_X1 port map( B1 => n15115, B2 => n15230, A => n62196, ZN => 
                           n15240);
   U2261 : INV_X1 port map( A => n15241, ZN => n60001);
   U2262 : OAI21_X1 port map( B1 => n15117, B2 => n15230, A => n62195, ZN => 
                           n15241);
   U2263 : INV_X1 port map( A => n15242, ZN => n59992);
   U2264 : OAI21_X1 port map( B1 => n15119, B2 => n15230, A => n62196, ZN => 
                           n15242);
   U2265 : INV_X1 port map( A => n15243, ZN => n59983);
   U2266 : OAI21_X1 port map( B1 => n15121, B2 => n15230, A => n62196, ZN => 
                           n15243);
   U2267 : INV_X1 port map( A => n15244, ZN => n59974);
   U2268 : OAI21_X1 port map( B1 => n15123, B2 => n15230, A => n62196, ZN => 
                           n15244);
   U2269 : INV_X1 port map( A => n15245, ZN => n59965);
   U2270 : OAI21_X1 port map( B1 => n15125, B2 => n15230, A => n62196, ZN => 
                           n15245);
   U2271 : INV_X1 port map( A => n15246, ZN => n59956);
   U2272 : OAI21_X1 port map( B1 => n15095, B2 => n15247, A => n62196, ZN => 
                           n15246);
   U2273 : INV_X1 port map( A => n15248, ZN => n59947);
   U2274 : OAI21_X1 port map( B1 => n15097, B2 => n15247, A => n62196, ZN => 
                           n15248);
   U2275 : INV_X1 port map( A => n15249, ZN => n59938);
   U2276 : OAI21_X1 port map( B1 => n15099, B2 => n15247, A => n62196, ZN => 
                           n15249);
   U2277 : INV_X1 port map( A => n15251, ZN => n59920);
   U2278 : OAI21_X1 port map( B1 => n15103, B2 => n15247, A => n62196, ZN => 
                           n15251);
   U2279 : INV_X1 port map( A => n15252, ZN => n59911);
   U2280 : OAI21_X1 port map( B1 => n15105, B2 => n15247, A => n62196, ZN => 
                           n15252);
   U2281 : INV_X1 port map( A => n15253, ZN => n59902);
   U2282 : OAI21_X1 port map( B1 => n15107, B2 => n15247, A => n62196, ZN => 
                           n15253);
   U2283 : INV_X1 port map( A => n15254, ZN => n59893);
   U2284 : OAI21_X1 port map( B1 => n15109, B2 => n15247, A => n62197, ZN => 
                           n15254);
   U2285 : INV_X1 port map( A => n15255, ZN => n59884);
   U2286 : OAI21_X1 port map( B1 => n15111, B2 => n15247, A => n62197, ZN => 
                           n15255);
   U2287 : INV_X1 port map( A => n15258, ZN => n59875);
   U2288 : OAI21_X1 port map( B1 => n15113, B2 => n15247, A => n62196, ZN => 
                           n15258);
   U2289 : INV_X1 port map( A => n15262, ZN => n59857);
   U2290 : OAI21_X1 port map( B1 => n15117, B2 => n15247, A => n62197, ZN => 
                           n15262);
   U2291 : INV_X1 port map( A => n15264, ZN => n59848);
   U2292 : OAI21_X1 port map( B1 => n15119, B2 => n15247, A => n62197, ZN => 
                           n15264);
   U2293 : INV_X1 port map( A => n15268, ZN => n59821);
   U2294 : OAI21_X1 port map( B1 => n15125, B2 => n15247, A => n62197, ZN => 
                           n15268);
   U2295 : INV_X1 port map( A => n15189, ZN => n60379);
   U2296 : OAI21_X1 port map( B1 => n15097, B2 => n15188, A => n62187, ZN => 
                           n15189);
   U2297 : INV_X1 port map( A => n15190, ZN => n60370);
   U2298 : OAI21_X1 port map( B1 => n15099, B2 => n15188, A => n62187, ZN => 
                           n15190);
   U2299 : INV_X1 port map( A => n15191, ZN => n60361);
   U2300 : OAI21_X1 port map( B1 => n15101, B2 => n15188, A => n62190, ZN => 
                           n15191);
   U2301 : INV_X1 port map( A => n15192, ZN => n60352);
   U2302 : OAI21_X1 port map( B1 => n15103, B2 => n15188, A => n62193, ZN => 
                           n15192);
   U2303 : INV_X1 port map( A => n15193, ZN => n60343);
   U2304 : OAI21_X1 port map( B1 => n15105, B2 => n15188, A => n62193, ZN => 
                           n15193);
   U2305 : INV_X1 port map( A => n15200, ZN => n60280);
   U2306 : OAI21_X1 port map( B1 => n15119, B2 => n15188, A => n62193, ZN => 
                           n15200);
   U2307 : INV_X1 port map( A => n15201, ZN => n60271);
   U2308 : OAI21_X1 port map( B1 => n15121, B2 => n15188, A => n62193, ZN => 
                           n15201);
   U2309 : INV_X1 port map( A => n15215, ZN => n60226);
   U2310 : OAI21_X1 port map( B1 => n15099, B2 => n15213, A => n62194, ZN => 
                           n15215);
   U2311 : INV_X1 port map( A => n15216, ZN => n60217);
   U2312 : OAI21_X1 port map( B1 => n15101, B2 => n15213, A => n62194, ZN => 
                           n15216);
   U2313 : INV_X1 port map( A => n15222, ZN => n60163);
   U2314 : OAI21_X1 port map( B1 => n15113, B2 => n15213, A => n62194, ZN => 
                           n15222);
   U2315 : INV_X1 port map( A => n15223, ZN => n60154);
   U2316 : OAI21_X1 port map( B1 => n15115, B2 => n15213, A => n62194, ZN => 
                           n15223);
   U2317 : INV_X1 port map( A => n15187, ZN => n60388);
   U2318 : OAI21_X1 port map( B1 => n15095, B2 => n15188, A => n62187, ZN => 
                           n15187);
   U2319 : INV_X1 port map( A => n15194, ZN => n60334);
   U2320 : OAI21_X1 port map( B1 => n15107, B2 => n15188, A => n62193, ZN => 
                           n15194);
   U2321 : INV_X1 port map( A => n15195, ZN => n60325);
   U2322 : OAI21_X1 port map( B1 => n15109, B2 => n15188, A => n62193, ZN => 
                           n15195);
   U2323 : INV_X1 port map( A => n15196, ZN => n60316);
   U2324 : OAI21_X1 port map( B1 => n15111, B2 => n15188, A => n62193, ZN => 
                           n15196);
   U2325 : INV_X1 port map( A => n15197, ZN => n60307);
   U2326 : OAI21_X1 port map( B1 => n15113, B2 => n15188, A => n62193, ZN => 
                           n15197);
   U2327 : INV_X1 port map( A => n15198, ZN => n60298);
   U2328 : OAI21_X1 port map( B1 => n15115, B2 => n15188, A => n62193, ZN => 
                           n15198);
   U2329 : INV_X1 port map( A => n15199, ZN => n60289);
   U2330 : OAI21_X1 port map( B1 => n15117, B2 => n15188, A => n62193, ZN => 
                           n15199);
   U2331 : INV_X1 port map( A => n15202, ZN => n60262);
   U2332 : OAI21_X1 port map( B1 => n15123, B2 => n15188, A => n62193, ZN => 
                           n15202);
   U2333 : INV_X1 port map( A => n15211, ZN => n60253);
   U2334 : OAI21_X1 port map( B1 => n15125, B2 => n15188, A => n62193, ZN => 
                           n15211);
   U2335 : INV_X1 port map( A => n15212, ZN => n60244);
   U2336 : OAI21_X1 port map( B1 => n15095, B2 => n15213, A => n62193, ZN => 
                           n15212);
   U2337 : INV_X1 port map( A => n15214, ZN => n60235);
   U2338 : OAI21_X1 port map( B1 => n15097, B2 => n15213, A => n62194, ZN => 
                           n15214);
   U2339 : INV_X1 port map( A => n15217, ZN => n60208);
   U2340 : OAI21_X1 port map( B1 => n15103, B2 => n15213, A => n62194, ZN => 
                           n15217);
   U2341 : INV_X1 port map( A => n15218, ZN => n60199);
   U2342 : OAI21_X1 port map( B1 => n15105, B2 => n15213, A => n62194, ZN => 
                           n15218);
   U2343 : INV_X1 port map( A => n15219, ZN => n60190);
   U2344 : OAI21_X1 port map( B1 => n15107, B2 => n15213, A => n62194, ZN => 
                           n15219);
   U2345 : INV_X1 port map( A => n15220, ZN => n60181);
   U2346 : OAI21_X1 port map( B1 => n15109, B2 => n15213, A => n62194, ZN => 
                           n15220);
   U2347 : INV_X1 port map( A => n15221, ZN => n60172);
   U2348 : OAI21_X1 port map( B1 => n15111, B2 => n15213, A => n62194, ZN => 
                           n15221);
   U2349 : INV_X1 port map( A => n15224, ZN => n60145);
   U2350 : OAI21_X1 port map( B1 => n15117, B2 => n15213, A => n62194, ZN => 
                           n15224);
   U2351 : INV_X1 port map( A => n15225, ZN => n60136);
   U2352 : OAI21_X1 port map( B1 => n15119, B2 => n15213, A => n62194, ZN => 
                           n15225);
   U2353 : INV_X1 port map( A => n15226, ZN => n60127);
   U2354 : OAI21_X1 port map( B1 => n15121, B2 => n15213, A => n62194, ZN => 
                           n15226);
   U2355 : INV_X1 port map( A => n15227, ZN => n60118);
   U2356 : OAI21_X1 port map( B1 => n15123, B2 => n15213, A => n62195, ZN => 
                           n15227);
   U2357 : INV_X1 port map( A => n15228, ZN => n60109);
   U2358 : OAI21_X1 port map( B1 => n15125, B2 => n15213, A => n62195, ZN => 
                           n15228);
   U2359 : INV_X1 port map( A => n15149, ZN => n60658);
   U2360 : OAI21_X1 port map( B1 => n15099, B2 => n15147, A => n62190, ZN => 
                           n15149);
   U2361 : INV_X1 port map( A => n15150, ZN => n60649);
   U2362 : OAI21_X1 port map( B1 => n15101, B2 => n15147, A => n62190, ZN => 
                           n15150);
   U2363 : INV_X1 port map( A => n15153, ZN => n60622);
   U2364 : OAI21_X1 port map( B1 => n15107, B2 => n15147, A => n62189, ZN => 
                           n15153);
   U2365 : INV_X1 port map( A => n15154, ZN => n60613);
   U2366 : OAI21_X1 port map( B1 => n15109, B2 => n15147, A => n62189, ZN => 
                           n15154);
   U2367 : INV_X1 port map( A => n15157, ZN => n60586);
   U2368 : OAI21_X1 port map( B1 => n15115, B2 => n15147, A => n62189, ZN => 
                           n15157);
   U2369 : INV_X1 port map( A => n15158, ZN => n60577);
   U2370 : OAI21_X1 port map( B1 => n15117, B2 => n15147, A => n62189, ZN => 
                           n15158);
   U2371 : INV_X1 port map( A => n15161, ZN => n60550);
   U2372 : OAI21_X1 port map( B1 => n15123, B2 => n15147, A => n62189, ZN => 
                           n15161);
   U2373 : INV_X1 port map( A => n15162, ZN => n60541);
   U2374 : OAI21_X1 port map( B1 => n15125, B2 => n15147, A => n62189, ZN => 
                           n15162);
   U2375 : INV_X1 port map( A => n15169, ZN => n60487);
   U2376 : OAI21_X1 port map( B1 => n15105, B2 => n15164, A => n62188, ZN => 
                           n15169);
   U2377 : INV_X1 port map( A => n15178, ZN => n60469);
   U2378 : OAI21_X1 port map( B1 => n15109, B2 => n15164, A => n62188, ZN => 
                           n15178);
   U2379 : INV_X1 port map( A => n15179, ZN => n60460);
   U2380 : OAI21_X1 port map( B1 => n15111, B2 => n15164, A => n62188, ZN => 
                           n15179);
   U2381 : INV_X1 port map( A => n15184, ZN => n60415);
   U2382 : OAI21_X1 port map( B1 => n15121, B2 => n15164, A => n62188, ZN => 
                           n15184);
   U2383 : INV_X1 port map( A => n15185, ZN => n60406);
   U2384 : OAI21_X1 port map( B1 => n15123, B2 => n15164, A => n62188, ZN => 
                           n15185);
   U2385 : INV_X1 port map( A => n15146, ZN => n60676);
   U2386 : OAI21_X1 port map( B1 => n15095, B2 => n15147, A => n62190, ZN => 
                           n15146);
   U2387 : INV_X1 port map( A => n15148, ZN => n60667);
   U2388 : OAI21_X1 port map( B1 => n15097, B2 => n15147, A => n62190, ZN => 
                           n15148);
   U2389 : INV_X1 port map( A => n15151, ZN => n60640);
   U2390 : OAI21_X1 port map( B1 => n15103, B2 => n15147, A => n62190, ZN => 
                           n15151);
   U2391 : INV_X1 port map( A => n15152, ZN => n60631);
   U2392 : OAI21_X1 port map( B1 => n15105, B2 => n15147, A => n62189, ZN => 
                           n15152);
   U2393 : INV_X1 port map( A => n15155, ZN => n60604);
   U2394 : OAI21_X1 port map( B1 => n15111, B2 => n15147, A => n62192, ZN => 
                           n15155);
   U2395 : INV_X1 port map( A => n15156, ZN => n60595);
   U2396 : OAI21_X1 port map( B1 => n15113, B2 => n15147, A => n62189, ZN => 
                           n15156);
   U2397 : INV_X1 port map( A => n15159, ZN => n60568);
   U2398 : OAI21_X1 port map( B1 => n15119, B2 => n15147, A => n62189, ZN => 
                           n15159);
   U2399 : INV_X1 port map( A => n15160, ZN => n60559);
   U2400 : OAI21_X1 port map( B1 => n15121, B2 => n15147, A => n62189, ZN => 
                           n15160);
   U2401 : INV_X1 port map( A => n15163, ZN => n60532);
   U2402 : OAI21_X1 port map( B1 => n15095, B2 => n15164, A => n62189, ZN => 
                           n15163);
   U2403 : INV_X1 port map( A => n15165, ZN => n60523);
   U2404 : OAI21_X1 port map( B1 => n15097, B2 => n15164, A => n62189, ZN => 
                           n15165);
   U2405 : INV_X1 port map( A => n15166, ZN => n60514);
   U2406 : OAI21_X1 port map( B1 => n15099, B2 => n15164, A => n62189, ZN => 
                           n15166);
   U2407 : INV_X1 port map( A => n15167, ZN => n60505);
   U2408 : OAI21_X1 port map( B1 => n15101, B2 => n15164, A => n62188, ZN => 
                           n15167);
   U2409 : INV_X1 port map( A => n15168, ZN => n60496);
   U2410 : OAI21_X1 port map( B1 => n15103, B2 => n15164, A => n62188, ZN => 
                           n15168);
   U2411 : INV_X1 port map( A => n15170, ZN => n60478);
   U2412 : OAI21_X1 port map( B1 => n15107, B2 => n15164, A => n62188, ZN => 
                           n15170);
   U2413 : INV_X1 port map( A => n15180, ZN => n60451);
   U2414 : OAI21_X1 port map( B1 => n15113, B2 => n15164, A => n62188, ZN => 
                           n15180);
   U2415 : INV_X1 port map( A => n15181, ZN => n60442);
   U2416 : OAI21_X1 port map( B1 => n15115, B2 => n15164, A => n62188, ZN => 
                           n15181);
   U2417 : INV_X1 port map( A => n15182, ZN => n60433);
   U2418 : OAI21_X1 port map( B1 => n15117, B2 => n15164, A => n62188, ZN => 
                           n15182);
   U2419 : INV_X1 port map( A => n15183, ZN => n60424);
   U2420 : OAI21_X1 port map( B1 => n15119, B2 => n15164, A => n62188, ZN => 
                           n15183);
   U2421 : INV_X1 port map( A => n15186, ZN => n60397);
   U2422 : OAI21_X1 port map( B1 => n15125, B2 => n15164, A => n62188, ZN => 
                           n15186);
   U2423 : INV_X1 port map( A => n15133, ZN => n60784);
   U2424 : OAI21_X1 port map( B1 => n15103, B2 => n15129, A => n62191, ZN => 
                           n15133);
   U2425 : INV_X1 port map( A => n15130, ZN => n60811);
   U2426 : OAI21_X1 port map( B1 => n15097, B2 => n15129, A => n62191, ZN => 
                           n15130);
   U2427 : INV_X1 port map( A => n15131, ZN => n60802);
   U2428 : OAI21_X1 port map( B1 => n15099, B2 => n15129, A => n62191, ZN => 
                           n15131);
   U2429 : INV_X1 port map( A => n15108, ZN => n60901);
   U2430 : OAI21_X1 port map( B1 => n15109, B2 => n15094, A => n62192, ZN => 
                           n15108);
   U2431 : INV_X1 port map( A => n15128, ZN => n60820);
   U2432 : OAI21_X1 port map( B1 => n15095, B2 => n15129, A => n62191, ZN => 
                           n15128);
   U2433 : INV_X1 port map( A => n15132, ZN => n60793);
   U2434 : OAI21_X1 port map( B1 => n15101, B2 => n15129, A => n62191, ZN => 
                           n15132);
   U2435 : INV_X1 port map( A => n15134, ZN => n60775);
   U2436 : OAI21_X1 port map( B1 => n15105, B2 => n15129, A => n62191, ZN => 
                           n15134);
   U2437 : INV_X1 port map( A => n15135, ZN => n60766);
   U2438 : OAI21_X1 port map( B1 => n15107, B2 => n15129, A => n62191, ZN => 
                           n15135);
   U2439 : INV_X1 port map( A => n15136, ZN => n60757);
   U2440 : OAI21_X1 port map( B1 => n15109, B2 => n15129, A => n62191, ZN => 
                           n15136);
   U2441 : INV_X1 port map( A => n15102, ZN => n60928);
   U2442 : OAI21_X1 port map( B1 => n15094, B2 => n15103, A => n62192, ZN => 
                           n15102);
   U2443 : INV_X1 port map( A => n15104, ZN => n60919);
   U2444 : OAI21_X1 port map( B1 => n15094, B2 => n15105, A => n62192, ZN => 
                           n15104);
   U2445 : INV_X1 port map( A => n15110, ZN => n60892);
   U2446 : OAI21_X1 port map( B1 => n15094, B2 => n15111, A => n62192, ZN => 
                           n15110);
   U2447 : INV_X1 port map( A => n15112, ZN => n60883);
   U2448 : OAI21_X1 port map( B1 => n15094, B2 => n15113, A => n62192, ZN => 
                           n15112);
   U2449 : INV_X1 port map( A => n15118, ZN => n60856);
   U2450 : OAI21_X1 port map( B1 => n15094, B2 => n15119, A => n62191, ZN => 
                           n15118);
   U2451 : INV_X1 port map( A => n15120, ZN => n60847);
   U2452 : OAI21_X1 port map( B1 => n15094, B2 => n15121, A => n62191, ZN => 
                           n15120);
   U2453 : INV_X1 port map( A => n15122, ZN => n60838);
   U2454 : OAI21_X1 port map( B1 => n15094, B2 => n15123, A => n62191, ZN => 
                           n15122);
   U2455 : INV_X1 port map( A => n15124, ZN => n60829);
   U2456 : OAI21_X1 port map( B1 => n15094, B2 => n15125, A => n62191, ZN => 
                           n15124);
   U2457 : INV_X1 port map( A => n15098, ZN => n60946);
   U2458 : OAI21_X1 port map( B1 => n15094, B2 => n15099, A => n62192, ZN => 
                           n15098);
   U2459 : INV_X1 port map( A => n15100, ZN => n60937);
   U2460 : OAI21_X1 port map( B1 => n15094, B2 => n15101, A => n62192, ZN => 
                           n15100);
   U2461 : INV_X1 port map( A => n15073, ZN => n61244);
   U2462 : OAI21_X1 port map( B1 => n15094, B2 => n15095, A => n62192, ZN => 
                           n15073);
   U2463 : INV_X1 port map( A => n15096, ZN => n60955);
   U2464 : OAI21_X1 port map( B1 => n15094, B2 => n15097, A => n62192, ZN => 
                           n15096);
   U2465 : INV_X1 port map( A => n15106, ZN => n60910);
   U2466 : OAI21_X1 port map( B1 => n15094, B2 => n15107, A => n62192, ZN => 
                           n15106);
   U2467 : INV_X1 port map( A => n15114, ZN => n60874);
   U2468 : OAI21_X1 port map( B1 => n15094, B2 => n15115, A => n62192, ZN => 
                           n15114);
   U2469 : INV_X1 port map( A => n15116, ZN => n60865);
   U2470 : OAI21_X1 port map( B1 => n15094, B2 => n15117, A => n62192, ZN => 
                           n15116);
   U2471 : INV_X1 port map( A => n15140, ZN => n60721);
   U2472 : OAI21_X1 port map( B1 => n15117, B2 => n15129, A => n62190, ZN => 
                           n15140);
   U2473 : INV_X1 port map( A => n15144, ZN => n60685);
   U2474 : OAI21_X1 port map( B1 => n15125, B2 => n15129, A => n62190, ZN => 
                           n15144);
   U2475 : INV_X1 port map( A => n15141, ZN => n60712);
   U2476 : OAI21_X1 port map( B1 => n15119, B2 => n15129, A => n62190, ZN => 
                           n15141);
   U2477 : INV_X1 port map( A => n15137, ZN => n60748);
   U2478 : OAI21_X1 port map( B1 => n15111, B2 => n15129, A => n62191, ZN => 
                           n15137);
   U2479 : INV_X1 port map( A => n15138, ZN => n60739);
   U2480 : OAI21_X1 port map( B1 => n15113, B2 => n15129, A => n62190, ZN => 
                           n15138);
   U2481 : INV_X1 port map( A => n15139, ZN => n60730);
   U2482 : OAI21_X1 port map( B1 => n15115, B2 => n15129, A => n62190, ZN => 
                           n15139);
   U2483 : INV_X1 port map( A => n15142, ZN => n60703);
   U2484 : OAI21_X1 port map( B1 => n15121, B2 => n15129, A => n62190, ZN => 
                           n15142);
   U2485 : INV_X1 port map( A => n15143, ZN => n60694);
   U2486 : OAI21_X1 port map( B1 => n15123, B2 => n15129, A => n62190, ZN => 
                           n15143);
   U2487 : INV_X1 port map( A => n15286, ZN => n59758);
   U2488 : BUF_X1 port map( A => n60998, Z => n61003);
   U2489 : BUF_X1 port map( A => n61012, Z => n61017);
   U2490 : BUF_X1 port map( A => n61026, Z => n61031);
   U2491 : BUF_X1 port map( A => n61040, Z => n61045);
   U2492 : BUF_X1 port map( A => n61054, Z => n61059);
   U2493 : BUF_X1 port map( A => n61068, Z => n61073);
   U2494 : BUF_X1 port map( A => n61082, Z => n61087);
   U2495 : BUF_X1 port map( A => n61096, Z => n61101);
   U2496 : BUF_X1 port map( A => n61110, Z => n61115);
   U2497 : BUF_X1 port map( A => n61124, Z => n61129);
   U2498 : BUF_X1 port map( A => n62103, Z => n62108);
   U2499 : BUF_X1 port map( A => n60956, Z => n60961);
   U2500 : BUF_X1 port map( A => n60970, Z => n60975);
   U2501 : BUF_X1 port map( A => n60984, Z => n60989);
   U2502 : BUF_X1 port map( A => n61963, Z => n61968);
   U2503 : BUF_X1 port map( A => n61977, Z => n61982);
   U2504 : BUF_X1 port map( A => n61991, Z => n61996);
   U2505 : BUF_X1 port map( A => n62005, Z => n62010);
   U2506 : BUF_X1 port map( A => n62019, Z => n62024);
   U2507 : BUF_X1 port map( A => n62033, Z => n62038);
   U2508 : BUF_X1 port map( A => n62047, Z => n62052);
   U2509 : BUF_X1 port map( A => n62061, Z => n62066);
   U2510 : BUF_X1 port map( A => n62075, Z => n62080);
   U2511 : BUF_X1 port map( A => n62089, Z => n62094);
   U2512 : BUF_X1 port map( A => n61963, Z => n61969);
   U2513 : BUF_X1 port map( A => n61977, Z => n61983);
   U2514 : BUF_X1 port map( A => n61991, Z => n61997);
   U2515 : BUF_X1 port map( A => n62005, Z => n62011);
   U2516 : BUF_X1 port map( A => n62019, Z => n62025);
   U2517 : BUF_X1 port map( A => n62033, Z => n62039);
   U2518 : BUF_X1 port map( A => n62047, Z => n62053);
   U2519 : BUF_X1 port map( A => n62061, Z => n62067);
   U2520 : BUF_X1 port map( A => n62075, Z => n62081);
   U2521 : BUF_X1 port map( A => n62089, Z => n62095);
   U2522 : BUF_X1 port map( A => n62103, Z => n62109);
   U2523 : BUF_X1 port map( A => n60956, Z => n60962);
   U2524 : BUF_X1 port map( A => n60970, Z => n60976);
   U2525 : BUF_X1 port map( A => n60984, Z => n60990);
   U2526 : BUF_X1 port map( A => n60998, Z => n61004);
   U2527 : BUF_X1 port map( A => n61012, Z => n61018);
   U2528 : BUF_X1 port map( A => n61026, Z => n61032);
   U2529 : BUF_X1 port map( A => n61040, Z => n61046);
   U2530 : BUF_X1 port map( A => n61054, Z => n61060);
   U2531 : BUF_X1 port map( A => n61068, Z => n61074);
   U2532 : BUF_X1 port map( A => n61082, Z => n61088);
   U2533 : BUF_X1 port map( A => n61096, Z => n61102);
   U2534 : BUF_X1 port map( A => n61110, Z => n61116);
   U2535 : BUF_X1 port map( A => n61124, Z => n61130);
   U2536 : BUF_X1 port map( A => n61963, Z => n61965);
   U2537 : BUF_X1 port map( A => n61977, Z => n61979);
   U2538 : BUF_X1 port map( A => n61991, Z => n61993);
   U2539 : BUF_X1 port map( A => n62005, Z => n62007);
   U2540 : BUF_X1 port map( A => n62019, Z => n62021);
   U2541 : BUF_X1 port map( A => n62033, Z => n62035);
   U2542 : BUF_X1 port map( A => n62047, Z => n62049);
   U2543 : BUF_X1 port map( A => n62061, Z => n62063);
   U2544 : BUF_X1 port map( A => n62075, Z => n62077);
   U2545 : BUF_X1 port map( A => n62089, Z => n62091);
   U2546 : BUF_X1 port map( A => n62103, Z => n62105);
   U2547 : BUF_X1 port map( A => n60956, Z => n60958);
   U2548 : BUF_X1 port map( A => n60970, Z => n60972);
   U2549 : BUF_X1 port map( A => n60984, Z => n60986);
   U2550 : BUF_X1 port map( A => n60998, Z => n61000);
   U2551 : BUF_X1 port map( A => n61012, Z => n61014);
   U2552 : BUF_X1 port map( A => n61026, Z => n61028);
   U2553 : BUF_X1 port map( A => n61040, Z => n61042);
   U2554 : BUF_X1 port map( A => n61054, Z => n61056);
   U2555 : BUF_X1 port map( A => n61068, Z => n61070);
   U2556 : BUF_X1 port map( A => n61082, Z => n61084);
   U2557 : BUF_X1 port map( A => n61096, Z => n61098);
   U2558 : BUF_X1 port map( A => n61110, Z => n61112);
   U2559 : BUF_X1 port map( A => n61124, Z => n61126);
   U2560 : BUF_X1 port map( A => n61963, Z => n61970);
   U2561 : BUF_X1 port map( A => n61977, Z => n61984);
   U2562 : BUF_X1 port map( A => n61991, Z => n61998);
   U2563 : BUF_X1 port map( A => n62005, Z => n62012);
   U2564 : BUF_X1 port map( A => n62019, Z => n62026);
   U2565 : BUF_X1 port map( A => n62033, Z => n62040);
   U2566 : BUF_X1 port map( A => n62047, Z => n62054);
   U2567 : BUF_X1 port map( A => n62061, Z => n62068);
   U2568 : BUF_X1 port map( A => n62075, Z => n62082);
   U2569 : BUF_X1 port map( A => n62089, Z => n62096);
   U2570 : BUF_X1 port map( A => n62103, Z => n62110);
   U2571 : BUF_X1 port map( A => n60956, Z => n60963);
   U2572 : BUF_X1 port map( A => n60970, Z => n60977);
   U2573 : BUF_X1 port map( A => n60984, Z => n60991);
   U2574 : BUF_X1 port map( A => n60998, Z => n61005);
   U2575 : BUF_X1 port map( A => n61012, Z => n61019);
   U2576 : BUF_X1 port map( A => n61026, Z => n61033);
   U2577 : BUF_X1 port map( A => n61040, Z => n61047);
   U2578 : BUF_X1 port map( A => n61054, Z => n61061);
   U2579 : BUF_X1 port map( A => n61068, Z => n61075);
   U2580 : BUF_X1 port map( A => n61082, Z => n61089);
   U2581 : BUF_X1 port map( A => n61096, Z => n61103);
   U2582 : BUF_X1 port map( A => n61110, Z => n61117);
   U2583 : BUF_X1 port map( A => n61124, Z => n61131);
   U2584 : BUF_X1 port map( A => n61963, Z => n61966);
   U2585 : BUF_X1 port map( A => n61977, Z => n61980);
   U2586 : BUF_X1 port map( A => n61991, Z => n61994);
   U2587 : BUF_X1 port map( A => n62005, Z => n62008);
   U2588 : BUF_X1 port map( A => n62019, Z => n62022);
   U2589 : BUF_X1 port map( A => n62033, Z => n62036);
   U2590 : BUF_X1 port map( A => n62047, Z => n62050);
   U2591 : BUF_X1 port map( A => n62061, Z => n62064);
   U2592 : BUF_X1 port map( A => n62075, Z => n62078);
   U2593 : BUF_X1 port map( A => n62089, Z => n62092);
   U2594 : BUF_X1 port map( A => n62103, Z => n62106);
   U2595 : BUF_X1 port map( A => n60956, Z => n60959);
   U2596 : BUF_X1 port map( A => n60970, Z => n60973);
   U2597 : BUF_X1 port map( A => n60984, Z => n60987);
   U2598 : BUF_X1 port map( A => n60998, Z => n61001);
   U2599 : BUF_X1 port map( A => n61012, Z => n61015);
   U2600 : BUF_X1 port map( A => n61026, Z => n61029);
   U2601 : BUF_X1 port map( A => n61040, Z => n61043);
   U2602 : BUF_X1 port map( A => n61054, Z => n61057);
   U2603 : BUF_X1 port map( A => n61068, Z => n61071);
   U2604 : BUF_X1 port map( A => n61082, Z => n61085);
   U2605 : BUF_X1 port map( A => n61096, Z => n61099);
   U2606 : BUF_X1 port map( A => n61110, Z => n61113);
   U2607 : BUF_X1 port map( A => n61124, Z => n61127);
   U2608 : BUF_X1 port map( A => n61963, Z => n61967);
   U2609 : BUF_X1 port map( A => n61977, Z => n61981);
   U2610 : BUF_X1 port map( A => n61991, Z => n61995);
   U2611 : BUF_X1 port map( A => n62005, Z => n62009);
   U2612 : BUF_X1 port map( A => n62019, Z => n62023);
   U2613 : BUF_X1 port map( A => n62033, Z => n62037);
   U2614 : BUF_X1 port map( A => n62047, Z => n62051);
   U2615 : BUF_X1 port map( A => n62061, Z => n62065);
   U2616 : BUF_X1 port map( A => n62075, Z => n62079);
   U2617 : BUF_X1 port map( A => n62089, Z => n62093);
   U2618 : BUF_X1 port map( A => n62103, Z => n62107);
   U2619 : BUF_X1 port map( A => n60956, Z => n60960);
   U2620 : BUF_X1 port map( A => n60970, Z => n60974);
   U2621 : BUF_X1 port map( A => n60984, Z => n60988);
   U2622 : BUF_X1 port map( A => n60998, Z => n61002);
   U2623 : BUF_X1 port map( A => n61012, Z => n61016);
   U2624 : BUF_X1 port map( A => n61026, Z => n61030);
   U2625 : BUF_X1 port map( A => n61040, Z => n61044);
   U2626 : BUF_X1 port map( A => n61054, Z => n61058);
   U2627 : BUF_X1 port map( A => n61068, Z => n61072);
   U2628 : BUF_X1 port map( A => n61082, Z => n61086);
   U2629 : BUF_X1 port map( A => n61096, Z => n61100);
   U2630 : BUF_X1 port map( A => n61110, Z => n61114);
   U2631 : BUF_X1 port map( A => n61124, Z => n61128);
   U2632 : BUF_X1 port map( A => n61138, Z => n61143);
   U2633 : BUF_X1 port map( A => n61152, Z => n61157);
   U2634 : BUF_X1 port map( A => n61166, Z => n61171);
   U2635 : BUF_X1 port map( A => n61180, Z => n61185);
   U2636 : BUF_X1 port map( A => n61194, Z => n61199);
   U2637 : BUF_X1 port map( A => n61208, Z => n61213);
   U2638 : BUF_X1 port map( A => n61222, Z => n61227);
   U2639 : BUF_X1 port map( A => n61245, Z => n61250);
   U2640 : BUF_X1 port map( A => n61138, Z => n61144);
   U2641 : BUF_X1 port map( A => n61152, Z => n61158);
   U2642 : BUF_X1 port map( A => n61166, Z => n61172);
   U2643 : BUF_X1 port map( A => n61180, Z => n61186);
   U2644 : BUF_X1 port map( A => n61194, Z => n61200);
   U2645 : BUF_X1 port map( A => n61208, Z => n61214);
   U2646 : BUF_X1 port map( A => n61222, Z => n61228);
   U2647 : BUF_X1 port map( A => n61245, Z => n61251);
   U2648 : BUF_X1 port map( A => n61138, Z => n61140);
   U2649 : BUF_X1 port map( A => n61152, Z => n61154);
   U2650 : BUF_X1 port map( A => n61166, Z => n61168);
   U2651 : BUF_X1 port map( A => n61180, Z => n61182);
   U2652 : BUF_X1 port map( A => n61194, Z => n61196);
   U2653 : BUF_X1 port map( A => n61208, Z => n61210);
   U2654 : BUF_X1 port map( A => n61222, Z => n61224);
   U2655 : BUF_X1 port map( A => n61245, Z => n61247);
   U2656 : BUF_X1 port map( A => n61138, Z => n61145);
   U2657 : BUF_X1 port map( A => n61152, Z => n61159);
   U2658 : BUF_X1 port map( A => n61166, Z => n61173);
   U2659 : BUF_X1 port map( A => n61180, Z => n61187);
   U2660 : BUF_X1 port map( A => n61194, Z => n61201);
   U2661 : BUF_X1 port map( A => n61208, Z => n61215);
   U2662 : BUF_X1 port map( A => n61222, Z => n61229);
   U2663 : BUF_X1 port map( A => n61245, Z => n61252);
   U2664 : BUF_X1 port map( A => n61138, Z => n61141);
   U2665 : BUF_X1 port map( A => n61152, Z => n61155);
   U2666 : BUF_X1 port map( A => n61166, Z => n61169);
   U2667 : BUF_X1 port map( A => n61180, Z => n61183);
   U2668 : BUF_X1 port map( A => n61194, Z => n61197);
   U2669 : BUF_X1 port map( A => n61208, Z => n61211);
   U2670 : BUF_X1 port map( A => n61222, Z => n61225);
   U2671 : BUF_X1 port map( A => n61245, Z => n61248);
   U2672 : BUF_X1 port map( A => n61138, Z => n61142);
   U2673 : BUF_X1 port map( A => n61152, Z => n61156);
   U2674 : BUF_X1 port map( A => n61166, Z => n61170);
   U2675 : BUF_X1 port map( A => n61180, Z => n61184);
   U2676 : BUF_X1 port map( A => n61194, Z => n61198);
   U2677 : BUF_X1 port map( A => n61208, Z => n61212);
   U2678 : BUF_X1 port map( A => n61222, Z => n61226);
   U2679 : BUF_X1 port map( A => n61245, Z => n61249);
   U2680 : BUF_X1 port map( A => n60957, Z => n60966);
   U2681 : BUF_X1 port map( A => n61083, Z => n61092);
   U2682 : BUF_X1 port map( A => n61097, Z => n61106);
   U2683 : BUF_X1 port map( A => n61111, Z => n61120);
   U2684 : BUF_X1 port map( A => n61125, Z => n61134);
   U2685 : BUF_X1 port map( A => n60971, Z => n60980);
   U2686 : BUF_X1 port map( A => n60985, Z => n60994);
   U2687 : BUF_X1 port map( A => n60999, Z => n61008);
   U2688 : BUF_X1 port map( A => n61013, Z => n61022);
   U2689 : BUF_X1 port map( A => n61027, Z => n61036);
   U2690 : BUF_X1 port map( A => n61041, Z => n61050);
   U2691 : BUF_X1 port map( A => n61055, Z => n61064);
   U2692 : BUF_X1 port map( A => n61069, Z => n61078);
   U2693 : BUF_X1 port map( A => n61964, Z => n61973);
   U2694 : BUF_X1 port map( A => n61978, Z => n61987);
   U2695 : BUF_X1 port map( A => n61992, Z => n62001);
   U2696 : BUF_X1 port map( A => n62006, Z => n62015);
   U2697 : BUF_X1 port map( A => n62020, Z => n62029);
   U2698 : BUF_X1 port map( A => n62034, Z => n62043);
   U2699 : BUF_X1 port map( A => n62048, Z => n62057);
   U2700 : BUF_X1 port map( A => n62062, Z => n62071);
   U2701 : BUF_X1 port map( A => n62076, Z => n62085);
   U2702 : BUF_X1 port map( A => n62090, Z => n62099);
   U2703 : BUF_X1 port map( A => n62104, Z => n62113);
   U2704 : BUF_X1 port map( A => n60957, Z => n60967);
   U2705 : BUF_X1 port map( A => n60971, Z => n60981);
   U2706 : BUF_X1 port map( A => n60985, Z => n60995);
   U2707 : BUF_X1 port map( A => n60999, Z => n61009);
   U2708 : BUF_X1 port map( A => n61013, Z => n61023);
   U2709 : BUF_X1 port map( A => n61027, Z => n61037);
   U2710 : BUF_X1 port map( A => n61041, Z => n61051);
   U2711 : BUF_X1 port map( A => n61055, Z => n61065);
   U2712 : BUF_X1 port map( A => n61069, Z => n61079);
   U2713 : BUF_X1 port map( A => n61083, Z => n61093);
   U2714 : BUF_X1 port map( A => n61097, Z => n61107);
   U2715 : BUF_X1 port map( A => n61111, Z => n61121);
   U2716 : BUF_X1 port map( A => n61125, Z => n61135);
   U2717 : BUF_X1 port map( A => n61964, Z => n61974);
   U2718 : BUF_X1 port map( A => n61978, Z => n61988);
   U2719 : BUF_X1 port map( A => n61992, Z => n62002);
   U2720 : BUF_X1 port map( A => n62006, Z => n62016);
   U2721 : BUF_X1 port map( A => n62020, Z => n62030);
   U2722 : BUF_X1 port map( A => n62034, Z => n62044);
   U2723 : BUF_X1 port map( A => n62048, Z => n62058);
   U2724 : BUF_X1 port map( A => n62062, Z => n62072);
   U2725 : BUF_X1 port map( A => n62076, Z => n62086);
   U2726 : BUF_X1 port map( A => n62090, Z => n62100);
   U2727 : BUF_X1 port map( A => n62104, Z => n62114);
   U2728 : BUF_X1 port map( A => n61964, Z => n61971);
   U2729 : BUF_X1 port map( A => n61978, Z => n61985);
   U2730 : BUF_X1 port map( A => n61992, Z => n61999);
   U2731 : BUF_X1 port map( A => n62006, Z => n62013);
   U2732 : BUF_X1 port map( A => n62020, Z => n62027);
   U2733 : BUF_X1 port map( A => n62034, Z => n62041);
   U2734 : BUF_X1 port map( A => n62048, Z => n62055);
   U2735 : BUF_X1 port map( A => n62062, Z => n62069);
   U2736 : BUF_X1 port map( A => n62076, Z => n62083);
   U2737 : BUF_X1 port map( A => n62090, Z => n62097);
   U2738 : BUF_X1 port map( A => n62104, Z => n62111);
   U2739 : BUF_X1 port map( A => n60957, Z => n60964);
   U2740 : BUF_X1 port map( A => n60971, Z => n60978);
   U2741 : BUF_X1 port map( A => n60985, Z => n60992);
   U2742 : BUF_X1 port map( A => n60999, Z => n61006);
   U2743 : BUF_X1 port map( A => n61013, Z => n61020);
   U2744 : BUF_X1 port map( A => n61027, Z => n61034);
   U2745 : BUF_X1 port map( A => n61041, Z => n61048);
   U2746 : BUF_X1 port map( A => n61055, Z => n61062);
   U2747 : BUF_X1 port map( A => n61069, Z => n61076);
   U2748 : BUF_X1 port map( A => n61083, Z => n61090);
   U2749 : BUF_X1 port map( A => n61097, Z => n61104);
   U2750 : BUF_X1 port map( A => n61111, Z => n61118);
   U2751 : BUF_X1 port map( A => n61125, Z => n61132);
   U2752 : BUF_X1 port map( A => n61964, Z => n61972);
   U2753 : BUF_X1 port map( A => n61978, Z => n61986);
   U2754 : BUF_X1 port map( A => n61992, Z => n62000);
   U2755 : BUF_X1 port map( A => n62006, Z => n62014);
   U2756 : BUF_X1 port map( A => n62020, Z => n62028);
   U2757 : BUF_X1 port map( A => n62034, Z => n62042);
   U2758 : BUF_X1 port map( A => n62048, Z => n62056);
   U2759 : BUF_X1 port map( A => n62062, Z => n62070);
   U2760 : BUF_X1 port map( A => n62076, Z => n62084);
   U2761 : BUF_X1 port map( A => n62090, Z => n62098);
   U2762 : BUF_X1 port map( A => n62104, Z => n62112);
   U2763 : BUF_X1 port map( A => n60957, Z => n60965);
   U2764 : BUF_X1 port map( A => n60971, Z => n60979);
   U2765 : BUF_X1 port map( A => n60985, Z => n60993);
   U2766 : BUF_X1 port map( A => n60999, Z => n61007);
   U2767 : BUF_X1 port map( A => n61013, Z => n61021);
   U2768 : BUF_X1 port map( A => n61027, Z => n61035);
   U2769 : BUF_X1 port map( A => n61041, Z => n61049);
   U2770 : BUF_X1 port map( A => n61055, Z => n61063);
   U2771 : BUF_X1 port map( A => n61069, Z => n61077);
   U2772 : BUF_X1 port map( A => n61083, Z => n61091);
   U2773 : BUF_X1 port map( A => n61097, Z => n61105);
   U2774 : BUF_X1 port map( A => n61111, Z => n61119);
   U2775 : BUF_X1 port map( A => n61125, Z => n61133);
   U2776 : BUF_X1 port map( A => n60957, Z => n60968);
   U2777 : BUF_X1 port map( A => n60971, Z => n60982);
   U2778 : BUF_X1 port map( A => n60985, Z => n60996);
   U2779 : BUF_X1 port map( A => n60999, Z => n61010);
   U2780 : BUF_X1 port map( A => n61013, Z => n61024);
   U2781 : BUF_X1 port map( A => n61027, Z => n61038);
   U2782 : BUF_X1 port map( A => n61041, Z => n61052);
   U2783 : BUF_X1 port map( A => n61055, Z => n61066);
   U2784 : BUF_X1 port map( A => n61069, Z => n61080);
   U2785 : BUF_X1 port map( A => n61083, Z => n61094);
   U2786 : BUF_X1 port map( A => n61097, Z => n61108);
   U2787 : BUF_X1 port map( A => n61111, Z => n61122);
   U2788 : BUF_X1 port map( A => n61125, Z => n61136);
   U2789 : BUF_X1 port map( A => n61964, Z => n61975);
   U2790 : BUF_X1 port map( A => n61978, Z => n61989);
   U2791 : BUF_X1 port map( A => n61992, Z => n62003);
   U2792 : BUF_X1 port map( A => n62006, Z => n62017);
   U2793 : BUF_X1 port map( A => n62020, Z => n62031);
   U2794 : BUF_X1 port map( A => n62034, Z => n62045);
   U2795 : BUF_X1 port map( A => n62048, Z => n62059);
   U2796 : BUF_X1 port map( A => n62062, Z => n62073);
   U2797 : BUF_X1 port map( A => n62076, Z => n62087);
   U2798 : BUF_X1 port map( A => n62090, Z => n62101);
   U2799 : BUF_X1 port map( A => n62104, Z => n62115);
   U2800 : BUF_X1 port map( A => n61139, Z => n61148);
   U2801 : BUF_X1 port map( A => n61153, Z => n61162);
   U2802 : BUF_X1 port map( A => n61167, Z => n61176);
   U2803 : BUF_X1 port map( A => n61181, Z => n61190);
   U2804 : BUF_X1 port map( A => n61195, Z => n61204);
   U2805 : BUF_X1 port map( A => n61209, Z => n61218);
   U2806 : BUF_X1 port map( A => n61223, Z => n61232);
   U2807 : BUF_X1 port map( A => n61246, Z => n61255);
   U2808 : BUF_X1 port map( A => n61139, Z => n61149);
   U2809 : BUF_X1 port map( A => n61153, Z => n61163);
   U2810 : BUF_X1 port map( A => n61167, Z => n61177);
   U2811 : BUF_X1 port map( A => n61181, Z => n61191);
   U2812 : BUF_X1 port map( A => n61195, Z => n61205);
   U2813 : BUF_X1 port map( A => n61209, Z => n61219);
   U2814 : BUF_X1 port map( A => n61223, Z => n61233);
   U2815 : BUF_X1 port map( A => n61246, Z => n61256);
   U2816 : BUF_X1 port map( A => n61139, Z => n61146);
   U2817 : BUF_X1 port map( A => n61153, Z => n61160);
   U2818 : BUF_X1 port map( A => n61167, Z => n61174);
   U2819 : BUF_X1 port map( A => n61181, Z => n61188);
   U2820 : BUF_X1 port map( A => n61195, Z => n61202);
   U2821 : BUF_X1 port map( A => n61209, Z => n61216);
   U2822 : BUF_X1 port map( A => n61223, Z => n61230);
   U2823 : BUF_X1 port map( A => n61246, Z => n61253);
   U2824 : BUF_X1 port map( A => n61139, Z => n61147);
   U2825 : BUF_X1 port map( A => n61153, Z => n61161);
   U2826 : BUF_X1 port map( A => n61167, Z => n61175);
   U2827 : BUF_X1 port map( A => n61181, Z => n61189);
   U2828 : BUF_X1 port map( A => n61195, Z => n61203);
   U2829 : BUF_X1 port map( A => n61209, Z => n61217);
   U2830 : BUF_X1 port map( A => n61223, Z => n61231);
   U2831 : BUF_X1 port map( A => n61246, Z => n61254);
   U2832 : BUF_X1 port map( A => n61139, Z => n61150);
   U2833 : BUF_X1 port map( A => n61153, Z => n61164);
   U2834 : BUF_X1 port map( A => n61167, Z => n61178);
   U2835 : BUF_X1 port map( A => n61181, Z => n61192);
   U2836 : BUF_X1 port map( A => n61195, Z => n61206);
   U2837 : BUF_X1 port map( A => n61209, Z => n61220);
   U2838 : BUF_X1 port map( A => n61223, Z => n61234);
   U2839 : BUF_X1 port map( A => n61246, Z => n61257);
   U2840 : BUF_X1 port map( A => n62183, Z => n62196);
   U2841 : BUF_X1 port map( A => n62182, Z => n62189);
   U2842 : BUF_X1 port map( A => n62182, Z => n62188);
   U2843 : BUF_X1 port map( A => n62183, Z => n62192);
   U2844 : BUF_X1 port map( A => n62183, Z => n62193);
   U2845 : BUF_X1 port map( A => n62183, Z => n62194);
   U2846 : BUF_X1 port map( A => n62183, Z => n62195);
   U2847 : BUF_X1 port map( A => n62183, Z => n62191);
   U2848 : BUF_X1 port map( A => n62182, Z => n62190);
   U2849 : BUF_X1 port map( A => n62184, Z => n62197);
   U2850 : BUF_X1 port map( A => n62182, Z => n62185);
   U2851 : BUF_X1 port map( A => n62182, Z => n62186);
   U2852 : BUF_X1 port map( A => n62182, Z => n62187);
   U2853 : INV_X1 port map( A => ADDR_WR(7), ZN => n5277);
   U2854 : NOR4_X1 port map( A1 => n6754, A2 => n6755, A3 => n6756, A4 => n6757
                           , ZN => n6753);
   U2855 : OAI221_X1 port map( B1 => n61859, B2 => n2482, C1 => n61856, C2 => 
                           n2534, A => n6760, ZN => n6755);
   U2856 : OAI221_X1 port map( B1 => n61693, B2 => n2606, C1 => n61696, C2 => 
                           n2630, A => n6759, ZN => n6756);
   U2857 : OAI221_X1 port map( B1 => n61847, B2 => n2234, C1 => n61844, C2 => 
                           n2294, A => n6761, ZN => n6754);
   U2858 : NOR4_X1 port map( A1 => n6679, A2 => n6680, A3 => n6681, A4 => n6682
                           , ZN => n6678);
   U2859 : OAI221_X1 port map( B1 => n61859, B2 => n2481, C1 => n61856, C2 => 
                           n2533, A => n6685, ZN => n6680);
   U2860 : OAI221_X1 port map( B1 => n6073, B2 => n2605, C1 => n61696, C2 => 
                           n2629, A => n6684, ZN => n6681);
   U2861 : OAI221_X1 port map( B1 => n61847, B2 => n2233, C1 => n61844, C2 => 
                           n2293, A => n6686, ZN => n6679);
   U2862 : NOR4_X1 port map( A1 => n6604, A2 => n6605, A3 => n6606, A4 => n6607
                           , ZN => n6603);
   U2863 : OAI221_X1 port map( B1 => n61859, B2 => n2480, C1 => n61856, C2 => 
                           n2532, A => n6610, ZN => n6605);
   U2864 : OAI221_X1 port map( B1 => n6073, B2 => n2604, C1 => n61696, C2 => 
                           n2628, A => n6609, ZN => n6606);
   U2865 : OAI221_X1 port map( B1 => n61847, B2 => n2232, C1 => n61844, C2 => 
                           n2292, A => n6611, ZN => n6604);
   U2866 : NOR4_X1 port map( A1 => n6529, A2 => n6530, A3 => n6531, A4 => n6532
                           , ZN => n6528);
   U2867 : OAI221_X1 port map( B1 => n61859, B2 => n2479, C1 => n61856, C2 => 
                           n2531, A => n6535, ZN => n6530);
   U2868 : OAI221_X1 port map( B1 => n6073, B2 => n2603, C1 => n61696, C2 => 
                           n2627, A => n6534, ZN => n6531);
   U2869 : OAI221_X1 port map( B1 => n61847, B2 => n2231, C1 => n61844, C2 => 
                           n2291, A => n6536, ZN => n6529);
   U2870 : NOR4_X1 port map( A1 => n6454, A2 => n6455, A3 => n6456, A4 => n6457
                           , ZN => n6453);
   U2871 : OAI221_X1 port map( B1 => n61859, B2 => n2478, C1 => n61856, C2 => 
                           n2530, A => n6460, ZN => n6455);
   U2872 : OAI221_X1 port map( B1 => n6073, B2 => n2602, C1 => n61696, C2 => 
                           n2626, A => n6459, ZN => n6456);
   U2873 : OAI221_X1 port map( B1 => n61847, B2 => n2230, C1 => n61844, C2 => 
                           n2290, A => n6461, ZN => n6454);
   U2874 : NOR4_X1 port map( A1 => n6379, A2 => n6380, A3 => n6381, A4 => n6382
                           , ZN => n6378);
   U2875 : OAI221_X1 port map( B1 => n61859, B2 => n2477, C1 => n61856, C2 => 
                           n2529, A => n6385, ZN => n6380);
   U2876 : OAI221_X1 port map( B1 => n6073, B2 => n2601, C1 => n61696, C2 => 
                           n2625, A => n6384, ZN => n6381);
   U2877 : OAI221_X1 port map( B1 => n61847, B2 => n2229, C1 => n61844, C2 => 
                           n2289, A => n6386, ZN => n6379);
   U2878 : NOR4_X1 port map( A1 => n6304, A2 => n6305, A3 => n6306, A4 => n6307
                           , ZN => n6303);
   U2879 : OAI221_X1 port map( B1 => n61859, B2 => n2476, C1 => n61856, C2 => 
                           n2528, A => n6310, ZN => n6305);
   U2880 : OAI221_X1 port map( B1 => n6073, B2 => n2600, C1 => n61696, C2 => 
                           n2624, A => n6309, ZN => n6306);
   U2881 : OAI221_X1 port map( B1 => n61847, B2 => n2228, C1 => n61844, C2 => 
                           n2288, A => n6311, ZN => n6304);
   U2882 : NOR4_X1 port map( A1 => n6229, A2 => n6230, A3 => n6231, A4 => n6232
                           , ZN => n6228);
   U2883 : OAI221_X1 port map( B1 => n61859, B2 => n2475, C1 => n61856, C2 => 
                           n2527, A => n6235, ZN => n6230);
   U2884 : OAI221_X1 port map( B1 => n6073, B2 => n2599, C1 => n61696, C2 => 
                           n2623, A => n6234, ZN => n6231);
   U2885 : OAI221_X1 port map( B1 => n61847, B2 => n2227, C1 => n61844, C2 => 
                           n2287, A => n6236, ZN => n6229);
   U2886 : NOR4_X1 port map( A1 => n6154, A2 => n6155, A3 => n6156, A4 => n6157
                           , ZN => n6153);
   U2887 : OAI221_X1 port map( B1 => n61859, B2 => n2474, C1 => n61856, C2 => 
                           n2526, A => n6160, ZN => n6155);
   U2888 : OAI221_X1 port map( B1 => n6073, B2 => n2598, C1 => n61696, C2 => 
                           n2622, A => n6159, ZN => n6156);
   U2889 : OAI221_X1 port map( B1 => n61847, B2 => n2226, C1 => n61844, C2 => 
                           n2286, A => n6161, ZN => n6154);
   U2890 : NOR4_X1 port map( A1 => n7129, A2 => n7130, A3 => n7131, A4 => n7132
                           , ZN => n7128);
   U2891 : OAI221_X1 port map( B1 => n61858, B2 => n2515, C1 => n61855, C2 => 
                           n2539, A => n7135, ZN => n7130);
   U2892 : OAI221_X1 port map( B1 => n61693, B2 => n2611, C1 => n61695, C2 => 
                           n2635, A => n7134, ZN => n7131);
   U2893 : OAI221_X1 port map( B1 => n61846, B2 => n2275, C1 => n61843, C2 => 
                           n2391, A => n7136, ZN => n7129);
   U2894 : NOR4_X1 port map( A1 => n7054, A2 => n7055, A3 => n7056, A4 => n7057
                           , ZN => n7053);
   U2895 : OAI221_X1 port map( B1 => n61858, B2 => n2514, C1 => n61855, C2 => 
                           n2538, A => n7060, ZN => n7055);
   U2896 : OAI221_X1 port map( B1 => n61693, B2 => n2610, C1 => n61695, C2 => 
                           n2634, A => n7059, ZN => n7056);
   U2897 : OAI221_X1 port map( B1 => n61846, B2 => n2274, C1 => n61843, C2 => 
                           n2298, A => n7061, ZN => n7054);
   U2898 : NOR4_X1 port map( A1 => n6904, A2 => n6905, A3 => n6906, A4 => n6907
                           , ZN => n6903);
   U2899 : OAI221_X1 port map( B1 => n61859, B2 => n2512, C1 => n61856, C2 => 
                           n2536, A => n6910, ZN => n6905);
   U2900 : OAI221_X1 port map( B1 => n6073, B2 => n2608, C1 => n61696, C2 => 
                           n2632, A => n6909, ZN => n6906);
   U2901 : OAI221_X1 port map( B1 => n61847, B2 => n2272, C1 => n61844, C2 => 
                           n2296, A => n6911, ZN => n6904);
   U2902 : NOR4_X1 port map( A1 => n6829, A2 => n6830, A3 => n6831, A4 => n6832
                           , ZN => n6828);
   U2903 : OAI221_X1 port map( B1 => n61859, B2 => n2511, C1 => n61856, C2 => 
                           n2535, A => n6835, ZN => n6830);
   U2904 : OAI221_X1 port map( B1 => n6073, B2 => n2607, C1 => n61696, C2 => 
                           n2631, A => n6834, ZN => n6831);
   U2905 : OAI221_X1 port map( B1 => n61847, B2 => n2271, C1 => n61844, C2 => 
                           n2295, A => n6836, ZN => n6829);
   U2906 : NOR4_X1 port map( A1 => n7279, A2 => n7280, A3 => n7281, A4 => n7282
                           , ZN => n7278);
   U2907 : OAI221_X1 port map( B1 => n61858, B2 => n2517, C1 => n61855, C2 => 
                           n2541, A => n7285, ZN => n7280);
   U2908 : OAI221_X1 port map( B1 => n61693, B2 => n2613, C1 => n61695, C2 => 
                           n2637, A => n7284, ZN => n7281);
   U2909 : OAI221_X1 port map( B1 => n61846, B2 => n2277, C1 => n61843, C2 => 
                           n2393, A => n7286, ZN => n7279);
   U2910 : NOR4_X1 port map( A1 => n7904, A2 => n7905, A3 => n7906, A4 => n7907
                           , ZN => n7903);
   U2911 : OAI221_X1 port map( B1 => n61858, B2 => n2525, C1 => n61855, C2 => 
                           n2549, A => n7911, ZN => n7905);
   U2912 : OAI221_X1 port map( B1 => n61693, B2 => n2621, C1 => n61695, C2 => 
                           n2652, A => n7909, ZN => n7906);
   U2913 : OAI221_X1 port map( B1 => n61846, B2 => n2285, C1 => n61843, C2 => 
                           n2401, A => n7913, ZN => n7904);
   U2914 : NOR4_X1 port map( A1 => n7804, A2 => n7805, A3 => n7806, A4 => n7807
                           , ZN => n7803);
   U2915 : OAI221_X1 port map( B1 => n61858, B2 => n2524, C1 => n61855, C2 => 
                           n2548, A => n7810, ZN => n7805);
   U2916 : OAI221_X1 port map( B1 => n61693, B2 => n2620, C1 => n61695, C2 => 
                           n2644, A => n7809, ZN => n7806);
   U2917 : OAI221_X1 port map( B1 => n61846, B2 => n2284, C1 => n61843, C2 => 
                           n2400, A => n7811, ZN => n7804);
   U2918 : NOR4_X1 port map( A1 => n7729, A2 => n7730, A3 => n7731, A4 => n7732
                           , ZN => n7728);
   U2919 : OAI221_X1 port map( B1 => n61858, B2 => n2523, C1 => n61855, C2 => 
                           n2547, A => n7735, ZN => n7730);
   U2920 : OAI221_X1 port map( B1 => n61693, B2 => n2619, C1 => n61695, C2 => 
                           n2643, A => n7734, ZN => n7731);
   U2921 : OAI221_X1 port map( B1 => n61846, B2 => n2283, C1 => n61843, C2 => 
                           n2399, A => n7736, ZN => n7729);
   U2922 : NOR4_X1 port map( A1 => n7654, A2 => n7655, A3 => n7656, A4 => n7657
                           , ZN => n7653);
   U2923 : OAI221_X1 port map( B1 => n61858, B2 => n2522, C1 => n61855, C2 => 
                           n2546, A => n7660, ZN => n7655);
   U2924 : OAI221_X1 port map( B1 => n61693, B2 => n2618, C1 => n61695, C2 => 
                           n2642, A => n7659, ZN => n7656);
   U2925 : OAI221_X1 port map( B1 => n61846, B2 => n2282, C1 => n61843, C2 => 
                           n2398, A => n7661, ZN => n7654);
   U2926 : NOR4_X1 port map( A1 => n7579, A2 => n7580, A3 => n7581, A4 => n7582
                           , ZN => n7578);
   U2927 : OAI221_X1 port map( B1 => n61858, B2 => n2521, C1 => n61855, C2 => 
                           n2545, A => n7585, ZN => n7580);
   U2928 : OAI221_X1 port map( B1 => n61693, B2 => n2617, C1 => n61695, C2 => 
                           n2641, A => n7584, ZN => n7581);
   U2929 : OAI221_X1 port map( B1 => n61846, B2 => n2281, C1 => n61843, C2 => 
                           n2397, A => n7586, ZN => n7579);
   U2930 : NOR4_X1 port map( A1 => n7504, A2 => n7505, A3 => n7506, A4 => n7507
                           , ZN => n7503);
   U2931 : OAI221_X1 port map( B1 => n61858, B2 => n2520, C1 => n61855, C2 => 
                           n2544, A => n7510, ZN => n7505);
   U2932 : OAI221_X1 port map( B1 => n61693, B2 => n2616, C1 => n61695, C2 => 
                           n2640, A => n7509, ZN => n7506);
   U2933 : OAI221_X1 port map( B1 => n61846, B2 => n2280, C1 => n61843, C2 => 
                           n2396, A => n7511, ZN => n7504);
   U2934 : NOR4_X1 port map( A1 => n7429, A2 => n7430, A3 => n7431, A4 => n7432
                           , ZN => n7428);
   U2935 : OAI221_X1 port map( B1 => n61858, B2 => n2519, C1 => n61855, C2 => 
                           n2543, A => n7435, ZN => n7430);
   U2936 : OAI221_X1 port map( B1 => n61693, B2 => n2615, C1 => n61695, C2 => 
                           n2639, A => n7434, ZN => n7431);
   U2937 : OAI221_X1 port map( B1 => n61846, B2 => n2279, C1 => n61843, C2 => 
                           n2395, A => n7436, ZN => n7429);
   U2938 : NOR4_X1 port map( A1 => n7354, A2 => n7355, A3 => n7356, A4 => n7357
                           , ZN => n7353);
   U2939 : OAI221_X1 port map( B1 => n61858, B2 => n2518, C1 => n61855, C2 => 
                           n2542, A => n7360, ZN => n7355);
   U2940 : OAI221_X1 port map( B1 => n61693, B2 => n2614, C1 => n61695, C2 => 
                           n2638, A => n7359, ZN => n7356);
   U2941 : OAI221_X1 port map( B1 => n61846, B2 => n2278, C1 => n61843, C2 => 
                           n2394, A => n7361, ZN => n7354);
   U2942 : NOR4_X1 port map( A1 => n7204, A2 => n7205, A3 => n7206, A4 => n7207
                           , ZN => n7203);
   U2943 : OAI221_X1 port map( B1 => n61858, B2 => n2516, C1 => n61855, C2 => 
                           n2540, A => n7210, ZN => n7205);
   U2944 : OAI221_X1 port map( B1 => n61693, B2 => n2612, C1 => n61695, C2 => 
                           n2636, A => n7209, ZN => n7206);
   U2945 : OAI221_X1 port map( B1 => n61846, B2 => n2276, C1 => n61843, C2 => 
                           n2392, A => n7211, ZN => n7204);
   U2946 : NOR4_X1 port map( A1 => n6979, A2 => n6980, A3 => n6981, A4 => n6982
                           , ZN => n6978);
   U2947 : OAI221_X1 port map( B1 => n61859, B2 => n2513, C1 => n61856, C2 => 
                           n2537, A => n6985, ZN => n6980);
   U2948 : OAI221_X1 port map( B1 => n6073, B2 => n2609, C1 => n61696, C2 => 
                           n2633, A => n6984, ZN => n6981);
   U2949 : OAI221_X1 port map( B1 => n61847, B2 => n2273, C1 => n61844, C2 => 
                           n2297, A => n6986, ZN => n6979);
   U2950 : NOR4_X1 port map( A1 => n14408, A2 => n14409, A3 => n14410, A4 => 
                           n14411, ZN => n14407);
   U2951 : OAI221_X1 port map( B1 => n2393, B2 => n61436, C1 => n2277, C2 => 
                           n61433, A => n14414, ZN => n14409);
   U2952 : OAI221_X1 port map( B1 => n2517, B2 => n61448, C1 => n2541, C2 => 
                           n61445, A => n14413, ZN => n14410);
   U2953 : OAI221_X1 port map( B1 => n2637, B2 => n61460, C1 => n2613, C2 => 
                           n61457, A => n14412, ZN => n14411);
   U2954 : NOR4_X1 port map( A1 => n9917, A2 => n9918, A3 => n9919, A4 => n9920
                           , ZN => n9916);
   U2955 : OAI221_X1 port map( B1 => n2392, B2 => n61436, C1 => n2276, C2 => 
                           n61433, A => n9923, ZN => n9918);
   U2956 : OAI221_X1 port map( B1 => n2516, B2 => n61448, C1 => n2540, C2 => 
                           n61445, A => n9922, ZN => n9919);
   U2957 : OAI221_X1 port map( B1 => n2636, B2 => n61460, C1 => n2612, C2 => 
                           n61457, A => n9921, ZN => n9920);
   U2958 : NOR4_X1 port map( A1 => n9842, A2 => n9843, A3 => n9844, A4 => n9845
                           , ZN => n9841);
   U2959 : OAI221_X1 port map( B1 => n2391, B2 => n61436, C1 => n2275, C2 => 
                           n61433, A => n9848, ZN => n9843);
   U2960 : OAI221_X1 port map( B1 => n2515, B2 => n61448, C1 => n2539, C2 => 
                           n61445, A => n9847, ZN => n9844);
   U2961 : OAI221_X1 port map( B1 => n2635, B2 => n61460, C1 => n2611, C2 => 
                           n61457, A => n9846, ZN => n9845);
   U2962 : NOR4_X1 port map( A1 => n9703, A2 => n9704, A3 => n9705, A4 => n9706
                           , ZN => n9702);
   U2963 : OAI221_X1 port map( B1 => n2298, B2 => n61436, C1 => n2274, C2 => 
                           n61433, A => n9709, ZN => n9704);
   U2964 : OAI221_X1 port map( B1 => n2514, B2 => n61448, C1 => n2538, C2 => 
                           n61445, A => n9708, ZN => n9705);
   U2965 : OAI221_X1 port map( B1 => n2634, B2 => n61460, C1 => n2610, C2 => 
                           n61457, A => n9707, ZN => n9706);
   U2966 : NOR4_X1 port map( A1 => n9628, A2 => n9629, A3 => n9630, A4 => n9631
                           , ZN => n9627);
   U2967 : OAI221_X1 port map( B1 => n2297, B2 => n61437, C1 => n2273, C2 => 
                           n61434, A => n9634, ZN => n9629);
   U2968 : OAI221_X1 port map( B1 => n2513, B2 => n61449, C1 => n2537, C2 => 
                           n61446, A => n9633, ZN => n9630);
   U2969 : OAI221_X1 port map( B1 => n2633, B2 => n61461, C1 => n2609, C2 => 
                           n61458, A => n9632, ZN => n9631);
   U2970 : NOR4_X1 port map( A1 => n9537, A2 => n9538, A3 => n9539, A4 => n9540
                           , ZN => n9536);
   U2971 : OAI221_X1 port map( B1 => n2296, B2 => n61437, C1 => n2272, C2 => 
                           n61434, A => n9543, ZN => n9538);
   U2972 : OAI221_X1 port map( B1 => n2512, B2 => n61449, C1 => n2536, C2 => 
                           n61446, A => n9542, ZN => n9539);
   U2973 : OAI221_X1 port map( B1 => n2632, B2 => n61461, C1 => n2608, C2 => 
                           n61458, A => n9541, ZN => n9540);
   U2974 : NOR4_X1 port map( A1 => n9462, A2 => n9463, A3 => n9464, A4 => n9465
                           , ZN => n9461);
   U2975 : OAI221_X1 port map( B1 => n2295, B2 => n61437, C1 => n2271, C2 => 
                           n61434, A => n9468, ZN => n9463);
   U2976 : OAI221_X1 port map( B1 => n2511, B2 => n61449, C1 => n2535, C2 => 
                           n61446, A => n9467, ZN => n9464);
   U2977 : OAI221_X1 port map( B1 => n2631, B2 => n61461, C1 => n2607, C2 => 
                           n61458, A => n9466, ZN => n9465);
   U2978 : NOR4_X1 port map( A1 => n9387, A2 => n9388, A3 => n9389, A4 => n9390
                           , ZN => n9386);
   U2979 : OAI221_X1 port map( B1 => n2294, B2 => n61437, C1 => n2234, C2 => 
                           n61434, A => n9393, ZN => n9388);
   U2980 : OAI221_X1 port map( B1 => n2482, B2 => n61449, C1 => n2534, C2 => 
                           n61446, A => n9392, ZN => n9389);
   U2981 : OAI221_X1 port map( B1 => n2630, B2 => n61461, C1 => n2606, C2 => 
                           n61458, A => n9391, ZN => n9390);
   U2982 : NOR4_X1 port map( A1 => n9248, A2 => n9249, A3 => n9250, A4 => n9251
                           , ZN => n9247);
   U2983 : OAI221_X1 port map( B1 => n2293, B2 => n61437, C1 => n2233, C2 => 
                           n61434, A => n9254, ZN => n9249);
   U2984 : OAI221_X1 port map( B1 => n2481, B2 => n61449, C1 => n2533, C2 => 
                           n61446, A => n9253, ZN => n9250);
   U2985 : OAI221_X1 port map( B1 => n2629, B2 => n61461, C1 => n2605, C2 => 
                           n61458, A => n9252, ZN => n9251);
   U2986 : NOR4_X1 port map( A1 => n9173, A2 => n9174, A3 => n9175, A4 => n9176
                           , ZN => n9172);
   U2987 : OAI221_X1 port map( B1 => n2292, B2 => n61437, C1 => n2232, C2 => 
                           n61434, A => n9179, ZN => n9174);
   U2988 : OAI221_X1 port map( B1 => n2480, B2 => n61449, C1 => n2532, C2 => 
                           n61446, A => n9178, ZN => n9175);
   U2989 : OAI221_X1 port map( B1 => n2628, B2 => n61461, C1 => n2604, C2 => 
                           n61458, A => n9177, ZN => n9176);
   U2990 : NOR4_X1 port map( A1 => n9098, A2 => n9099, A3 => n9100, A4 => n9101
                           , ZN => n9097);
   U2991 : OAI221_X1 port map( B1 => n2291, B2 => n61437, C1 => n2231, C2 => 
                           n61434, A => n9104, ZN => n9099);
   U2992 : OAI221_X1 port map( B1 => n2479, B2 => n61449, C1 => n2531, C2 => 
                           n61446, A => n9103, ZN => n9100);
   U2993 : OAI221_X1 port map( B1 => n2627, B2 => n61461, C1 => n2603, C2 => 
                           n61458, A => n9102, ZN => n9101);
   U2994 : NOR4_X1 port map( A1 => n9023, A2 => n9024, A3 => n9025, A4 => n9026
                           , ZN => n9022);
   U2995 : OAI221_X1 port map( B1 => n2290, B2 => n61437, C1 => n2230, C2 => 
                           n61434, A => n9029, ZN => n9024);
   U2996 : OAI221_X1 port map( B1 => n2478, B2 => n61449, C1 => n2530, C2 => 
                           n61446, A => n9028, ZN => n9025);
   U2997 : OAI221_X1 port map( B1 => n2626, B2 => n61461, C1 => n2602, C2 => 
                           n61458, A => n9027, ZN => n9026);
   U2998 : NOR4_X1 port map( A1 => n8948, A2 => n8949, A3 => n8950, A4 => n8951
                           , ZN => n8947);
   U2999 : OAI221_X1 port map( B1 => n2289, B2 => n61437, C1 => n2229, C2 => 
                           n61434, A => n8954, ZN => n8949);
   U3000 : OAI221_X1 port map( B1 => n2477, B2 => n61449, C1 => n2529, C2 => 
                           n61446, A => n8953, ZN => n8950);
   U3001 : OAI221_X1 port map( B1 => n2625, B2 => n61461, C1 => n2601, C2 => 
                           n61458, A => n8952, ZN => n8951);
   U3002 : NOR4_X1 port map( A1 => n8873, A2 => n8874, A3 => n8875, A4 => n8876
                           , ZN => n8872);
   U3003 : OAI221_X1 port map( B1 => n2288, B2 => n61437, C1 => n2228, C2 => 
                           n61434, A => n8879, ZN => n8874);
   U3004 : OAI221_X1 port map( B1 => n2476, B2 => n61449, C1 => n2528, C2 => 
                           n61446, A => n8878, ZN => n8875);
   U3005 : OAI221_X1 port map( B1 => n2624, B2 => n61461, C1 => n2600, C2 => 
                           n61458, A => n8877, ZN => n8876);
   U3006 : NOR4_X1 port map( A1 => n8798, A2 => n8799, A3 => n8800, A4 => n8801
                           , ZN => n8797);
   U3007 : OAI221_X1 port map( B1 => n2287, B2 => n61437, C1 => n2227, C2 => 
                           n61434, A => n8804, ZN => n8799);
   U3008 : OAI221_X1 port map( B1 => n2475, B2 => n61449, C1 => n2527, C2 => 
                           n61446, A => n8803, ZN => n8800);
   U3009 : OAI221_X1 port map( B1 => n2623, B2 => n61461, C1 => n2599, C2 => 
                           n61458, A => n8802, ZN => n8801);
   U3010 : NOR4_X1 port map( A1 => n8723, A2 => n8724, A3 => n8725, A4 => n8726
                           , ZN => n8722);
   U3011 : OAI221_X1 port map( B1 => n2286, B2 => n61437, C1 => n2226, C2 => 
                           n61434, A => n8729, ZN => n8724);
   U3012 : OAI221_X1 port map( B1 => n2474, B2 => n61449, C1 => n2526, C2 => 
                           n61446, A => n8728, ZN => n8725);
   U3013 : OAI221_X1 port map( B1 => n2622, B2 => n61461, C1 => n2598, C2 => 
                           n61458, A => n8727, ZN => n8726);
   U3014 : NOR4_X1 port map( A1 => n15031, A2 => n15032, A3 => n15033, A4 => 
                           n15034, ZN => n15030);
   U3015 : OAI221_X1 port map( B1 => n2401, B2 => n61436, C1 => n2285, C2 => 
                           n61433, A => n15039, ZN => n15032);
   U3016 : OAI221_X1 port map( B1 => n2525, B2 => n61448, C1 => n2549, C2 => 
                           n61445, A => n15037, ZN => n15033);
   U3017 : OAI221_X1 port map( B1 => n2652, B2 => n61460, C1 => n2621, C2 => 
                           n61457, A => n15035, ZN => n15034);
   U3018 : NOR4_X1 port map( A1 => n14933, A2 => n14934, A3 => n14935, A4 => 
                           n14936, ZN => n14932);
   U3019 : OAI221_X1 port map( B1 => n2400, B2 => n61436, C1 => n2284, C2 => 
                           n61433, A => n14939, ZN => n14934);
   U3020 : OAI221_X1 port map( B1 => n2524, B2 => n61448, C1 => n2548, C2 => 
                           n61445, A => n14938, ZN => n14935);
   U3021 : OAI221_X1 port map( B1 => n2644, B2 => n61460, C1 => n2620, C2 => 
                           n61457, A => n14937, ZN => n14936);
   U3022 : NOR4_X1 port map( A1 => n14858, A2 => n14859, A3 => n14860, A4 => 
                           n14861, ZN => n14857);
   U3023 : OAI221_X1 port map( B1 => n2399, B2 => n61436, C1 => n2283, C2 => 
                           n61433, A => n14864, ZN => n14859);
   U3024 : OAI221_X1 port map( B1 => n2523, B2 => n61448, C1 => n2547, C2 => 
                           n61445, A => n14863, ZN => n14860);
   U3025 : OAI221_X1 port map( B1 => n2643, B2 => n61460, C1 => n2619, C2 => 
                           n61457, A => n14862, ZN => n14861);
   U3026 : NOR4_X1 port map( A1 => n14783, A2 => n14784, A3 => n14785, A4 => 
                           n14786, ZN => n14782);
   U3027 : OAI221_X1 port map( B1 => n2398, B2 => n61436, C1 => n2282, C2 => 
                           n61433, A => n14789, ZN => n14784);
   U3028 : OAI221_X1 port map( B1 => n2522, B2 => n61448, C1 => n2546, C2 => 
                           n61445, A => n14788, ZN => n14785);
   U3029 : OAI221_X1 port map( B1 => n2642, B2 => n61460, C1 => n2618, C2 => 
                           n61457, A => n14787, ZN => n14786);
   U3030 : NOR4_X1 port map( A1 => n14708, A2 => n14709, A3 => n14710, A4 => 
                           n14711, ZN => n14707);
   U3031 : OAI221_X1 port map( B1 => n2397, B2 => n61436, C1 => n2281, C2 => 
                           n61433, A => n14714, ZN => n14709);
   U3032 : OAI221_X1 port map( B1 => n2521, B2 => n61448, C1 => n2545, C2 => 
                           n61445, A => n14713, ZN => n14710);
   U3033 : OAI221_X1 port map( B1 => n2641, B2 => n61460, C1 => n2617, C2 => 
                           n61457, A => n14712, ZN => n14711);
   U3034 : NOR4_X1 port map( A1 => n14633, A2 => n14634, A3 => n14635, A4 => 
                           n14636, ZN => n14632);
   U3035 : OAI221_X1 port map( B1 => n2396, B2 => n61436, C1 => n2280, C2 => 
                           n61433, A => n14639, ZN => n14634);
   U3036 : OAI221_X1 port map( B1 => n2520, B2 => n61448, C1 => n2544, C2 => 
                           n61445, A => n14638, ZN => n14635);
   U3037 : OAI221_X1 port map( B1 => n2640, B2 => n61460, C1 => n2616, C2 => 
                           n61457, A => n14637, ZN => n14636);
   U3038 : NOR4_X1 port map( A1 => n14558, A2 => n14559, A3 => n14560, A4 => 
                           n14561, ZN => n14557);
   U3039 : OAI221_X1 port map( B1 => n2395, B2 => n61436, C1 => n2279, C2 => 
                           n61433, A => n14564, ZN => n14559);
   U3040 : OAI221_X1 port map( B1 => n2519, B2 => n61448, C1 => n2543, C2 => 
                           n61445, A => n14563, ZN => n14560);
   U3041 : OAI221_X1 port map( B1 => n2639, B2 => n61460, C1 => n2615, C2 => 
                           n61457, A => n14562, ZN => n14561);
   U3042 : NOR4_X1 port map( A1 => n14483, A2 => n14484, A3 => n14485, A4 => 
                           n14486, ZN => n14482);
   U3043 : OAI221_X1 port map( B1 => n2394, B2 => n61436, C1 => n2278, C2 => 
                           n61433, A => n14489, ZN => n14484);
   U3044 : OAI221_X1 port map( B1 => n2518, B2 => n61448, C1 => n2542, C2 => 
                           n61445, A => n14488, ZN => n14485);
   U3045 : OAI221_X1 port map( B1 => n2638, B2 => n61460, C1 => n2614, C2 => 
                           n61457, A => n14487, ZN => n14486);
   U3046 : NOR4_X1 port map( A1 => n8612, A2 => n8613, A3 => n8614, A4 => n8615
                           , ZN => n8611);
   U3047 : OAI221_X1 port map( B1 => n4139, B2 => n61642, C1 => n4147, C2 => 
                           n61639, A => n8618, ZN => n8613);
   U3048 : OAI221_X1 port map( B1 => n4155, B2 => n61654, C1 => n4163, C2 => 
                           n61651, A => n8617, ZN => n8614);
   U3049 : OAI221_X1 port map( B1 => n478, B2 => n61666, C1 => n486, C2 => 
                           n61663, A => n8616, ZN => n8615);
   U3050 : NOR4_X1 port map( A1 => n8648, A2 => n8649, A3 => n8650, A4 => n8651
                           , ZN => n8647);
   U3051 : OAI221_X1 port map( B1 => n4059, B2 => n61438, C1 => n4051, C2 => 
                           n61435, A => n8654, ZN => n8649);
   U3052 : OAI221_X1 port map( B1 => n324, B2 => n61450, C1 => n332, C2 => 
                           n61447, A => n8653, ZN => n8650);
   U3053 : OAI221_X1 port map( B1 => n4075, B2 => n61462, C1 => n4067, C2 => 
                           n61459, A => n8652, ZN => n8651);
   U3054 : NOR4_X1 port map( A1 => n8537, A2 => n8538, A3 => n8539, A4 => n8540
                           , ZN => n8536);
   U3055 : OAI221_X1 port map( B1 => n4138, B2 => n61642, C1 => n4146, C2 => 
                           n61639, A => n8543, ZN => n8538);
   U3056 : OAI221_X1 port map( B1 => n4154, B2 => n61654, C1 => n4162, C2 => 
                           n61651, A => n8542, ZN => n8539);
   U3057 : OAI221_X1 port map( B1 => n477, B2 => n61666, C1 => n485, C2 => 
                           n61663, A => n8541, ZN => n8540);
   U3058 : NOR4_X1 port map( A1 => n8573, A2 => n8574, A3 => n8575, A4 => n8576
                           , ZN => n8572);
   U3059 : OAI221_X1 port map( B1 => n4058, B2 => n61438, C1 => n4050, C2 => 
                           n61435, A => n8579, ZN => n8574);
   U3060 : OAI221_X1 port map( B1 => n323, B2 => n61450, C1 => n331, C2 => 
                           n61447, A => n8578, ZN => n8575);
   U3061 : OAI221_X1 port map( B1 => n4074, B2 => n61462, C1 => n4066, C2 => 
                           n61459, A => n8577, ZN => n8576);
   U3062 : NOR4_X1 port map( A1 => n8462, A2 => n8463, A3 => n8464, A4 => n8465
                           , ZN => n8461);
   U3063 : OAI221_X1 port map( B1 => n4137, B2 => n61642, C1 => n4145, C2 => 
                           n61639, A => n8468, ZN => n8463);
   U3064 : OAI221_X1 port map( B1 => n4153, B2 => n61654, C1 => n4161, C2 => 
                           n61651, A => n8467, ZN => n8464);
   U3065 : OAI221_X1 port map( B1 => n476, B2 => n61666, C1 => n484, C2 => 
                           n61663, A => n8466, ZN => n8465);
   U3066 : NOR4_X1 port map( A1 => n8498, A2 => n8499, A3 => n8500, A4 => n8501
                           , ZN => n8497);
   U3067 : OAI221_X1 port map( B1 => n4057, B2 => n61438, C1 => n4049, C2 => 
                           n61435, A => n8504, ZN => n8499);
   U3068 : OAI221_X1 port map( B1 => n322, B2 => n61450, C1 => n330, C2 => 
                           n61447, A => n8503, ZN => n8500);
   U3069 : OAI221_X1 port map( B1 => n4073, B2 => n61462, C1 => n4065, C2 => 
                           n61459, A => n8502, ZN => n8501);
   U3070 : NOR4_X1 port map( A1 => n8387, A2 => n8388, A3 => n8389, A4 => n8390
                           , ZN => n8386);
   U3071 : OAI221_X1 port map( B1 => n4136, B2 => n61642, C1 => n4144, C2 => 
                           n61639, A => n8393, ZN => n8388);
   U3072 : OAI221_X1 port map( B1 => n4152, B2 => n61654, C1 => n4160, C2 => 
                           n61651, A => n8392, ZN => n8389);
   U3073 : OAI221_X1 port map( B1 => n473, B2 => n61666, C1 => n483, C2 => 
                           n61663, A => n8391, ZN => n8390);
   U3074 : NOR4_X1 port map( A1 => n8423, A2 => n8424, A3 => n8425, A4 => n8426
                           , ZN => n8422);
   U3075 : OAI221_X1 port map( B1 => n4056, B2 => n61438, C1 => n4048, C2 => 
                           n61435, A => n8429, ZN => n8424);
   U3076 : OAI221_X1 port map( B1 => n321, B2 => n61450, C1 => n329, C2 => 
                           n61447, A => n8428, ZN => n8425);
   U3077 : OAI221_X1 port map( B1 => n4072, B2 => n61462, C1 => n4064, C2 => 
                           n61459, A => n8427, ZN => n8426);
   U3078 : NOR4_X1 port map( A1 => n8312, A2 => n8313, A3 => n8314, A4 => n8315
                           , ZN => n8311);
   U3079 : OAI221_X1 port map( B1 => n4135, B2 => n61642, C1 => n4143, C2 => 
                           n61639, A => n8318, ZN => n8313);
   U3080 : OAI221_X1 port map( B1 => n4151, B2 => n61654, C1 => n4159, C2 => 
                           n61651, A => n8317, ZN => n8314);
   U3081 : OAI221_X1 port map( B1 => n472, B2 => n61666, C1 => n482, C2 => 
                           n61663, A => n8316, ZN => n8315);
   U3082 : NOR4_X1 port map( A1 => n8348, A2 => n8349, A3 => n8350, A4 => n8351
                           , ZN => n8347);
   U3083 : OAI221_X1 port map( B1 => n4055, B2 => n61438, C1 => n4047, C2 => 
                           n61435, A => n8354, ZN => n8349);
   U3084 : OAI221_X1 port map( B1 => n320, B2 => n61450, C1 => n328, C2 => 
                           n61447, A => n8353, ZN => n8350);
   U3085 : OAI221_X1 port map( B1 => n4071, B2 => n61462, C1 => n4063, C2 => 
                           n61459, A => n8352, ZN => n8351);
   U3086 : NOR4_X1 port map( A1 => n8237, A2 => n8238, A3 => n8239, A4 => n8240
                           , ZN => n8236);
   U3087 : OAI221_X1 port map( B1 => n4134, B2 => n61642, C1 => n4142, C2 => 
                           n61639, A => n8243, ZN => n8238);
   U3088 : OAI221_X1 port map( B1 => n4150, B2 => n61654, C1 => n4158, C2 => 
                           n61651, A => n8242, ZN => n8239);
   U3089 : OAI221_X1 port map( B1 => n471, B2 => n61666, C1 => n481, C2 => 
                           n61663, A => n8241, ZN => n8240);
   U3090 : NOR4_X1 port map( A1 => n8273, A2 => n8274, A3 => n8275, A4 => n8276
                           , ZN => n8272);
   U3091 : OAI221_X1 port map( B1 => n4054, B2 => n61438, C1 => n4046, C2 => 
                           n61435, A => n8279, ZN => n8274);
   U3092 : OAI221_X1 port map( B1 => n319, B2 => n61450, C1 => n327, C2 => 
                           n61447, A => n8278, ZN => n8275);
   U3093 : OAI221_X1 port map( B1 => n4070, B2 => n61462, C1 => n4062, C2 => 
                           n61459, A => n8277, ZN => n8276);
   U3094 : NOR4_X1 port map( A1 => n8162, A2 => n8163, A3 => n8164, A4 => n8165
                           , ZN => n8161);
   U3095 : OAI221_X1 port map( B1 => n4133, B2 => n61642, C1 => n4141, C2 => 
                           n61639, A => n8168, ZN => n8163);
   U3096 : OAI221_X1 port map( B1 => n4149, B2 => n61654, C1 => n4157, C2 => 
                           n61651, A => n8167, ZN => n8164);
   U3097 : OAI221_X1 port map( B1 => n470, B2 => n61666, C1 => n480, C2 => 
                           n61663, A => n8166, ZN => n8165);
   U3098 : NOR4_X1 port map( A1 => n8198, A2 => n8199, A3 => n8200, A4 => n8201
                           , ZN => n8197);
   U3099 : OAI221_X1 port map( B1 => n4053, B2 => n61438, C1 => n4045, C2 => 
                           n61435, A => n8204, ZN => n8199);
   U3100 : OAI221_X1 port map( B1 => n318, B2 => n61450, C1 => n326, C2 => 
                           n61447, A => n8203, ZN => n8200);
   U3101 : OAI221_X1 port map( B1 => n4069, B2 => n61462, C1 => n4061, C2 => 
                           n61459, A => n8202, ZN => n8201);
   U3102 : NOR4_X1 port map( A1 => n7951, A2 => n7952, A3 => n7953, A4 => n7954
                           , ZN => n7950);
   U3103 : OAI221_X1 port map( B1 => n4132, B2 => n61642, C1 => n4140, C2 => 
                           n61639, A => n7967, ZN => n7952);
   U3104 : OAI221_X1 port map( B1 => n4148, B2 => n61654, C1 => n4156, C2 => 
                           n61651, A => n7962, ZN => n7953);
   U3105 : OAI221_X1 port map( B1 => n469, B2 => n61666, C1 => n479, C2 => 
                           n61663, A => n7957, ZN => n7954);
   U3106 : NOR4_X1 port map( A1 => n8055, A2 => n8056, A3 => n8057, A4 => n8058
                           , ZN => n8054);
   U3107 : OAI221_X1 port map( B1 => n4052, B2 => n61438, C1 => n4044, C2 => 
                           n61435, A => n8071, ZN => n8056);
   U3108 : OAI221_X1 port map( B1 => n317, B2 => n61450, C1 => n325, C2 => 
                           n61447, A => n8066, ZN => n8057);
   U3109 : OAI221_X1 port map( B1 => n4068, B2 => n61462, C1 => n4060, C2 => 
                           n61459, A => n8061, ZN => n8058);
   U3110 : OAI21_X1 port map( B1 => n15270, B2 => n15109, A => n62187, ZN => 
                           n5362);
   U3111 : NOR4_X1 port map( A1 => n14416, A2 => n14417, A3 => n14418, A4 => 
                           n14419, ZN => n14406);
   U3112 : OAI221_X1 port map( B1 => n1917, B2 => n61397, C1 => n1941, C2 => 
                           n61394, A => n14421, ZN => n14418);
   U3113 : OAI221_X1 port map( B1 => n2037, B2 => n61409, C1 => n1989, C2 => 
                           n61406, A => n14420, ZN => n14419);
   U3114 : OAI221_X1 port map( B1 => n1845, B2 => n61385, C1 => n1821, C2 => 
                           n61382, A => n14422, ZN => n14417);
   U3115 : NOR4_X1 port map( A1 => n14341, A2 => n14342, A3 => n14343, A4 => 
                           n14344, ZN => n9915);
   U3116 : OAI221_X1 port map( B1 => n1916, B2 => n61397, C1 => n1940, C2 => 
                           n61394, A => n14346, ZN => n14343);
   U3117 : OAI221_X1 port map( B1 => n2036, B2 => n61409, C1 => n1988, C2 => 
                           n61406, A => n14345, ZN => n14344);
   U3118 : OAI221_X1 port map( B1 => n1844, B2 => n61385, C1 => n1820, C2 => 
                           n61382, A => n14347, ZN => n14342);
   U3119 : NOR4_X1 port map( A1 => n9850, A2 => n9851, A3 => n9852, A4 => n9853
                           , ZN => n9840);
   U3120 : OAI221_X1 port map( B1 => n1915, B2 => n61397, C1 => n1939, C2 => 
                           n61394, A => n9855, ZN => n9852);
   U3121 : OAI221_X1 port map( B1 => n2035, B2 => n61409, C1 => n1987, C2 => 
                           n61406, A => n9854, ZN => n9853);
   U3122 : OAI221_X1 port map( B1 => n1843, B2 => n61385, C1 => n1819, C2 => 
                           n61382, A => n9856, ZN => n9851);
   U3123 : NOR4_X1 port map( A1 => n9711, A2 => n9712, A3 => n9713, A4 => n9714
                           , ZN => n9701);
   U3124 : OAI221_X1 port map( B1 => n1914, B2 => n61397, C1 => n1938, C2 => 
                           n61394, A => n9716, ZN => n9713);
   U3125 : OAI221_X1 port map( B1 => n2034, B2 => n61409, C1 => n1986, C2 => 
                           n61406, A => n9715, ZN => n9714);
   U3126 : OAI221_X1 port map( B1 => n1842, B2 => n61385, C1 => n1818, C2 => 
                           n61382, A => n9717, ZN => n9712);
   U3127 : NOR4_X1 port map( A1 => n9636, A2 => n9637, A3 => n9638, A4 => n9639
                           , ZN => n9626);
   U3128 : OAI221_X1 port map( B1 => n1913, B2 => n61398, C1 => n1937, C2 => 
                           n61395, A => n9641, ZN => n9638);
   U3129 : OAI221_X1 port map( B1 => n2033, B2 => n61410, C1 => n1985, C2 => 
                           n61407, A => n9640, ZN => n9639);
   U3130 : OAI221_X1 port map( B1 => n1841, B2 => n61386, C1 => n1817, C2 => 
                           n61383, A => n9642, ZN => n9637);
   U3131 : NOR4_X1 port map( A1 => n9545, A2 => n9546, A3 => n9547, A4 => n9548
                           , ZN => n9535);
   U3132 : OAI221_X1 port map( B1 => n1912, B2 => n61398, C1 => n1936, C2 => 
                           n61395, A => n9550, ZN => n9547);
   U3133 : OAI221_X1 port map( B1 => n2032, B2 => n61410, C1 => n1984, C2 => 
                           n61407, A => n9549, ZN => n9548);
   U3134 : OAI221_X1 port map( B1 => n1840, B2 => n61386, C1 => n1816, C2 => 
                           n61383, A => n9551, ZN => n9546);
   U3135 : NOR4_X1 port map( A1 => n9470, A2 => n9471, A3 => n9472, A4 => n9473
                           , ZN => n9460);
   U3136 : OAI221_X1 port map( B1 => n1911, B2 => n61398, C1 => n1935, C2 => 
                           n61395, A => n9475, ZN => n9472);
   U3137 : OAI221_X1 port map( B1 => n2031, B2 => n61410, C1 => n1983, C2 => 
                           n61407, A => n9474, ZN => n9473);
   U3138 : OAI221_X1 port map( B1 => n1839, B2 => n61386, C1 => n1815, C2 => 
                           n61383, A => n9476, ZN => n9471);
   U3139 : NOR4_X1 port map( A1 => n9395, A2 => n9396, A3 => n9397, A4 => n9398
                           , ZN => n9385);
   U3140 : OAI221_X1 port map( B1 => n1910, B2 => n61398, C1 => n1934, C2 => 
                           n61395, A => n9400, ZN => n9397);
   U3141 : OAI221_X1 port map( B1 => n2030, B2 => n61410, C1 => n1982, C2 => 
                           n61407, A => n9399, ZN => n9398);
   U3142 : OAI221_X1 port map( B1 => n1838, B2 => n61386, C1 => n1814, C2 => 
                           n61383, A => n9401, ZN => n9396);
   U3143 : NOR4_X1 port map( A1 => n9256, A2 => n9257, A3 => n9258, A4 => n9259
                           , ZN => n9246);
   U3144 : OAI221_X1 port map( B1 => n1909, B2 => n61398, C1 => n1933, C2 => 
                           n61395, A => n9261, ZN => n9258);
   U3145 : OAI221_X1 port map( B1 => n2029, B2 => n61410, C1 => n1981, C2 => 
                           n61407, A => n9260, ZN => n9259);
   U3146 : OAI221_X1 port map( B1 => n1837, B2 => n61386, C1 => n1813, C2 => 
                           n61383, A => n9262, ZN => n9257);
   U3147 : NOR4_X1 port map( A1 => n14641, A2 => n14642, A3 => n14643, A4 => 
                           n14644, ZN => n14631);
   U3148 : OAI221_X1 port map( B1 => n1920, B2 => n61397, C1 => n1944, C2 => 
                           n61394, A => n14646, ZN => n14643);
   U3149 : OAI221_X1 port map( B1 => n2040, B2 => n61409, C1 => n1992, C2 => 
                           n61406, A => n14645, ZN => n14644);
   U3150 : OAI221_X1 port map( B1 => n1848, B2 => n61385, C1 => n1824, C2 => 
                           n61382, A => n14647, ZN => n14642);
   U3151 : NOR4_X1 port map( A1 => n14566, A2 => n14567, A3 => n14568, A4 => 
                           n14569, ZN => n14556);
   U3152 : OAI221_X1 port map( B1 => n1919, B2 => n61397, C1 => n1943, C2 => 
                           n61394, A => n14571, ZN => n14568);
   U3153 : OAI221_X1 port map( B1 => n2039, B2 => n61409, C1 => n1991, C2 => 
                           n61406, A => n14570, ZN => n14569);
   U3154 : OAI221_X1 port map( B1 => n1847, B2 => n61385, C1 => n1823, C2 => 
                           n61382, A => n14572, ZN => n14567);
   U3155 : NOR4_X1 port map( A1 => n14491, A2 => n14492, A3 => n14493, A4 => 
                           n14494, ZN => n14481);
   U3156 : OAI221_X1 port map( B1 => n1918, B2 => n61397, C1 => n1942, C2 => 
                           n61394, A => n14496, ZN => n14493);
   U3157 : OAI221_X1 port map( B1 => n2038, B2 => n61409, C1 => n1990, C2 => 
                           n61406, A => n14495, ZN => n14494);
   U3158 : OAI221_X1 port map( B1 => n1846, B2 => n61385, C1 => n1822, C2 => 
                           n61382, A => n14497, ZN => n14492);
   U3159 : NOR4_X1 port map( A1 => n8656, A2 => n8657, A3 => n8658, A4 => n8659
                           , ZN => n8646);
   U3160 : OAI221_X1 port map( B1 => n4019, B2 => n61399, C1 => n4027, C2 => 
                           n61396, A => n8661, ZN => n8658);
   U3161 : OAI221_X1 port map( B1 => n260, B2 => n61411, C1 => n252, C2 => 
                           n61408, A => n8660, ZN => n8659);
   U3162 : OAI221_X1 port map( B1 => n159, B2 => n61387, C1 => n151, C2 => 
                           n61384, A => n8662, ZN => n8657);
   U3163 : NOR4_X1 port map( A1 => n8581, A2 => n8582, A3 => n8583, A4 => n8584
                           , ZN => n8571);
   U3164 : OAI221_X1 port map( B1 => n4018, B2 => n61399, C1 => n4026, C2 => 
                           n61396, A => n8586, ZN => n8583);
   U3165 : OAI221_X1 port map( B1 => n259, B2 => n61411, C1 => n251, C2 => 
                           n61408, A => n8585, ZN => n8584);
   U3166 : OAI221_X1 port map( B1 => n158, B2 => n61387, C1 => n150, C2 => 
                           n61384, A => n8587, ZN => n8582);
   U3167 : NOR4_X1 port map( A1 => n8506, A2 => n8507, A3 => n8508, A4 => n8509
                           , ZN => n8496);
   U3168 : OAI221_X1 port map( B1 => n4017, B2 => n61399, C1 => n4025, C2 => 
                           n61396, A => n8511, ZN => n8508);
   U3169 : OAI221_X1 port map( B1 => n258, B2 => n61411, C1 => n250, C2 => 
                           n61408, A => n8510, ZN => n8509);
   U3170 : OAI221_X1 port map( B1 => n157, B2 => n61387, C1 => n149, C2 => 
                           n61384, A => n8512, ZN => n8507);
   U3171 : NOR4_X1 port map( A1 => n8431, A2 => n8432, A3 => n8433, A4 => n8434
                           , ZN => n8421);
   U3172 : OAI221_X1 port map( B1 => n4016, B2 => n61399, C1 => n4024, C2 => 
                           n61396, A => n8436, ZN => n8433);
   U3173 : OAI221_X1 port map( B1 => n257, B2 => n61411, C1 => n249, C2 => 
                           n61408, A => n8435, ZN => n8434);
   U3174 : OAI221_X1 port map( B1 => n156, B2 => n61387, C1 => n148, C2 => 
                           n61384, A => n8437, ZN => n8432);
   U3175 : NOR4_X1 port map( A1 => n8356, A2 => n8357, A3 => n8358, A4 => n8359
                           , ZN => n8346);
   U3176 : OAI221_X1 port map( B1 => n4015, B2 => n61399, C1 => n4023, C2 => 
                           n61396, A => n8361, ZN => n8358);
   U3177 : OAI221_X1 port map( B1 => n256, B2 => n61411, C1 => n248, C2 => 
                           n61408, A => n8360, ZN => n8359);
   U3178 : OAI221_X1 port map( B1 => n155, B2 => n61387, C1 => n147, C2 => 
                           n61384, A => n8362, ZN => n8357);
   U3179 : NOR4_X1 port map( A1 => n8281, A2 => n8282, A3 => n8283, A4 => n8284
                           , ZN => n8271);
   U3180 : OAI221_X1 port map( B1 => n4014, B2 => n61399, C1 => n4022, C2 => 
                           n61396, A => n8286, ZN => n8283);
   U3181 : OAI221_X1 port map( B1 => n255, B2 => n61411, C1 => n247, C2 => 
                           n61408, A => n8285, ZN => n8284);
   U3182 : OAI221_X1 port map( B1 => n154, B2 => n61387, C1 => n146, C2 => 
                           n61384, A => n8287, ZN => n8282);
   U3183 : NOR4_X1 port map( A1 => n8206, A2 => n8207, A3 => n8208, A4 => n8209
                           , ZN => n8196);
   U3184 : OAI221_X1 port map( B1 => n4013, B2 => n61399, C1 => n4021, C2 => 
                           n61396, A => n8211, ZN => n8208);
   U3185 : OAI221_X1 port map( B1 => n254, B2 => n61411, C1 => n246, C2 => 
                           n61408, A => n8210, ZN => n8209);
   U3186 : OAI221_X1 port map( B1 => n153, B2 => n61387, C1 => n145, C2 => 
                           n61384, A => n8212, ZN => n8207);
   U3187 : NOR4_X1 port map( A1 => n8080, A2 => n8081, A3 => n8082, A4 => n8083
                           , ZN => n8053);
   U3188 : OAI221_X1 port map( B1 => n4012, B2 => n61399, C1 => n4020, C2 => 
                           n61396, A => n8091, ZN => n8082);
   U3189 : OAI221_X1 port map( B1 => n253, B2 => n61411, C1 => n245, C2 => 
                           n61408, A => n8086, ZN => n8083);
   U3190 : OAI221_X1 port map( B1 => n152, B2 => n61387, C1 => n144, C2 => 
                           n61384, A => n8096, ZN => n8081);
   U3191 : NOR4_X1 port map( A1 => n6093, A2 => n6094, A3 => n6095, A4 => n6096
                           , ZN => n6064);
   U3192 : OAI221_X1 port map( B1 => n61798, B2 => n1154, C1 => n61797, C2 => 
                           n1162, A => n6099, ZN => n6094);
   U3193 : OAI221_X1 port map( B1 => n5516, B2 => n1170, C1 => n5517, C2 => 
                           n1178, A => n6098, ZN => n6095);
   U3194 : OAI221_X1 port map( B1 => n61818, B2 => n1186, C1 => n61815, C2 => 
                           n1194, A => n6097, ZN => n6096);
   U3195 : NOR4_X1 port map( A1 => n5989, A2 => n5990, A3 => n5991, A4 => n5992
                           , ZN => n5970);
   U3196 : OAI221_X1 port map( B1 => n61798, B2 => n1153, C1 => n61797, C2 => 
                           n1161, A => n5995, ZN => n5990);
   U3197 : OAI221_X1 port map( B1 => n5516, B2 => n1169, C1 => n5517, C2 => 
                           n1177, A => n5994, ZN => n5991);
   U3198 : OAI221_X1 port map( B1 => n61818, B2 => n1185, C1 => n61815, C2 => 
                           n1193, A => n5993, ZN => n5992);
   U3199 : NOR4_X1 port map( A1 => n5914, A2 => n5915, A3 => n5916, A4 => n5917
                           , ZN => n5895);
   U3200 : OAI221_X1 port map( B1 => n61798, B2 => n1152, C1 => n61797, C2 => 
                           n1160, A => n5920, ZN => n5915);
   U3201 : OAI221_X1 port map( B1 => n5516, B2 => n1168, C1 => n5517, C2 => 
                           n1176, A => n5919, ZN => n5916);
   U3202 : OAI221_X1 port map( B1 => n61818, B2 => n1184, C1 => n61815, C2 => 
                           n1192, A => n5918, ZN => n5917);
   U3203 : NOR4_X1 port map( A1 => n5839, A2 => n5840, A3 => n5841, A4 => n5842
                           , ZN => n5820);
   U3204 : OAI221_X1 port map( B1 => n61798, B2 => n1151, C1 => n61797, C2 => 
                           n1159, A => n5845, ZN => n5840);
   U3205 : OAI221_X1 port map( B1 => n5516, B2 => n1167, C1 => n5517, C2 => 
                           n1175, A => n5844, ZN => n5841);
   U3206 : OAI221_X1 port map( B1 => n61818, B2 => n1183, C1 => n61815, C2 => 
                           n1191, A => n5843, ZN => n5842);
   U3207 : NOR4_X1 port map( A1 => n5764, A2 => n5765, A3 => n5766, A4 => n5767
                           , ZN => n5745);
   U3208 : OAI221_X1 port map( B1 => n61798, B2 => n1150, C1 => n61797, C2 => 
                           n1158, A => n5770, ZN => n5765);
   U3209 : OAI221_X1 port map( B1 => n5516, B2 => n1166, C1 => n5517, C2 => 
                           n1174, A => n5769, ZN => n5766);
   U3210 : OAI221_X1 port map( B1 => n61818, B2 => n1182, C1 => n61815, C2 => 
                           n1190, A => n5768, ZN => n5767);
   U3211 : NOR4_X1 port map( A1 => n5689, A2 => n5690, A3 => n5691, A4 => n5692
                           , ZN => n5670);
   U3212 : OAI221_X1 port map( B1 => n61798, B2 => n1149, C1 => n61797, C2 => 
                           n1157, A => n5695, ZN => n5690);
   U3213 : OAI221_X1 port map( B1 => n5516, B2 => n1165, C1 => n5517, C2 => 
                           n1173, A => n5694, ZN => n5691);
   U3214 : OAI221_X1 port map( B1 => n61818, B2 => n1181, C1 => n61815, C2 => 
                           n1189, A => n5693, ZN => n5692);
   U3215 : NOR4_X1 port map( A1 => n5614, A2 => n5615, A3 => n5616, A4 => n5617
                           , ZN => n5595);
   U3216 : OAI221_X1 port map( B1 => n61798, B2 => n1148, C1 => n61797, C2 => 
                           n1156, A => n5620, ZN => n5615);
   U3217 : OAI221_X1 port map( B1 => n5516, B2 => n1164, C1 => n5517, C2 => 
                           n1172, A => n5619, ZN => n5616);
   U3218 : OAI221_X1 port map( B1 => n61818, B2 => n1180, C1 => n61815, C2 => 
                           n1188, A => n5618, ZN => n5617);
   U3219 : NOR4_X1 port map( A1 => n5507, A2 => n5508, A3 => n5509, A4 => n5510
                           , ZN => n5464);
   U3220 : OAI221_X1 port map( B1 => n61798, B2 => n1147, C1 => n61797, C2 => 
                           n1155, A => n5523, ZN => n5508);
   U3221 : OAI221_X1 port map( B1 => n5516, B2 => n1163, C1 => n5517, C2 => 
                           n1171, A => n5518, ZN => n5509);
   U3222 : OAI221_X1 port map( B1 => n61818, B2 => n1179, C1 => n61815, C2 => 
                           n1187, A => n5513, ZN => n5510);
   U3223 : NOR4_X1 port map( A1 => n6770, A2 => n6771, A3 => n6772, A4 => n6773
                           , ZN => n6751);
   U3224 : OAI221_X1 port map( B1 => n61817, B2 => n3687, C1 => n61814, C2 => 
                           n3711, A => n6775, ZN => n6772);
   U3225 : OAI221_X1 port map( B1 => n6092, B2 => n3879, C1 => n61680, C2 => 
                           n3807, A => n6774, ZN => n6773);
   U3226 : OAI221_X1 port map( B1 => n61787, B2 => n3581, C1 => n61784, C2 => 
                           n3557, A => n6777, ZN => n6770);
   U3227 : NOR4_X1 port map( A1 => n6695, A2 => n6696, A3 => n6697, A4 => n6698
                           , ZN => n6676);
   U3228 : OAI221_X1 port map( B1 => n61817, B2 => n3686, C1 => n61814, C2 => 
                           n3710, A => n6700, ZN => n6697);
   U3229 : OAI221_X1 port map( B1 => n6092, B2 => n3878, C1 => n61680, C2 => 
                           n3806, A => n6699, ZN => n6698);
   U3230 : OAI221_X1 port map( B1 => n61787, B2 => n3580, C1 => n61784, C2 => 
                           n3556, A => n6702, ZN => n6695);
   U3231 : NOR4_X1 port map( A1 => n6620, A2 => n6621, A3 => n6622, A4 => n6623
                           , ZN => n6601);
   U3232 : OAI221_X1 port map( B1 => n61817, B2 => n3685, C1 => n61814, C2 => 
                           n3709, A => n6625, ZN => n6622);
   U3233 : OAI221_X1 port map( B1 => n6092, B2 => n3877, C1 => n61680, C2 => 
                           n3805, A => n6624, ZN => n6623);
   U3234 : OAI221_X1 port map( B1 => n61787, B2 => n3579, C1 => n61784, C2 => 
                           n3555, A => n6627, ZN => n6620);
   U3235 : NOR4_X1 port map( A1 => n6545, A2 => n6546, A3 => n6547, A4 => n6548
                           , ZN => n6526);
   U3236 : OAI221_X1 port map( B1 => n61817, B2 => n3684, C1 => n61814, C2 => 
                           n3708, A => n6550, ZN => n6547);
   U3237 : OAI221_X1 port map( B1 => n6092, B2 => n3876, C1 => n61680, C2 => 
                           n3804, A => n6549, ZN => n6548);
   U3238 : OAI221_X1 port map( B1 => n61787, B2 => n3578, C1 => n61784, C2 => 
                           n3554, A => n6552, ZN => n6545);
   U3239 : NOR4_X1 port map( A1 => n6470, A2 => n6471, A3 => n6472, A4 => n6473
                           , ZN => n6451);
   U3240 : OAI221_X1 port map( B1 => n61817, B2 => n3683, C1 => n61814, C2 => 
                           n3707, A => n6475, ZN => n6472);
   U3241 : OAI221_X1 port map( B1 => n6092, B2 => n3875, C1 => n61680, C2 => 
                           n3803, A => n6474, ZN => n6473);
   U3242 : OAI221_X1 port map( B1 => n61787, B2 => n3577, C1 => n61784, C2 => 
                           n3553, A => n6477, ZN => n6470);
   U3243 : NOR4_X1 port map( A1 => n6395, A2 => n6396, A3 => n6397, A4 => n6398
                           , ZN => n6376);
   U3244 : OAI221_X1 port map( B1 => n61817, B2 => n3682, C1 => n61814, C2 => 
                           n3706, A => n6400, ZN => n6397);
   U3245 : OAI221_X1 port map( B1 => n6092, B2 => n3874, C1 => n61680, C2 => 
                           n3802, A => n6399, ZN => n6398);
   U3246 : OAI221_X1 port map( B1 => n61787, B2 => n3576, C1 => n61784, C2 => 
                           n3552, A => n6402, ZN => n6395);
   U3247 : NOR4_X1 port map( A1 => n6320, A2 => n6321, A3 => n6322, A4 => n6323
                           , ZN => n6301);
   U3248 : OAI221_X1 port map( B1 => n61817, B2 => n3681, C1 => n61814, C2 => 
                           n3705, A => n6325, ZN => n6322);
   U3249 : OAI221_X1 port map( B1 => n6092, B2 => n3873, C1 => n61680, C2 => 
                           n3801, A => n6324, ZN => n6323);
   U3250 : OAI221_X1 port map( B1 => n61787, B2 => n3575, C1 => n61784, C2 => 
                           n3551, A => n6327, ZN => n6320);
   U3251 : NOR4_X1 port map( A1 => n6245, A2 => n6246, A3 => n6247, A4 => n6248
                           , ZN => n6226);
   U3252 : OAI221_X1 port map( B1 => n61817, B2 => n3680, C1 => n61814, C2 => 
                           n3704, A => n6250, ZN => n6247);
   U3253 : OAI221_X1 port map( B1 => n6092, B2 => n3872, C1 => n61680, C2 => 
                           n3800, A => n6249, ZN => n6248);
   U3254 : OAI221_X1 port map( B1 => n61787, B2 => n3574, C1 => n61784, C2 => 
                           n3550, A => n6252, ZN => n6245);
   U3255 : NOR4_X1 port map( A1 => n6170, A2 => n6171, A3 => n6172, A4 => n6173
                           , ZN => n6151);
   U3256 : OAI221_X1 port map( B1 => n61817, B2 => n3679, C1 => n61814, C2 => 
                           n3703, A => n6175, ZN => n6172);
   U3257 : OAI221_X1 port map( B1 => n6092, B2 => n3871, C1 => n61680, C2 => 
                           n3799, A => n6174, ZN => n6173);
   U3258 : OAI221_X1 port map( B1 => n61787, B2 => n3573, C1 => n61784, C2 => 
                           n3549, A => n6177, ZN => n6170);
   U3259 : NOR4_X1 port map( A1 => n7145, A2 => n7146, A3 => n7147, A4 => n7148
                           , ZN => n7126);
   U3260 : OAI221_X1 port map( B1 => n61816, B2 => n3692, C1 => n61813, C2 => 
                           n3716, A => n7150, ZN => n7147);
   U3261 : OAI221_X1 port map( B1 => n61677, B2 => n3884, C1 => n61679, C2 => 
                           n3812, A => n7149, ZN => n7148);
   U3262 : OAI221_X1 port map( B1 => n61786, B2 => n3586, C1 => n61783, C2 => 
                           n3562, A => n7152, ZN => n7145);
   U3263 : NOR4_X1 port map( A1 => n7070, A2 => n7071, A3 => n7072, A4 => n7073
                           , ZN => n7051);
   U3264 : OAI221_X1 port map( B1 => n61816, B2 => n3691, C1 => n61813, C2 => 
                           n3715, A => n7075, ZN => n7072);
   U3265 : OAI221_X1 port map( B1 => n61677, B2 => n3883, C1 => n61679, C2 => 
                           n3811, A => n7074, ZN => n7073);
   U3266 : OAI221_X1 port map( B1 => n61786, B2 => n3585, C1 => n61783, C2 => 
                           n3561, A => n7077, ZN => n7070);
   U3267 : NOR4_X1 port map( A1 => n6920, A2 => n6921, A3 => n6922, A4 => n6923
                           , ZN => n6901);
   U3268 : OAI221_X1 port map( B1 => n61817, B2 => n3689, C1 => n61814, C2 => 
                           n3713, A => n6925, ZN => n6922);
   U3269 : OAI221_X1 port map( B1 => n6092, B2 => n3881, C1 => n61680, C2 => 
                           n3809, A => n6924, ZN => n6923);
   U3270 : OAI221_X1 port map( B1 => n61787, B2 => n3583, C1 => n61784, C2 => 
                           n3559, A => n6927, ZN => n6920);
   U3271 : NOR4_X1 port map( A1 => n6845, A2 => n6846, A3 => n6847, A4 => n6848
                           , ZN => n6826);
   U3272 : OAI221_X1 port map( B1 => n61817, B2 => n3688, C1 => n61814, C2 => 
                           n3712, A => n6850, ZN => n6847);
   U3273 : OAI221_X1 port map( B1 => n6092, B2 => n3880, C1 => n61680, C2 => 
                           n3808, A => n6849, ZN => n6848);
   U3274 : OAI221_X1 port map( B1 => n61787, B2 => n3582, C1 => n61784, C2 => 
                           n3558, A => n6852, ZN => n6845);
   U3275 : NOR4_X1 port map( A1 => n7295, A2 => n7296, A3 => n7297, A4 => n7298
                           , ZN => n7276);
   U3276 : OAI221_X1 port map( B1 => n61816, B2 => n3694, C1 => n61813, C2 => 
                           n3718, A => n7300, ZN => n7297);
   U3277 : OAI221_X1 port map( B1 => n61677, B2 => n3886, C1 => n61679, C2 => 
                           n3814, A => n7299, ZN => n7298);
   U3278 : OAI221_X1 port map( B1 => n61786, B2 => n3588, C1 => n61783, C2 => 
                           n3564, A => n7302, ZN => n7295);
   U3279 : NOR4_X1 port map( A1 => n7925, A2 => n7926, A3 => n7927, A4 => n7928
                           , ZN => n7901);
   U3280 : OAI221_X1 port map( B1 => n61816, B2 => n3702, C1 => n61813, C2 => 
                           n3726, A => n7930, ZN => n7927);
   U3281 : OAI221_X1 port map( B1 => n61677, B2 => n3894, C1 => n61679, C2 => 
                           n3822, A => n7929, ZN => n7928);
   U3282 : OAI221_X1 port map( B1 => n61786, B2 => n3596, C1 => n61783, C2 => 
                           n3572, A => n7933, ZN => n7925);
   U3283 : NOR4_X1 port map( A1 => n7820, A2 => n7821, A3 => n7822, A4 => n7823
                           , ZN => n7801);
   U3284 : OAI221_X1 port map( B1 => n61816, B2 => n3701, C1 => n61813, C2 => 
                           n3725, A => n7825, ZN => n7822);
   U3285 : OAI221_X1 port map( B1 => n61677, B2 => n3893, C1 => n61679, C2 => 
                           n3821, A => n7824, ZN => n7823);
   U3286 : OAI221_X1 port map( B1 => n61786, B2 => n3595, C1 => n61783, C2 => 
                           n3571, A => n7827, ZN => n7820);
   U3287 : NOR4_X1 port map( A1 => n7745, A2 => n7746, A3 => n7747, A4 => n7748
                           , ZN => n7726);
   U3288 : OAI221_X1 port map( B1 => n61816, B2 => n3700, C1 => n61813, C2 => 
                           n3724, A => n7750, ZN => n7747);
   U3289 : OAI221_X1 port map( B1 => n61677, B2 => n3892, C1 => n61679, C2 => 
                           n3820, A => n7749, ZN => n7748);
   U3290 : OAI221_X1 port map( B1 => n61786, B2 => n3594, C1 => n61783, C2 => 
                           n3570, A => n7752, ZN => n7745);
   U3291 : NOR4_X1 port map( A1 => n7670, A2 => n7671, A3 => n7672, A4 => n7673
                           , ZN => n7651);
   U3292 : OAI221_X1 port map( B1 => n61816, B2 => n3699, C1 => n61813, C2 => 
                           n3723, A => n7675, ZN => n7672);
   U3293 : OAI221_X1 port map( B1 => n61677, B2 => n3891, C1 => n61679, C2 => 
                           n3819, A => n7674, ZN => n7673);
   U3294 : OAI221_X1 port map( B1 => n61786, B2 => n3593, C1 => n61783, C2 => 
                           n3569, A => n7677, ZN => n7670);
   U3295 : NOR4_X1 port map( A1 => n7595, A2 => n7596, A3 => n7597, A4 => n7598
                           , ZN => n7576);
   U3296 : OAI221_X1 port map( B1 => n61816, B2 => n3698, C1 => n61813, C2 => 
                           n3722, A => n7600, ZN => n7597);
   U3297 : OAI221_X1 port map( B1 => n61677, B2 => n3890, C1 => n61679, C2 => 
                           n3818, A => n7599, ZN => n7598);
   U3298 : OAI221_X1 port map( B1 => n61786, B2 => n3592, C1 => n61783, C2 => 
                           n3568, A => n7602, ZN => n7595);
   U3299 : NOR4_X1 port map( A1 => n7520, A2 => n7521, A3 => n7522, A4 => n7523
                           , ZN => n7501);
   U3300 : OAI221_X1 port map( B1 => n61816, B2 => n3697, C1 => n61813, C2 => 
                           n3721, A => n7525, ZN => n7522);
   U3301 : OAI221_X1 port map( B1 => n61677, B2 => n3889, C1 => n61679, C2 => 
                           n3817, A => n7524, ZN => n7523);
   U3302 : OAI221_X1 port map( B1 => n61786, B2 => n3591, C1 => n61783, C2 => 
                           n3567, A => n7527, ZN => n7520);
   U3303 : NOR4_X1 port map( A1 => n7445, A2 => n7446, A3 => n7447, A4 => n7448
                           , ZN => n7426);
   U3304 : OAI221_X1 port map( B1 => n61816, B2 => n3696, C1 => n61813, C2 => 
                           n3720, A => n7450, ZN => n7447);
   U3305 : OAI221_X1 port map( B1 => n61677, B2 => n3888, C1 => n61679, C2 => 
                           n3816, A => n7449, ZN => n7448);
   U3306 : OAI221_X1 port map( B1 => n61786, B2 => n3590, C1 => n61783, C2 => 
                           n3566, A => n7452, ZN => n7445);
   U3307 : NOR4_X1 port map( A1 => n7370, A2 => n7371, A3 => n7372, A4 => n7373
                           , ZN => n7351);
   U3308 : OAI221_X1 port map( B1 => n61816, B2 => n3695, C1 => n61813, C2 => 
                           n3719, A => n7375, ZN => n7372);
   U3309 : OAI221_X1 port map( B1 => n61677, B2 => n3887, C1 => n61679, C2 => 
                           n3815, A => n7374, ZN => n7373);
   U3310 : OAI221_X1 port map( B1 => n61786, B2 => n3589, C1 => n61783, C2 => 
                           n3565, A => n7377, ZN => n7370);
   U3311 : NOR4_X1 port map( A1 => n7220, A2 => n7221, A3 => n7222, A4 => n7223
                           , ZN => n7201);
   U3312 : OAI221_X1 port map( B1 => n61816, B2 => n3693, C1 => n61813, C2 => 
                           n3717, A => n7225, ZN => n7222);
   U3313 : OAI221_X1 port map( B1 => n61677, B2 => n3885, C1 => n61679, C2 => 
                           n3813, A => n7224, ZN => n7223);
   U3314 : OAI221_X1 port map( B1 => n61786, B2 => n3587, C1 => n61783, C2 => 
                           n3563, A => n7227, ZN => n7220);
   U3315 : NOR4_X1 port map( A1 => n6995, A2 => n6996, A3 => n6997, A4 => n6998
                           , ZN => n6976);
   U3316 : OAI221_X1 port map( B1 => n61817, B2 => n3690, C1 => n61814, C2 => 
                           n3714, A => n7000, ZN => n6997);
   U3317 : OAI221_X1 port map( B1 => n6092, B2 => n3882, C1 => n61680, C2 => 
                           n3810, A => n6999, ZN => n6998);
   U3318 : OAI221_X1 port map( B1 => n61787, B2 => n3584, C1 => n61784, C2 => 
                           n3560, A => n7002, ZN => n6995);
   U3319 : NOR4_X1 port map( A1 => n8628, A2 => n8629, A3 => n8630, A4 => n8631
                           , ZN => n8609);
   U3320 : OAI221_X1 port map( B1 => n4240, B2 => n61540, C1 => n993, C2 => 
                           n61537, A => n8634, ZN => n8629);
   U3321 : OAI221_X1 port map( B1 => n1005, B2 => n61552, C1 => n1013, C2 => 
                           n61549, A => n8633, ZN => n8630);
   U3322 : OAI221_X1 port map( B1 => n1021, B2 => n61564, C1 => n1029, C2 => 
                           n61561, A => n8632, ZN => n8631);
   U3323 : NOR4_X1 port map( A1 => n8664, A2 => n8665, A3 => n8666, A4 => n8667
                           , ZN => n8645);
   U3324 : OAI221_X1 port map( B1 => n1122, B2 => n61336, C1 => n1130, C2 => 
                           n61333, A => n8670, ZN => n8665);
   U3325 : OAI221_X1 port map( B1 => n1154, B2 => n61348, C1 => n1162, C2 => 
                           n61345, A => n8669, ZN => n8666);
   U3326 : OAI221_X1 port map( B1 => n1186, B2 => n61360, C1 => n1194, C2 => 
                           n61357, A => n8668, ZN => n8667);
   U3327 : NOR4_X1 port map( A1 => n8553, A2 => n8554, A3 => n8555, A4 => n8556
                           , ZN => n8534);
   U3328 : OAI221_X1 port map( B1 => n4239, B2 => n61540, C1 => n992, C2 => 
                           n61537, A => n8559, ZN => n8554);
   U3329 : OAI221_X1 port map( B1 => n1004, B2 => n61552, C1 => n1012, C2 => 
                           n61549, A => n8558, ZN => n8555);
   U3330 : OAI221_X1 port map( B1 => n1020, B2 => n61564, C1 => n1028, C2 => 
                           n61561, A => n8557, ZN => n8556);
   U3331 : NOR4_X1 port map( A1 => n8589, A2 => n8590, A3 => n8591, A4 => n8592
                           , ZN => n8570);
   U3332 : OAI221_X1 port map( B1 => n1121, B2 => n61336, C1 => n1129, C2 => 
                           n61333, A => n8595, ZN => n8590);
   U3333 : OAI221_X1 port map( B1 => n1153, B2 => n61348, C1 => n1161, C2 => 
                           n61345, A => n8594, ZN => n8591);
   U3334 : OAI221_X1 port map( B1 => n1185, B2 => n61360, C1 => n1193, C2 => 
                           n61357, A => n8593, ZN => n8592);
   U3335 : NOR4_X1 port map( A1 => n8478, A2 => n8479, A3 => n8480, A4 => n8481
                           , ZN => n8459);
   U3336 : OAI221_X1 port map( B1 => n4238, B2 => n61540, C1 => n991, C2 => 
                           n61537, A => n8484, ZN => n8479);
   U3337 : OAI221_X1 port map( B1 => n1003, B2 => n61552, C1 => n1011, C2 => 
                           n61549, A => n8483, ZN => n8480);
   U3338 : OAI221_X1 port map( B1 => n1019, B2 => n61564, C1 => n1027, C2 => 
                           n61561, A => n8482, ZN => n8481);
   U3339 : NOR4_X1 port map( A1 => n8514, A2 => n8515, A3 => n8516, A4 => n8517
                           , ZN => n8495);
   U3340 : OAI221_X1 port map( B1 => n1120, B2 => n61336, C1 => n1128, C2 => 
                           n61333, A => n8520, ZN => n8515);
   U3341 : OAI221_X1 port map( B1 => n1152, B2 => n61348, C1 => n1160, C2 => 
                           n61345, A => n8519, ZN => n8516);
   U3342 : OAI221_X1 port map( B1 => n1184, B2 => n61360, C1 => n1192, C2 => 
                           n61357, A => n8518, ZN => n8517);
   U3343 : NOR4_X1 port map( A1 => n8403, A2 => n8404, A3 => n8405, A4 => n8406
                           , ZN => n8384);
   U3344 : OAI221_X1 port map( B1 => n4237, B2 => n61540, C1 => n990, C2 => 
                           n61537, A => n8409, ZN => n8404);
   U3345 : OAI221_X1 port map( B1 => n1002, B2 => n61552, C1 => n1010, C2 => 
                           n61549, A => n8408, ZN => n8405);
   U3346 : OAI221_X1 port map( B1 => n1018, B2 => n61564, C1 => n1026, C2 => 
                           n61561, A => n8407, ZN => n8406);
   U3347 : NOR4_X1 port map( A1 => n8439, A2 => n8440, A3 => n8441, A4 => n8442
                           , ZN => n8420);
   U3348 : OAI221_X1 port map( B1 => n1119, B2 => n61336, C1 => n1127, C2 => 
                           n61333, A => n8445, ZN => n8440);
   U3349 : OAI221_X1 port map( B1 => n1151, B2 => n61348, C1 => n1159, C2 => 
                           n61345, A => n8444, ZN => n8441);
   U3350 : OAI221_X1 port map( B1 => n1183, B2 => n61360, C1 => n1191, C2 => 
                           n61357, A => n8443, ZN => n8442);
   U3351 : NOR4_X1 port map( A1 => n8328, A2 => n8329, A3 => n8330, A4 => n8331
                           , ZN => n8309);
   U3352 : OAI221_X1 port map( B1 => n4236, B2 => n61540, C1 => n989, C2 => 
                           n61537, A => n8334, ZN => n8329);
   U3353 : OAI221_X1 port map( B1 => n1001, B2 => n61552, C1 => n1009, C2 => 
                           n61549, A => n8333, ZN => n8330);
   U3354 : OAI221_X1 port map( B1 => n1017, B2 => n61564, C1 => n1025, C2 => 
                           n61561, A => n8332, ZN => n8331);
   U3355 : NOR4_X1 port map( A1 => n8364, A2 => n8365, A3 => n8366, A4 => n8367
                           , ZN => n8345);
   U3356 : OAI221_X1 port map( B1 => n1118, B2 => n61336, C1 => n1126, C2 => 
                           n61333, A => n8370, ZN => n8365);
   U3357 : OAI221_X1 port map( B1 => n1150, B2 => n61348, C1 => n1158, C2 => 
                           n61345, A => n8369, ZN => n8366);
   U3358 : OAI221_X1 port map( B1 => n1182, B2 => n61360, C1 => n1190, C2 => 
                           n61357, A => n8368, ZN => n8367);
   U3359 : NOR4_X1 port map( A1 => n8253, A2 => n8254, A3 => n8255, A4 => n8256
                           , ZN => n8234);
   U3360 : OAI221_X1 port map( B1 => n985, B2 => n61540, C1 => n988, C2 => 
                           n61537, A => n8259, ZN => n8254);
   U3361 : OAI221_X1 port map( B1 => n1000, B2 => n61552, C1 => n1008, C2 => 
                           n61549, A => n8258, ZN => n8255);
   U3362 : OAI221_X1 port map( B1 => n1016, B2 => n61564, C1 => n1024, C2 => 
                           n61561, A => n8257, ZN => n8256);
   U3363 : NOR4_X1 port map( A1 => n8289, A2 => n8290, A3 => n8291, A4 => n8292
                           , ZN => n8270);
   U3364 : OAI221_X1 port map( B1 => n1117, B2 => n61336, C1 => n1125, C2 => 
                           n61333, A => n8295, ZN => n8290);
   U3365 : OAI221_X1 port map( B1 => n1149, B2 => n61348, C1 => n1157, C2 => 
                           n61345, A => n8294, ZN => n8291);
   U3366 : OAI221_X1 port map( B1 => n1181, B2 => n61360, C1 => n1189, C2 => 
                           n61357, A => n8293, ZN => n8292);
   U3367 : NOR4_X1 port map( A1 => n8178, A2 => n8179, A3 => n8180, A4 => n8181
                           , ZN => n8159);
   U3368 : OAI221_X1 port map( B1 => n984, B2 => n61540, C1 => n987, C2 => 
                           n61537, A => n8184, ZN => n8179);
   U3369 : OAI221_X1 port map( B1 => n995, B2 => n61552, C1 => n1007, C2 => 
                           n61549, A => n8183, ZN => n8180);
   U3370 : OAI221_X1 port map( B1 => n1015, B2 => n61564, C1 => n1023, C2 => 
                           n61561, A => n8182, ZN => n8181);
   U3371 : NOR4_X1 port map( A1 => n8214, A2 => n8215, A3 => n8216, A4 => n8217
                           , ZN => n8195);
   U3372 : OAI221_X1 port map( B1 => n1116, B2 => n61336, C1 => n1124, C2 => 
                           n61333, A => n8220, ZN => n8215);
   U3373 : OAI221_X1 port map( B1 => n1148, B2 => n61348, C1 => n1156, C2 => 
                           n61345, A => n8219, ZN => n8216);
   U3374 : OAI221_X1 port map( B1 => n1180, B2 => n61360, C1 => n1188, C2 => 
                           n61357, A => n8218, ZN => n8217);
   U3375 : NOR4_X1 port map( A1 => n8001, A2 => n8002, A3 => n8003, A4 => n8004
                           , ZN => n7948);
   U3376 : OAI221_X1 port map( B1 => n983, B2 => n61540, C1 => n986, C2 => 
                           n61537, A => n8017, ZN => n8002);
   U3377 : OAI221_X1 port map( B1 => n994, B2 => n61552, C1 => n1006, C2 => 
                           n61549, A => n8012, ZN => n8003);
   U3378 : OAI221_X1 port map( B1 => n1014, B2 => n61564, C1 => n1022, C2 => 
                           n61561, A => n8007, ZN => n8004);
   U3379 : NOR4_X1 port map( A1 => n8105, A2 => n8106, A3 => n8107, A4 => n8108
                           , ZN => n8052);
   U3380 : OAI221_X1 port map( B1 => n1115, B2 => n61336, C1 => n1123, C2 => 
                           n61333, A => n8121, ZN => n8106);
   U3381 : OAI221_X1 port map( B1 => n1147, B2 => n61348, C1 => n1155, C2 => 
                           n61345, A => n8116, ZN => n8107);
   U3382 : OAI221_X1 port map( B1 => n1179, B2 => n61360, C1 => n1187, C2 => 
                           n61357, A => n8111, ZN => n8108);
   U3383 : NOR2_X1 port map( A1 => ADDR_WR(1), A2 => ADDR_WR(0), ZN => n15257);
   U3384 : NOR4_X1 port map( A1 => n7267, A2 => n7268, A3 => n7269, A4 => n7270
                           , ZN => n7239);
   U3385 : OAI221_X1 port map( B1 => n61709, B2 => n3200, C1 => n61711, C2 => 
                           n3142, A => n7272, ZN => n7269);
   U3386 : OAI221_X1 port map( B1 => n61705, B2 => n2926, C1 => n61707, C2 => 
                           n2950, A => n7273, ZN => n7268);
   U3387 : OAI221_X1 port map( B1 => n61948, B2 => n2770, C1 => n61947, C2 => 
                           n2764, A => n7271, ZN => n7270);
   U3388 : NOR4_X1 port map( A1 => n7642, A2 => n7643, A3 => n7644, A4 => n7645
                           , ZN => n7614);
   U3389 : OAI221_X1 port map( B1 => n61709, B2 => n3205, C1 => n61711, C2 => 
                           n3147, A => n7647, ZN => n7644);
   U3390 : OAI221_X1 port map( B1 => n61705, B2 => n2931, C1 => n61707, C2 => 
                           n2955, A => n7648, ZN => n7643);
   U3391 : OAI221_X1 port map( B1 => n61948, B2 => n2775, C1 => n61947, C2 => 
                           n2769, A => n7646, ZN => n7645);
   U3392 : NOR4_X1 port map( A1 => n7567, A2 => n7568, A3 => n7569, A4 => n7570
                           , ZN => n7539);
   U3393 : OAI221_X1 port map( B1 => n61709, B2 => n3204, C1 => n61711, C2 => 
                           n3146, A => n7572, ZN => n7569);
   U3394 : OAI221_X1 port map( B1 => n61705, B2 => n2930, C1 => n61707, C2 => 
                           n2954, A => n7573, ZN => n7568);
   U3395 : OAI221_X1 port map( B1 => n61948, B2 => n2774, C1 => n61947, C2 => 
                           n2768, A => n7571, ZN => n7570);
   U3396 : NOR4_X1 port map( A1 => n7492, A2 => n7493, A3 => n7494, A4 => n7495
                           , ZN => n7464);
   U3397 : OAI221_X1 port map( B1 => n61709, B2 => n3203, C1 => n61711, C2 => 
                           n3145, A => n7497, ZN => n7494);
   U3398 : OAI221_X1 port map( B1 => n61705, B2 => n2929, C1 => n61707, C2 => 
                           n2953, A => n7498, ZN => n7493);
   U3399 : OAI221_X1 port map( B1 => n61948, B2 => n2773, C1 => n61947, C2 => 
                           n2767, A => n7496, ZN => n7495);
   U3400 : NOR4_X1 port map( A1 => n7417, A2 => n7418, A3 => n7419, A4 => n7420
                           , ZN => n7389);
   U3401 : OAI221_X1 port map( B1 => n61709, B2 => n3202, C1 => n61711, C2 => 
                           n3144, A => n7422, ZN => n7419);
   U3402 : OAI221_X1 port map( B1 => n61705, B2 => n2928, C1 => n61707, C2 => 
                           n2952, A => n7423, ZN => n7418);
   U3403 : OAI221_X1 port map( B1 => n61948, B2 => n2772, C1 => n61947, C2 => 
                           n2766, A => n7421, ZN => n7420);
   U3404 : NOR4_X1 port map( A1 => n7342, A2 => n7343, A3 => n7344, A4 => n7345
                           , ZN => n7314);
   U3405 : OAI221_X1 port map( B1 => n61709, B2 => n3201, C1 => n61711, C2 => 
                           n3143, A => n7347, ZN => n7344);
   U3406 : OAI221_X1 port map( B1 => n61705, B2 => n2927, C1 => n61707, C2 => 
                           n2951, A => n7348, ZN => n7343);
   U3407 : OAI221_X1 port map( B1 => n61948, B2 => n2771, C1 => n61947, C2 => 
                           n2765, A => n7346, ZN => n7345);
   U3408 : NOR4_X1 port map( A1 => n6778, A2 => n6779, A3 => n6780, A4 => n6781
                           , ZN => n6750);
   U3409 : OAI221_X1 port map( B1 => n61748, B2 => n1358, C1 => n61745, C2 => 
                           n1323, A => n6785, ZN => n6778);
   U3410 : OAI221_X1 port map( B1 => n61760, B2 => n1395, C1 => n61757, C2 => 
                           n1371, A => n6784, ZN => n6779);
   U3411 : OAI221_X1 port map( B1 => n61772, B2 => n3365, C1 => n61769, C2 => 
                           n3341, A => n6783, ZN => n6780);
   U3412 : NOR4_X1 port map( A1 => n6703, A2 => n6704, A3 => n6705, A4 => n6706
                           , ZN => n6675);
   U3413 : OAI221_X1 port map( B1 => n61748, B2 => n1357, C1 => n61745, C2 => 
                           n1322, A => n6710, ZN => n6703);
   U3414 : OAI221_X1 port map( B1 => n61760, B2 => n1394, C1 => n61757, C2 => 
                           n1370, A => n6709, ZN => n6704);
   U3415 : OAI221_X1 port map( B1 => n61772, B2 => n3364, C1 => n61769, C2 => 
                           n3340, A => n6708, ZN => n6705);
   U3416 : NOR4_X1 port map( A1 => n6628, A2 => n6629, A3 => n6630, A4 => n6631
                           , ZN => n6600);
   U3417 : OAI221_X1 port map( B1 => n61748, B2 => n1356, C1 => n61745, C2 => 
                           n1321, A => n6635, ZN => n6628);
   U3418 : OAI221_X1 port map( B1 => n61760, B2 => n1393, C1 => n61757, C2 => 
                           n1369, A => n6634, ZN => n6629);
   U3419 : OAI221_X1 port map( B1 => n61772, B2 => n3363, C1 => n61769, C2 => 
                           n3339, A => n6633, ZN => n6630);
   U3420 : NOR4_X1 port map( A1 => n6553, A2 => n6554, A3 => n6555, A4 => n6556
                           , ZN => n6525);
   U3421 : OAI221_X1 port map( B1 => n61748, B2 => n1355, C1 => n61745, C2 => 
                           n1320, A => n6560, ZN => n6553);
   U3422 : OAI221_X1 port map( B1 => n61760, B2 => n1392, C1 => n61757, C2 => 
                           n1368, A => n6559, ZN => n6554);
   U3423 : OAI221_X1 port map( B1 => n61772, B2 => n3362, C1 => n61769, C2 => 
                           n3338, A => n6558, ZN => n6555);
   U3424 : NOR4_X1 port map( A1 => n6478, A2 => n6479, A3 => n6480, A4 => n6481
                           , ZN => n6450);
   U3425 : OAI221_X1 port map( B1 => n61748, B2 => n1354, C1 => n61745, C2 => 
                           n1319, A => n6485, ZN => n6478);
   U3426 : OAI221_X1 port map( B1 => n61760, B2 => n1391, C1 => n61757, C2 => 
                           n1367, A => n6484, ZN => n6479);
   U3427 : OAI221_X1 port map( B1 => n61772, B2 => n3361, C1 => n61769, C2 => 
                           n3337, A => n6483, ZN => n6480);
   U3428 : NOR4_X1 port map( A1 => n6403, A2 => n6404, A3 => n6405, A4 => n6406
                           , ZN => n6375);
   U3429 : OAI221_X1 port map( B1 => n61748, B2 => n1353, C1 => n61745, C2 => 
                           n1318, A => n6410, ZN => n6403);
   U3430 : OAI221_X1 port map( B1 => n61760, B2 => n1390, C1 => n61757, C2 => 
                           n1366, A => n6409, ZN => n6404);
   U3431 : OAI221_X1 port map( B1 => n61772, B2 => n3360, C1 => n61768, C2 => 
                           n3336, A => n6408, ZN => n6405);
   U3432 : NOR4_X1 port map( A1 => n6328, A2 => n6329, A3 => n6330, A4 => n6331
                           , ZN => n6300);
   U3433 : OAI221_X1 port map( B1 => n61748, B2 => n1352, C1 => n61745, C2 => 
                           n1317, A => n6335, ZN => n6328);
   U3434 : OAI221_X1 port map( B1 => n61760, B2 => n1389, C1 => n61757, C2 => 
                           n1365, A => n6334, ZN => n6329);
   U3435 : OAI221_X1 port map( B1 => n61772, B2 => n3359, C1 => n61768, C2 => 
                           n3335, A => n6333, ZN => n6330);
   U3436 : NOR4_X1 port map( A1 => n6253, A2 => n6254, A3 => n6255, A4 => n6256
                           , ZN => n6225);
   U3437 : OAI221_X1 port map( B1 => n61748, B2 => n1351, C1 => n61745, C2 => 
                           n1316, A => n6260, ZN => n6253);
   U3438 : OAI221_X1 port map( B1 => n61760, B2 => n1388, C1 => n61757, C2 => 
                           n1364, A => n6259, ZN => n6254);
   U3439 : OAI221_X1 port map( B1 => n61772, B2 => n3358, C1 => n61768, C2 => 
                           n3334, A => n6258, ZN => n6255);
   U3440 : NOR4_X1 port map( A1 => n6178, A2 => n6179, A3 => n6180, A4 => n6181
                           , ZN => n6150);
   U3441 : OAI221_X1 port map( B1 => n61748, B2 => n1350, C1 => n61745, C2 => 
                           n1315, A => n6185, ZN => n6178);
   U3442 : OAI221_X1 port map( B1 => n61760, B2 => n1387, C1 => n61757, C2 => 
                           n1363, A => n6184, ZN => n6179);
   U3443 : OAI221_X1 port map( B1 => n61772, B2 => n3357, C1 => n61768, C2 => 
                           n3333, A => n6183, ZN => n6180);
   U3444 : NOR4_X1 port map( A1 => n7153, A2 => n7154, A3 => n7155, A4 => n7156
                           , ZN => n7125);
   U3445 : OAI221_X1 port map( B1 => n61747, B2 => n1328, C1 => n61744, C2 => 
                           n1339, A => n7160, ZN => n7153);
   U3446 : OAI221_X1 port map( B1 => n61759, B2 => n1400, C1 => n61756, C2 => 
                           n1376, A => n7159, ZN => n7154);
   U3447 : OAI221_X1 port map( B1 => n61771, B2 => n3370, C1 => n61769, C2 => 
                           n3346, A => n7158, ZN => n7155);
   U3448 : NOR4_X1 port map( A1 => n7078, A2 => n7079, A3 => n7080, A4 => n7081
                           , ZN => n7050);
   U3449 : OAI221_X1 port map( B1 => n61747, B2 => n1362, C1 => n61744, C2 => 
                           n1327, A => n7085, ZN => n7078);
   U3450 : OAI221_X1 port map( B1 => n61759, B2 => n1399, C1 => n61756, C2 => 
                           n1375, A => n7084, ZN => n7079);
   U3451 : OAI221_X1 port map( B1 => n61771, B2 => n3369, C1 => n61769, C2 => 
                           n3345, A => n7083, ZN => n7080);
   U3452 : NOR4_X1 port map( A1 => n6928, A2 => n6929, A3 => n6930, A4 => n6931
                           , ZN => n6900);
   U3453 : OAI221_X1 port map( B1 => n61748, B2 => n1360, C1 => n61745, C2 => 
                           n1325, A => n6935, ZN => n6928);
   U3454 : OAI221_X1 port map( B1 => n61760, B2 => n1397, C1 => n61757, C2 => 
                           n1373, A => n6934, ZN => n6929);
   U3455 : OAI221_X1 port map( B1 => n61772, B2 => n3367, C1 => n61769, C2 => 
                           n3343, A => n6933, ZN => n6930);
   U3456 : NOR4_X1 port map( A1 => n6853, A2 => n6854, A3 => n6855, A4 => n6856
                           , ZN => n6825);
   U3457 : OAI221_X1 port map( B1 => n61748, B2 => n1359, C1 => n61745, C2 => 
                           n1324, A => n6860, ZN => n6853);
   U3458 : OAI221_X1 port map( B1 => n61760, B2 => n1396, C1 => n61757, C2 => 
                           n1372, A => n6859, ZN => n6854);
   U3459 : OAI221_X1 port map( B1 => n61772, B2 => n3366, C1 => n61769, C2 => 
                           n3342, A => n6858, ZN => n6855);
   U3460 : NOR4_X1 port map( A1 => n7303, A2 => n7304, A3 => n7305, A4 => n7306
                           , ZN => n7275);
   U3461 : OAI221_X1 port map( B1 => n61747, B2 => n1330, C1 => n61744, C2 => 
                           n1341, A => n7310, ZN => n7303);
   U3462 : OAI221_X1 port map( B1 => n61759, B2 => n1402, C1 => n61756, C2 => 
                           n1378, A => n7309, ZN => n7304);
   U3463 : OAI221_X1 port map( B1 => n61771, B2 => n3372, C1 => n61769, C2 => 
                           n3348, A => n7308, ZN => n7305);
   U3464 : NOR4_X1 port map( A1 => n7935, A2 => n7936, A3 => n7937, A4 => n7938
                           , ZN => n7900);
   U3465 : OAI221_X1 port map( B1 => n61747, B2 => n1338, C1 => n61744, C2 => 
                           n1349, A => n7942, ZN => n7935);
   U3466 : OAI221_X1 port map( B1 => n61759, B2 => n1410, C1 => n61756, C2 => 
                           n1386, A => n7941, ZN => n7936);
   U3467 : OAI221_X1 port map( B1 => n61771, B2 => n3380, C1 => n61770, C2 => 
                           n3356, A => n7940, ZN => n7937);
   U3468 : NOR4_X1 port map( A1 => n7828, A2 => n7829, A3 => n7830, A4 => n7831
                           , ZN => n7800);
   U3469 : OAI221_X1 port map( B1 => n61747, B2 => n1337, C1 => n61744, C2 => 
                           n1348, A => n7835, ZN => n7828);
   U3470 : OAI221_X1 port map( B1 => n61759, B2 => n1409, C1 => n61756, C2 => 
                           n1385, A => n7834, ZN => n7829);
   U3471 : OAI221_X1 port map( B1 => n61771, B2 => n3379, C1 => n61770, C2 => 
                           n3355, A => n7833, ZN => n7830);
   U3472 : NOR4_X1 port map( A1 => n7753, A2 => n7754, A3 => n7755, A4 => n7756
                           , ZN => n7725);
   U3473 : OAI221_X1 port map( B1 => n61747, B2 => n1336, C1 => n61744, C2 => 
                           n1347, A => n7760, ZN => n7753);
   U3474 : OAI221_X1 port map( B1 => n61759, B2 => n1408, C1 => n61756, C2 => 
                           n1384, A => n7759, ZN => n7754);
   U3475 : OAI221_X1 port map( B1 => n61771, B2 => n3378, C1 => n61770, C2 => 
                           n3354, A => n7758, ZN => n7755);
   U3476 : NOR4_X1 port map( A1 => n7678, A2 => n7679, A3 => n7680, A4 => n7681
                           , ZN => n7650);
   U3477 : OAI221_X1 port map( B1 => n61747, B2 => n1335, C1 => n61744, C2 => 
                           n1346, A => n7685, ZN => n7678);
   U3478 : OAI221_X1 port map( B1 => n61759, B2 => n1407, C1 => n61756, C2 => 
                           n1383, A => n7684, ZN => n7679);
   U3479 : OAI221_X1 port map( B1 => n61771, B2 => n3377, C1 => n61770, C2 => 
                           n3353, A => n7683, ZN => n7680);
   U3480 : NOR4_X1 port map( A1 => n7603, A2 => n7604, A3 => n7605, A4 => n7606
                           , ZN => n7575);
   U3481 : OAI221_X1 port map( B1 => n61747, B2 => n1334, C1 => n61744, C2 => 
                           n1345, A => n7610, ZN => n7603);
   U3482 : OAI221_X1 port map( B1 => n61759, B2 => n1406, C1 => n61756, C2 => 
                           n1382, A => n7609, ZN => n7604);
   U3483 : OAI221_X1 port map( B1 => n61771, B2 => n3376, C1 => n61770, C2 => 
                           n3352, A => n7608, ZN => n7605);
   U3484 : NOR4_X1 port map( A1 => n7528, A2 => n7529, A3 => n7530, A4 => n7531
                           , ZN => n7500);
   U3485 : OAI221_X1 port map( B1 => n61747, B2 => n1333, C1 => n61744, C2 => 
                           n1344, A => n7535, ZN => n7528);
   U3486 : OAI221_X1 port map( B1 => n61759, B2 => n1405, C1 => n61756, C2 => 
                           n1381, A => n7534, ZN => n7529);
   U3487 : OAI221_X1 port map( B1 => n61771, B2 => n3375, C1 => n61770, C2 => 
                           n3351, A => n7533, ZN => n7530);
   U3488 : NOR4_X1 port map( A1 => n7453, A2 => n7454, A3 => n7455, A4 => n7456
                           , ZN => n7425);
   U3489 : OAI221_X1 port map( B1 => n61747, B2 => n1332, C1 => n61744, C2 => 
                           n1343, A => n7460, ZN => n7453);
   U3490 : OAI221_X1 port map( B1 => n61759, B2 => n1404, C1 => n61756, C2 => 
                           n1380, A => n7459, ZN => n7454);
   U3491 : OAI221_X1 port map( B1 => n61771, B2 => n3374, C1 => n61770, C2 => 
                           n3350, A => n7458, ZN => n7455);
   U3492 : NOR4_X1 port map( A1 => n7378, A2 => n7379, A3 => n7380, A4 => n7381
                           , ZN => n7350);
   U3493 : OAI221_X1 port map( B1 => n61747, B2 => n1331, C1 => n61744, C2 => 
                           n1342, A => n7385, ZN => n7378);
   U3494 : OAI221_X1 port map( B1 => n61759, B2 => n1403, C1 => n61756, C2 => 
                           n1379, A => n7384, ZN => n7379);
   U3495 : OAI221_X1 port map( B1 => n61771, B2 => n3373, C1 => n61769, C2 => 
                           n3349, A => n7383, ZN => n7380);
   U3496 : NOR4_X1 port map( A1 => n7228, A2 => n7229, A3 => n7230, A4 => n7231
                           , ZN => n7200);
   U3497 : OAI221_X1 port map( B1 => n61747, B2 => n1329, C1 => n61744, C2 => 
                           n1340, A => n7235, ZN => n7228);
   U3498 : OAI221_X1 port map( B1 => n61759, B2 => n1401, C1 => n61756, C2 => 
                           n1377, A => n7234, ZN => n7229);
   U3499 : OAI221_X1 port map( B1 => n61771, B2 => n3371, C1 => n61769, C2 => 
                           n3347, A => n7233, ZN => n7230);
   U3500 : NOR4_X1 port map( A1 => n7003, A2 => n7004, A3 => n7005, A4 => n7006
                           , ZN => n6975);
   U3501 : OAI221_X1 port map( B1 => n61748, B2 => n1361, C1 => n61745, C2 => 
                           n1326, A => n7010, ZN => n7003);
   U3502 : OAI221_X1 port map( B1 => n61760, B2 => n1398, C1 => n61757, C2 => 
                           n1374, A => n7009, ZN => n7004);
   U3503 : OAI221_X1 port map( B1 => n61772, B2 => n3368, C1 => n61769, C2 => 
                           n3344, A => n7008, ZN => n7005);
   U3504 : NOR4_X1 port map( A1 => n6101, A2 => n6102, A3 => n6103, A4 => n6104
                           , ZN => n6063);
   U3505 : OAI221_X1 port map( B1 => n61749, B2 => n19, C1 => n61746, C2 => n11
                           , A => n6110, ZN => n6101);
   U3506 : OAI221_X1 port map( B1 => n5536, B2 => n1113, C1 => n5537, C2 => 
                           n1097, A => n6105, ZN => n6104);
   U3507 : OAI221_X1 port map( B1 => n61761, B2 => n35, C1 => n61758, C2 => n27
                           , A => n6109, ZN => n6102);
   U3508 : NOR4_X1 port map( A1 => n5997, A2 => n5998, A3 => n5999, A4 => n6000
                           , ZN => n5969);
   U3509 : OAI221_X1 port map( B1 => n61749, B2 => n18, C1 => n61746, C2 => n10
                           , A => n6004, ZN => n5997);
   U3510 : OAI221_X1 port map( B1 => n5536, B2 => n1112, C1 => n5537, C2 => 
                           n1096, A => n6001, ZN => n6000);
   U3511 : OAI221_X1 port map( B1 => n61761, B2 => n34, C1 => n61758, C2 => n26
                           , A => n6003, ZN => n5998);
   U3512 : NOR4_X1 port map( A1 => n5922, A2 => n5923, A3 => n5924, A4 => n5925
                           , ZN => n5894);
   U3513 : OAI221_X1 port map( B1 => n61749, B2 => n17, C1 => n61746, C2 => n9,
                           A => n5929, ZN => n5922);
   U3514 : OAI221_X1 port map( B1 => n5536, B2 => n1111, C1 => n5537, C2 => 
                           n1095, A => n5926, ZN => n5925);
   U3515 : OAI221_X1 port map( B1 => n61761, B2 => n33, C1 => n61758, C2 => n25
                           , A => n5928, ZN => n5923);
   U3516 : NOR4_X1 port map( A1 => n5847, A2 => n5848, A3 => n5849, A4 => n5850
                           , ZN => n5819);
   U3517 : OAI221_X1 port map( B1 => n61749, B2 => n16, C1 => n61746, C2 => n8,
                           A => n5854, ZN => n5847);
   U3518 : OAI221_X1 port map( B1 => n5536, B2 => n1110, C1 => n5537, C2 => 
                           n1094, A => n5851, ZN => n5850);
   U3519 : OAI221_X1 port map( B1 => n61761, B2 => n32, C1 => n61758, C2 => n24
                           , A => n5853, ZN => n5848);
   U3520 : NOR4_X1 port map( A1 => n5772, A2 => n5773, A3 => n5774, A4 => n5775
                           , ZN => n5744);
   U3521 : OAI221_X1 port map( B1 => n61749, B2 => n15, C1 => n61746, C2 => n7,
                           A => n5779, ZN => n5772);
   U3522 : OAI221_X1 port map( B1 => n5536, B2 => n1109, C1 => n5537, C2 => 
                           n1093, A => n5776, ZN => n5775);
   U3523 : OAI221_X1 port map( B1 => n61761, B2 => n31, C1 => n61758, C2 => n23
                           , A => n5778, ZN => n5773);
   U3524 : NOR4_X1 port map( A1 => n5697, A2 => n5698, A3 => n5699, A4 => n5700
                           , ZN => n5669);
   U3525 : OAI221_X1 port map( B1 => n61749, B2 => n14, C1 => n61746, C2 => n6,
                           A => n5704, ZN => n5697);
   U3526 : OAI221_X1 port map( B1 => n5536, B2 => n1108, C1 => n5537, C2 => 
                           n1092, A => n5701, ZN => n5700);
   U3527 : OAI221_X1 port map( B1 => n61761, B2 => n30, C1 => n61758, C2 => n22
                           , A => n5703, ZN => n5698);
   U3528 : NOR4_X1 port map( A1 => n5622, A2 => n5623, A3 => n5624, A4 => n5625
                           , ZN => n5594);
   U3529 : OAI221_X1 port map( B1 => n61749, B2 => n13, C1 => n61746, C2 => n5,
                           A => n5629, ZN => n5622);
   U3530 : OAI221_X1 port map( B1 => n5536, B2 => n1107, C1 => n5537, C2 => 
                           n1091, A => n5626, ZN => n5625);
   U3531 : OAI221_X1 port map( B1 => n61761, B2 => n29, C1 => n61758, C2 => n21
                           , A => n5628, ZN => n5623);
   U3532 : NOR4_X1 port map( A1 => n5532, A2 => n5533, A3 => n5534, A4 => n5535
                           , ZN => n5463);
   U3533 : OAI221_X1 port map( B1 => n61749, B2 => n12, C1 => n61746, C2 => n4,
                           A => n5551, ZN => n5532);
   U3534 : OAI221_X1 port map( B1 => n5536, B2 => n1106, C1 => n5537, C2 => 
                           n1090, A => n5538, ZN => n5535);
   U3535 : OAI221_X1 port map( B1 => n61761, B2 => n28, C1 => n61758, C2 => n20
                           , A => n5546, ZN => n5533);
   U3536 : NOR4_X1 port map( A1 => n14432, A2 => n14433, A3 => n14434, A4 => 
                           n14435, ZN => n14404);
   U3537 : OAI221_X1 port map( B1 => n1330, B2 => n61271, C1 => n1341, C2 => 
                           n61268, A => n14439, ZN => n14432);
   U3538 : OAI221_X1 port map( B1 => n1402, B2 => n61283, C1 => n1378, C2 => 
                           n61280, A => n14438, ZN => n14433);
   U3539 : OAI221_X1 port map( B1 => n3324, B2 => n61295, C1 => n3300, C2 => 
                           n61292, A => n14437, ZN => n14434);
   U3540 : NOR4_X1 port map( A1 => n14357, A2 => n14358, A3 => n14359, A4 => 
                           n14360, ZN => n9913);
   U3541 : OAI221_X1 port map( B1 => n1329, B2 => n61271, C1 => n1340, C2 => 
                           n61268, A => n14364, ZN => n14357);
   U3542 : OAI221_X1 port map( B1 => n1401, B2 => n61283, C1 => n1377, C2 => 
                           n61280, A => n14363, ZN => n14358);
   U3543 : OAI221_X1 port map( B1 => n3323, B2 => n61295, C1 => n3299, C2 => 
                           n61292, A => n14362, ZN => n14359);
   U3544 : NOR4_X1 port map( A1 => n9866, A2 => n9867, A3 => n9868, A4 => n9869
                           , ZN => n9838);
   U3545 : OAI221_X1 port map( B1 => n1328, B2 => n61271, C1 => n1339, C2 => 
                           n61268, A => n9873, ZN => n9866);
   U3546 : OAI221_X1 port map( B1 => n1400, B2 => n61283, C1 => n1376, C2 => 
                           n61280, A => n9872, ZN => n9867);
   U3547 : OAI221_X1 port map( B1 => n3322, B2 => n61295, C1 => n3298, C2 => 
                           n61292, A => n9871, ZN => n9868);
   U3548 : NOR4_X1 port map( A1 => n9727, A2 => n9728, A3 => n9729, A4 => n9730
                           , ZN => n9699);
   U3549 : OAI221_X1 port map( B1 => n1362, B2 => n61271, C1 => n1327, C2 => 
                           n61268, A => n9734, ZN => n9727);
   U3550 : OAI221_X1 port map( B1 => n1399, B2 => n61283, C1 => n1375, C2 => 
                           n61280, A => n9733, ZN => n9728);
   U3551 : OAI221_X1 port map( B1 => n3321, B2 => n61295, C1 => n3297, C2 => 
                           n61292, A => n9732, ZN => n9729);
   U3552 : NOR4_X1 port map( A1 => n9652, A2 => n9653, A3 => n9654, A4 => n9655
                           , ZN => n9624);
   U3553 : OAI221_X1 port map( B1 => n1361, B2 => n61272, C1 => n1326, C2 => 
                           n61269, A => n9659, ZN => n9652);
   U3554 : OAI221_X1 port map( B1 => n1398, B2 => n61284, C1 => n1374, C2 => 
                           n61281, A => n9658, ZN => n9653);
   U3555 : OAI221_X1 port map( B1 => n3320, B2 => n61296, C1 => n3296, C2 => 
                           n61293, A => n9657, ZN => n9654);
   U3556 : NOR4_X1 port map( A1 => n9561, A2 => n9562, A3 => n9563, A4 => n9564
                           , ZN => n9533);
   U3557 : OAI221_X1 port map( B1 => n1360, B2 => n61272, C1 => n1325, C2 => 
                           n61269, A => n9568, ZN => n9561);
   U3558 : OAI221_X1 port map( B1 => n1397, B2 => n61284, C1 => n1373, C2 => 
                           n61281, A => n9567, ZN => n9562);
   U3559 : OAI221_X1 port map( B1 => n3319, B2 => n61296, C1 => n3295, C2 => 
                           n61293, A => n9566, ZN => n9563);
   U3560 : NOR4_X1 port map( A1 => n9486, A2 => n9487, A3 => n9488, A4 => n9489
                           , ZN => n9458);
   U3561 : OAI221_X1 port map( B1 => n1359, B2 => n61272, C1 => n1324, C2 => 
                           n61269, A => n9493, ZN => n9486);
   U3562 : OAI221_X1 port map( B1 => n1396, B2 => n61284, C1 => n1372, C2 => 
                           n61281, A => n9492, ZN => n9487);
   U3563 : OAI221_X1 port map( B1 => n3318, B2 => n61296, C1 => n3294, C2 => 
                           n61293, A => n9491, ZN => n9488);
   U3564 : NOR4_X1 port map( A1 => n9411, A2 => n9412, A3 => n9413, A4 => n9414
                           , ZN => n9383);
   U3565 : OAI221_X1 port map( B1 => n1358, B2 => n61272, C1 => n1323, C2 => 
                           n61269, A => n9418, ZN => n9411);
   U3566 : OAI221_X1 port map( B1 => n1395, B2 => n61284, C1 => n1371, C2 => 
                           n61281, A => n9417, ZN => n9412);
   U3567 : OAI221_X1 port map( B1 => n3317, B2 => n61296, C1 => n3293, C2 => 
                           n61293, A => n9416, ZN => n9413);
   U3568 : NOR4_X1 port map( A1 => n9272, A2 => n9273, A3 => n9274, A4 => n9275
                           , ZN => n9244);
   U3569 : OAI221_X1 port map( B1 => n1357, B2 => n61272, C1 => n1322, C2 => 
                           n61269, A => n9279, ZN => n9272);
   U3570 : OAI221_X1 port map( B1 => n1394, B2 => n61284, C1 => n1370, C2 => 
                           n61281, A => n9278, ZN => n9273);
   U3571 : OAI221_X1 port map( B1 => n3316, B2 => n61296, C1 => n3292, C2 => 
                           n61293, A => n9277, ZN => n9274);
   U3572 : NOR4_X1 port map( A1 => n9197, A2 => n9198, A3 => n9199, A4 => n9200
                           , ZN => n9169);
   U3573 : OAI221_X1 port map( B1 => n1356, B2 => n61272, C1 => n1321, C2 => 
                           n61269, A => n9204, ZN => n9197);
   U3574 : OAI221_X1 port map( B1 => n1393, B2 => n61284, C1 => n1369, C2 => 
                           n61281, A => n9203, ZN => n9198);
   U3575 : OAI221_X1 port map( B1 => n3315, B2 => n61296, C1 => n3291, C2 => 
                           n61293, A => n9202, ZN => n9199);
   U3576 : NOR4_X1 port map( A1 => n9122, A2 => n9123, A3 => n9124, A4 => n9125
                           , ZN => n9094);
   U3577 : OAI221_X1 port map( B1 => n1355, B2 => n61272, C1 => n1320, C2 => 
                           n61269, A => n9129, ZN => n9122);
   U3578 : OAI221_X1 port map( B1 => n1392, B2 => n61284, C1 => n1368, C2 => 
                           n61281, A => n9128, ZN => n9123);
   U3579 : OAI221_X1 port map( B1 => n3314, B2 => n61296, C1 => n3290, C2 => 
                           n61293, A => n9127, ZN => n9124);
   U3580 : NOR4_X1 port map( A1 => n9047, A2 => n9048, A3 => n9049, A4 => n9050
                           , ZN => n9019);
   U3581 : OAI221_X1 port map( B1 => n1354, B2 => n61272, C1 => n1319, C2 => 
                           n61269, A => n9054, ZN => n9047);
   U3582 : OAI221_X1 port map( B1 => n1391, B2 => n61284, C1 => n1367, C2 => 
                           n61281, A => n9053, ZN => n9048);
   U3583 : OAI221_X1 port map( B1 => n3313, B2 => n61296, C1 => n3289, C2 => 
                           n61293, A => n9052, ZN => n9049);
   U3584 : NOR4_X1 port map( A1 => n8972, A2 => n8973, A3 => n8974, A4 => n8975
                           , ZN => n8944);
   U3585 : OAI221_X1 port map( B1 => n1353, B2 => n61272, C1 => n1318, C2 => 
                           n61269, A => n8979, ZN => n8972);
   U3586 : OAI221_X1 port map( B1 => n1390, B2 => n61284, C1 => n1366, C2 => 
                           n61281, A => n8978, ZN => n8973);
   U3587 : OAI221_X1 port map( B1 => n3312, B2 => n61296, C1 => n3288, C2 => 
                           n61293, A => n8977, ZN => n8974);
   U3588 : NOR4_X1 port map( A1 => n8897, A2 => n8898, A3 => n8899, A4 => n8900
                           , ZN => n8869);
   U3589 : OAI221_X1 port map( B1 => n1352, B2 => n61272, C1 => n1317, C2 => 
                           n61269, A => n8904, ZN => n8897);
   U3590 : OAI221_X1 port map( B1 => n1389, B2 => n61284, C1 => n1365, C2 => 
                           n61281, A => n8903, ZN => n8898);
   U3591 : OAI221_X1 port map( B1 => n3311, B2 => n61296, C1 => n3287, C2 => 
                           n61293, A => n8902, ZN => n8899);
   U3592 : NOR4_X1 port map( A1 => n8822, A2 => n8823, A3 => n8824, A4 => n8825
                           , ZN => n8794);
   U3593 : OAI221_X1 port map( B1 => n1351, B2 => n61272, C1 => n1316, C2 => 
                           n61269, A => n8829, ZN => n8822);
   U3594 : OAI221_X1 port map( B1 => n1388, B2 => n61284, C1 => n1364, C2 => 
                           n61281, A => n8828, ZN => n8823);
   U3595 : OAI221_X1 port map( B1 => n3310, B2 => n61296, C1 => n3286, C2 => 
                           n61293, A => n8827, ZN => n8824);
   U3596 : NOR4_X1 port map( A1 => n8747, A2 => n8748, A3 => n8749, A4 => n8750
                           , ZN => n8719);
   U3597 : OAI221_X1 port map( B1 => n1350, B2 => n61272, C1 => n1315, C2 => 
                           n61269, A => n8754, ZN => n8747);
   U3598 : OAI221_X1 port map( B1 => n1387, B2 => n61284, C1 => n1363, C2 => 
                           n61281, A => n8753, ZN => n8748);
   U3599 : OAI221_X1 port map( B1 => n3309, B2 => n61296, C1 => n3285, C2 => 
                           n61293, A => n8752, ZN => n8749);
   U3600 : NOR4_X1 port map( A1 => n15063, A2 => n15064, A3 => n15065, A4 => 
                           n15066, ZN => n15027);
   U3601 : OAI221_X1 port map( B1 => n1338, B2 => n61271, C1 => n1349, C2 => 
                           n61268, A => n15071, ZN => n15063);
   U3602 : OAI221_X1 port map( B1 => n1410, B2 => n61283, C1 => n1386, C2 => 
                           n61280, A => n15070, ZN => n15064);
   U3603 : OAI221_X1 port map( B1 => n3332, B2 => n61295, C1 => n3308, C2 => 
                           n61292, A => n15069, ZN => n15065);
   U3604 : NOR4_X1 port map( A1 => n14957, A2 => n14958, A3 => n14959, A4 => 
                           n14960, ZN => n14929);
   U3605 : OAI221_X1 port map( B1 => n1337, B2 => n61271, C1 => n1348, C2 => 
                           n61268, A => n14964, ZN => n14957);
   U3606 : OAI221_X1 port map( B1 => n1409, B2 => n61283, C1 => n1385, C2 => 
                           n61280, A => n14963, ZN => n14958);
   U3607 : OAI221_X1 port map( B1 => n3331, B2 => n61295, C1 => n3307, C2 => 
                           n61292, A => n14962, ZN => n14959);
   U3608 : NOR4_X1 port map( A1 => n14882, A2 => n14883, A3 => n14884, A4 => 
                           n14885, ZN => n14854);
   U3609 : OAI221_X1 port map( B1 => n1336, B2 => n61271, C1 => n1347, C2 => 
                           n61268, A => n14889, ZN => n14882);
   U3610 : OAI221_X1 port map( B1 => n1408, B2 => n61283, C1 => n1384, C2 => 
                           n61280, A => n14888, ZN => n14883);
   U3611 : OAI221_X1 port map( B1 => n3330, B2 => n61295, C1 => n3306, C2 => 
                           n61292, A => n14887, ZN => n14884);
   U3612 : NOR4_X1 port map( A1 => n14807, A2 => n14808, A3 => n14809, A4 => 
                           n14810, ZN => n14779);
   U3613 : OAI221_X1 port map( B1 => n1335, B2 => n61271, C1 => n1346, C2 => 
                           n61268, A => n14814, ZN => n14807);
   U3614 : OAI221_X1 port map( B1 => n1407, B2 => n61283, C1 => n1383, C2 => 
                           n61280, A => n14813, ZN => n14808);
   U3615 : OAI221_X1 port map( B1 => n3329, B2 => n61295, C1 => n3305, C2 => 
                           n61292, A => n14812, ZN => n14809);
   U3616 : NOR4_X1 port map( A1 => n14732, A2 => n14733, A3 => n14734, A4 => 
                           n14735, ZN => n14704);
   U3617 : OAI221_X1 port map( B1 => n1334, B2 => n61271, C1 => n1345, C2 => 
                           n61268, A => n14739, ZN => n14732);
   U3618 : OAI221_X1 port map( B1 => n1406, B2 => n61283, C1 => n1382, C2 => 
                           n61280, A => n14738, ZN => n14733);
   U3619 : OAI221_X1 port map( B1 => n3328, B2 => n61295, C1 => n3304, C2 => 
                           n61292, A => n14737, ZN => n14734);
   U3620 : NOR4_X1 port map( A1 => n14657, A2 => n14658, A3 => n14659, A4 => 
                           n14660, ZN => n14629);
   U3621 : OAI221_X1 port map( B1 => n1333, B2 => n61271, C1 => n1344, C2 => 
                           n61268, A => n14664, ZN => n14657);
   U3622 : OAI221_X1 port map( B1 => n1405, B2 => n61283, C1 => n1381, C2 => 
                           n61280, A => n14663, ZN => n14658);
   U3623 : OAI221_X1 port map( B1 => n3327, B2 => n61295, C1 => n3303, C2 => 
                           n61292, A => n14662, ZN => n14659);
   U3624 : NOR4_X1 port map( A1 => n14582, A2 => n14583, A3 => n14584, A4 => 
                           n14585, ZN => n14554);
   U3625 : OAI221_X1 port map( B1 => n1332, B2 => n61271, C1 => n1343, C2 => 
                           n61268, A => n14589, ZN => n14582);
   U3626 : OAI221_X1 port map( B1 => n1404, B2 => n61283, C1 => n1380, C2 => 
                           n61280, A => n14588, ZN => n14583);
   U3627 : OAI221_X1 port map( B1 => n3326, B2 => n61295, C1 => n3302, C2 => 
                           n61292, A => n14587, ZN => n14584);
   U3628 : NOR4_X1 port map( A1 => n14507, A2 => n14508, A3 => n14509, A4 => 
                           n14510, ZN => n14479);
   U3629 : OAI221_X1 port map( B1 => n1331, B2 => n61271, C1 => n1342, C2 => 
                           n61268, A => n14514, ZN => n14507);
   U3630 : OAI221_X1 port map( B1 => n1403, B2 => n61283, C1 => n1379, C2 => 
                           n61280, A => n14513, ZN => n14508);
   U3631 : OAI221_X1 port map( B1 => n3325, B2 => n61295, C1 => n3301, C2 => 
                           n61292, A => n14512, ZN => n14509);
   U3632 : NOR4_X1 port map( A1 => n8672, A2 => n8673, A3 => n8674, A4 => n8675
                           , ZN => n8644);
   U3633 : OAI221_X1 port map( B1 => n19, B2 => n61273, C1 => n11, C2 => n61270
                           , A => n8679, ZN => n8672);
   U3634 : OAI221_X1 port map( B1 => n35, B2 => n61285, C1 => n27, C2 => n61282
                           , A => n8678, ZN => n8673);
   U3635 : OAI221_X1 port map( B1 => n1069, B2 => n61297, C1 => n1061, C2 => 
                           n61294, A => n8677, ZN => n8674);
   U3636 : NOR4_X1 port map( A1 => n8597, A2 => n8598, A3 => n8599, A4 => n8600
                           , ZN => n8569);
   U3637 : OAI221_X1 port map( B1 => n18, B2 => n61273, C1 => n10, C2 => n61270
                           , A => n8604, ZN => n8597);
   U3638 : OAI221_X1 port map( B1 => n34, B2 => n61285, C1 => n26, C2 => n61282
                           , A => n8603, ZN => n8598);
   U3639 : OAI221_X1 port map( B1 => n1068, B2 => n61297, C1 => n1060, C2 => 
                           n61294, A => n8602, ZN => n8599);
   U3640 : NOR4_X1 port map( A1 => n8522, A2 => n8523, A3 => n8524, A4 => n8525
                           , ZN => n8494);
   U3641 : OAI221_X1 port map( B1 => n17, B2 => n61273, C1 => n9, C2 => n61270,
                           A => n8529, ZN => n8522);
   U3642 : OAI221_X1 port map( B1 => n33, B2 => n61285, C1 => n25, C2 => n61282
                           , A => n8528, ZN => n8523);
   U3643 : OAI221_X1 port map( B1 => n1067, B2 => n61297, C1 => n1059, C2 => 
                           n61294, A => n8527, ZN => n8524);
   U3644 : NOR4_X1 port map( A1 => n8447, A2 => n8448, A3 => n8449, A4 => n8450
                           , ZN => n8419);
   U3645 : OAI221_X1 port map( B1 => n16, B2 => n61273, C1 => n8, C2 => n61270,
                           A => n8454, ZN => n8447);
   U3646 : OAI221_X1 port map( B1 => n32, B2 => n61285, C1 => n24, C2 => n61282
                           , A => n8453, ZN => n8448);
   U3647 : OAI221_X1 port map( B1 => n1066, B2 => n61297, C1 => n1058, C2 => 
                           n61294, A => n8452, ZN => n8449);
   U3648 : NOR4_X1 port map( A1 => n8372, A2 => n8373, A3 => n8374, A4 => n8375
                           , ZN => n8344);
   U3649 : OAI221_X1 port map( B1 => n15, B2 => n61273, C1 => n7, C2 => n61270,
                           A => n8379, ZN => n8372);
   U3650 : OAI221_X1 port map( B1 => n31, B2 => n61285, C1 => n23, C2 => n61282
                           , A => n8378, ZN => n8373);
   U3651 : OAI221_X1 port map( B1 => n1065, B2 => n61297, C1 => n1057, C2 => 
                           n61294, A => n8377, ZN => n8374);
   U3652 : NOR4_X1 port map( A1 => n8297, A2 => n8298, A3 => n8299, A4 => n8300
                           , ZN => n8269);
   U3653 : OAI221_X1 port map( B1 => n14, B2 => n61273, C1 => n6, C2 => n61270,
                           A => n8304, ZN => n8297);
   U3654 : OAI221_X1 port map( B1 => n30, B2 => n61285, C1 => n22, C2 => n61282
                           , A => n8303, ZN => n8298);
   U3655 : OAI221_X1 port map( B1 => n1064, B2 => n61297, C1 => n1056, C2 => 
                           n61294, A => n8302, ZN => n8299);
   U3656 : NOR4_X1 port map( A1 => n8222, A2 => n8223, A3 => n8224, A4 => n8225
                           , ZN => n8194);
   U3657 : OAI221_X1 port map( B1 => n13, B2 => n61273, C1 => n5, C2 => n61270,
                           A => n8229, ZN => n8222);
   U3658 : OAI221_X1 port map( B1 => n29, B2 => n61285, C1 => n21, C2 => n61282
                           , A => n8228, ZN => n8223);
   U3659 : OAI221_X1 port map( B1 => n1063, B2 => n61297, C1 => n1055, C2 => 
                           n61294, A => n8227, ZN => n8224);
   U3660 : NOR4_X1 port map( A1 => n8130, A2 => n8131, A3 => n8132, A4 => n8133
                           , ZN => n8051);
   U3661 : OAI221_X1 port map( B1 => n12, B2 => n61273, C1 => n4, C2 => n61270,
                           A => n8151, ZN => n8130);
   U3662 : OAI221_X1 port map( B1 => n28, B2 => n61285, C1 => n20, C2 => n61282
                           , A => n8146, ZN => n8131);
   U3663 : OAI221_X1 port map( B1 => n1062, B2 => n61297, C1 => n1054, C2 => 
                           n61294, A => n8141, ZN => n8132);
   U3664 : NOR2_X1 port map( A1 => n5282, A2 => ADDR_WR(0), ZN => n15261);
   U3665 : NOR2_X1 port map( A1 => ADDR_WR(3), A2 => ADDR_WR(2), ZN => n15279);
   U3666 : NOR2_X1 port map( A1 => n5283, A2 => ADDR_WR(1), ZN => n15259);
   U3667 : NAND2_X1 port map( A1 => n15126, A2 => n15127, ZN => n15094);
   U3668 : INV_X1 port map( A => ADDR_RD2(0), ZN => n5361);
   U3669 : INV_X1 port map( A => ADDR_RD1(0), ZN => n5353);
   U3670 : INV_X1 port map( A => ADDR_RD2(1), ZN => n5360);
   U3671 : INV_X1 port map( A => ADDR_RD1(1), ZN => n5352);
   U3672 : INV_X1 port map( A => ADDR_RD2(2), ZN => n5359);
   U3673 : INV_X1 port map( A => ADDR_RD1(2), ZN => n5351);
   U3674 : OAI22_X1 port map( A1 => n60655, A2 => n61142, B1 => n4288, B2 => 
                           n60650, ZN => n13245);
   U3675 : OAI22_X1 port map( A1 => n60656, A2 => n61156, B1 => n4287, B2 => 
                           n60650, ZN => n13246);
   U3676 : OAI22_X1 port map( A1 => n60656, A2 => n61170, B1 => n4286, B2 => 
                           n60650, ZN => n13247);
   U3677 : OAI22_X1 port map( A1 => n60656, A2 => n61184, B1 => n4285, B2 => 
                           n60650, ZN => n13248);
   U3678 : OAI22_X1 port map( A1 => n60656, A2 => n61198, B1 => n4284, B2 => 
                           n15149, ZN => n13249);
   U3679 : OAI22_X1 port map( A1 => n60656, A2 => n61212, B1 => n4283, B2 => 
                           n15149, ZN => n13250);
   U3680 : OAI22_X1 port map( A1 => n60657, A2 => n61226, B1 => n4282, B2 => 
                           n15149, ZN => n13251);
   U3681 : OAI22_X1 port map( A1 => n60657, A2 => n61249, B1 => n4281, B2 => 
                           n15149, ZN => n13252);
   U3682 : OAI22_X1 port map( A1 => n60646, A2 => n61142, B1 => n4280, B2 => 
                           n60641, ZN => n13213);
   U3683 : OAI22_X1 port map( A1 => n60647, A2 => n61156, B1 => n4279, B2 => 
                           n60641, ZN => n13214);
   U3684 : OAI22_X1 port map( A1 => n60647, A2 => n61170, B1 => n4278, B2 => 
                           n60641, ZN => n13215);
   U3685 : OAI22_X1 port map( A1 => n60647, A2 => n61184, B1 => n4277, B2 => 
                           n60641, ZN => n13216);
   U3686 : OAI22_X1 port map( A1 => n60647, A2 => n61198, B1 => n4276, B2 => 
                           n15150, ZN => n13217);
   U3687 : OAI22_X1 port map( A1 => n60647, A2 => n61212, B1 => n4275, B2 => 
                           n15150, ZN => n13218);
   U3688 : OAI22_X1 port map( A1 => n60648, A2 => n61226, B1 => n4274, B2 => 
                           n15150, ZN => n13219);
   U3689 : OAI22_X1 port map( A1 => n60648, A2 => n61249, B1 => n4273, B2 => 
                           n15150, ZN => n13220);
   U3690 : OAI22_X1 port map( A1 => n60556, A2 => n61143, B1 => n4240, B2 => 
                           n60551, ZN => n12893);
   U3691 : OAI22_X1 port map( A1 => n60557, A2 => n61157, B1 => n4239, B2 => 
                           n60551, ZN => n12894);
   U3692 : OAI22_X1 port map( A1 => n60557, A2 => n61171, B1 => n4238, B2 => 
                           n60551, ZN => n12895);
   U3693 : OAI22_X1 port map( A1 => n60557, A2 => n61185, B1 => n4237, B2 => 
                           n60551, ZN => n12896);
   U3694 : OAI22_X1 port map( A1 => n60557, A2 => n61199, B1 => n4236, B2 => 
                           n15160, ZN => n12897);
   U3695 : OAI22_X1 port map( A1 => n60547, A2 => n61143, B1 => n4235, B2 => 
                           n60542, ZN => n12861);
   U3696 : OAI22_X1 port map( A1 => n60548, A2 => n61157, B1 => n4234, B2 => 
                           n60542, ZN => n12862);
   U3697 : OAI22_X1 port map( A1 => n60548, A2 => n61171, B1 => n4233, B2 => 
                           n60542, ZN => n12863);
   U3698 : OAI22_X1 port map( A1 => n60548, A2 => n61185, B1 => n4232, B2 => 
                           n60542, ZN => n12864);
   U3699 : OAI22_X1 port map( A1 => n60548, A2 => n61199, B1 => n4231, B2 => 
                           n15161, ZN => n12865);
   U3700 : OAI22_X1 port map( A1 => n60548, A2 => n61213, B1 => n4230, B2 => 
                           n15161, ZN => n12866);
   U3701 : OAI22_X1 port map( A1 => n60549, A2 => n61227, B1 => n4229, B2 => 
                           n15161, ZN => n12867);
   U3702 : OAI22_X1 port map( A1 => n60549, A2 => n61250, B1 => n4228, B2 => 
                           n15161, ZN => n12868);
   U3703 : OAI22_X1 port map( A1 => n60538, A2 => n61143, B1 => n4227, B2 => 
                           n60533, ZN => n12829);
   U3704 : OAI22_X1 port map( A1 => n60539, A2 => n61157, B1 => n4226, B2 => 
                           n60533, ZN => n12830);
   U3705 : OAI22_X1 port map( A1 => n60539, A2 => n61171, B1 => n4225, B2 => 
                           n60533, ZN => n12831);
   U3706 : OAI22_X1 port map( A1 => n60539, A2 => n61185, B1 => n4224, B2 => 
                           n60533, ZN => n12832);
   U3707 : OAI22_X1 port map( A1 => n60539, A2 => n61199, B1 => n4223, B2 => 
                           n15162, ZN => n12833);
   U3708 : OAI22_X1 port map( A1 => n60539, A2 => n61213, B1 => n4222, B2 => 
                           n15162, ZN => n12834);
   U3709 : OAI22_X1 port map( A1 => n60540, A2 => n61227, B1 => n4221, B2 => 
                           n15162, ZN => n12835);
   U3710 : OAI22_X1 port map( A1 => n60540, A2 => n61250, B1 => n4220, B2 => 
                           n15162, ZN => n12836);
   U3711 : OAI22_X1 port map( A1 => n60484, A2 => n61144, B1 => n4219, B2 => 
                           n60479, ZN => n12637);
   U3712 : OAI22_X1 port map( A1 => n60485, A2 => n61158, B1 => n4218, B2 => 
                           n60479, ZN => n12638);
   U3713 : OAI22_X1 port map( A1 => n60485, A2 => n61172, B1 => n4217, B2 => 
                           n60479, ZN => n12639);
   U3714 : OAI22_X1 port map( A1 => n60485, A2 => n61186, B1 => n4216, B2 => 
                           n60479, ZN => n12640);
   U3715 : OAI22_X1 port map( A1 => n60485, A2 => n61200, B1 => n4215, B2 => 
                           n15169, ZN => n12641);
   U3716 : OAI22_X1 port map( A1 => n60485, A2 => n61214, B1 => n4214, B2 => 
                           n15169, ZN => n12642);
   U3717 : OAI22_X1 port map( A1 => n60486, A2 => n61228, B1 => n4213, B2 => 
                           n15169, ZN => n12643);
   U3718 : OAI22_X1 port map( A1 => n60486, A2 => n61251, B1 => n4212, B2 => 
                           n15169, ZN => n12644);
   U3719 : OAI22_X1 port map( A1 => n60925, A2 => n61140, B1 => n4163, B2 => 
                           n60920, ZN => n14205);
   U3720 : OAI22_X1 port map( A1 => n60926, A2 => n61154, B1 => n4162, B2 => 
                           n60920, ZN => n14206);
   U3721 : OAI22_X1 port map( A1 => n60926, A2 => n61168, B1 => n4161, B2 => 
                           n60920, ZN => n14207);
   U3722 : OAI22_X1 port map( A1 => n60926, A2 => n61182, B1 => n4160, B2 => 
                           n60920, ZN => n14208);
   U3723 : OAI22_X1 port map( A1 => n60926, A2 => n61196, B1 => n4159, B2 => 
                           n15102, ZN => n14209);
   U3724 : OAI22_X1 port map( A1 => n60926, A2 => n61210, B1 => n4158, B2 => 
                           n15102, ZN => n14210);
   U3725 : OAI22_X1 port map( A1 => n60927, A2 => n61224, B1 => n4157, B2 => 
                           n15102, ZN => n14211);
   U3726 : OAI22_X1 port map( A1 => n60927, A2 => n61247, B1 => n4156, B2 => 
                           n15102, ZN => n14212);
   U3727 : OAI22_X1 port map( A1 => n60916, A2 => n61140, B1 => n4155, B2 => 
                           n60911, ZN => n14173);
   U3728 : OAI22_X1 port map( A1 => n60917, A2 => n61154, B1 => n4154, B2 => 
                           n60911, ZN => n14174);
   U3729 : OAI22_X1 port map( A1 => n60917, A2 => n61168, B1 => n4153, B2 => 
                           n60911, ZN => n14175);
   U3730 : OAI22_X1 port map( A1 => n60917, A2 => n61182, B1 => n4152, B2 => 
                           n60911, ZN => n14176);
   U3731 : OAI22_X1 port map( A1 => n60917, A2 => n61196, B1 => n4151, B2 => 
                           n15104, ZN => n14177);
   U3732 : OAI22_X1 port map( A1 => n60917, A2 => n61210, B1 => n4150, B2 => 
                           n15104, ZN => n14178);
   U3733 : OAI22_X1 port map( A1 => n60918, A2 => n61224, B1 => n4149, B2 => 
                           n15104, ZN => n14179);
   U3734 : OAI22_X1 port map( A1 => n60918, A2 => n61247, B1 => n4148, B2 => 
                           n15104, ZN => n14180);
   U3735 : OAI22_X1 port map( A1 => n60889, A2 => n61140, B1 => n4147, B2 => 
                           n60884, ZN => n14077);
   U3736 : OAI22_X1 port map( A1 => n60890, A2 => n61154, B1 => n4146, B2 => 
                           n60884, ZN => n14078);
   U3737 : OAI22_X1 port map( A1 => n60890, A2 => n61168, B1 => n4145, B2 => 
                           n60884, ZN => n14079);
   U3738 : OAI22_X1 port map( A1 => n60890, A2 => n61182, B1 => n4144, B2 => 
                           n60884, ZN => n14080);
   U3739 : OAI22_X1 port map( A1 => n60890, A2 => n61196, B1 => n4143, B2 => 
                           n15110, ZN => n14081);
   U3740 : OAI22_X1 port map( A1 => n60890, A2 => n61210, B1 => n4142, B2 => 
                           n15110, ZN => n14082);
   U3741 : OAI22_X1 port map( A1 => n60891, A2 => n61224, B1 => n4141, B2 => 
                           n15110, ZN => n14083);
   U3742 : OAI22_X1 port map( A1 => n60891, A2 => n61247, B1 => n4140, B2 => 
                           n15110, ZN => n14084);
   U3743 : OAI22_X1 port map( A1 => n60880, A2 => n61140, B1 => n4139, B2 => 
                           n60875, ZN => n14045);
   U3744 : OAI22_X1 port map( A1 => n60881, A2 => n61154, B1 => n4138, B2 => 
                           n60875, ZN => n14046);
   U3745 : OAI22_X1 port map( A1 => n60881, A2 => n61168, B1 => n4137, B2 => 
                           n60875, ZN => n14047);
   U3746 : OAI22_X1 port map( A1 => n60881, A2 => n61182, B1 => n4136, B2 => 
                           n60875, ZN => n14048);
   U3747 : OAI22_X1 port map( A1 => n60881, A2 => n61196, B1 => n4135, B2 => 
                           n15112, ZN => n14049);
   U3748 : OAI22_X1 port map( A1 => n60881, A2 => n61210, B1 => n4134, B2 => 
                           n15112, ZN => n14050);
   U3749 : OAI22_X1 port map( A1 => n60882, A2 => n61224, B1 => n4133, B2 => 
                           n15112, ZN => n14051);
   U3750 : OAI22_X1 port map( A1 => n60882, A2 => n61247, B1 => n4132, B2 => 
                           n15112, ZN => n14052);
   U3751 : OAI22_X1 port map( A1 => n60853, A2 => n61141, B1 => n4131, B2 => 
                           n60848, ZN => n13949);
   U3752 : OAI22_X1 port map( A1 => n60854, A2 => n61155, B1 => n4130, B2 => 
                           n60848, ZN => n13950);
   U3753 : OAI22_X1 port map( A1 => n60854, A2 => n61169, B1 => n4129, B2 => 
                           n60848, ZN => n13951);
   U3754 : OAI22_X1 port map( A1 => n60854, A2 => n61183, B1 => n4128, B2 => 
                           n60848, ZN => n13952);
   U3755 : OAI22_X1 port map( A1 => n60854, A2 => n61197, B1 => n4127, B2 => 
                           n15118, ZN => n13953);
   U3756 : OAI22_X1 port map( A1 => n60854, A2 => n61211, B1 => n4126, B2 => 
                           n15118, ZN => n13954);
   U3757 : OAI22_X1 port map( A1 => n60855, A2 => n61225, B1 => n4125, B2 => 
                           n15118, ZN => n13955);
   U3758 : OAI22_X1 port map( A1 => n60855, A2 => n61248, B1 => n4124, B2 => 
                           n15118, ZN => n13956);
   U3759 : OAI22_X1 port map( A1 => n60844, A2 => n61141, B1 => n4123, B2 => 
                           n60839, ZN => n13917);
   U3760 : OAI22_X1 port map( A1 => n60845, A2 => n61155, B1 => n4122, B2 => 
                           n60839, ZN => n13918);
   U3761 : OAI22_X1 port map( A1 => n60845, A2 => n61169, B1 => n4121, B2 => 
                           n60839, ZN => n13919);
   U3762 : OAI22_X1 port map( A1 => n60845, A2 => n61183, B1 => n4120, B2 => 
                           n60839, ZN => n13920);
   U3763 : OAI22_X1 port map( A1 => n60845, A2 => n61197, B1 => n4119, B2 => 
                           n15120, ZN => n13921);
   U3764 : OAI22_X1 port map( A1 => n60845, A2 => n61211, B1 => n4118, B2 => 
                           n15120, ZN => n13922);
   U3765 : OAI22_X1 port map( A1 => n60846, A2 => n61225, B1 => n4117, B2 => 
                           n15120, ZN => n13923);
   U3766 : OAI22_X1 port map( A1 => n60846, A2 => n61248, B1 => n4116, B2 => 
                           n15120, ZN => n13924);
   U3767 : OAI22_X1 port map( A1 => n60349, A2 => n61145, B1 => n4075, B2 => 
                           n60344, ZN => n12157);
   U3768 : OAI22_X1 port map( A1 => n60350, A2 => n61159, B1 => n4074, B2 => 
                           n60344, ZN => n12158);
   U3769 : OAI22_X1 port map( A1 => n60350, A2 => n61173, B1 => n4073, B2 => 
                           n60344, ZN => n12159);
   U3770 : OAI22_X1 port map( A1 => n60350, A2 => n61187, B1 => n4072, B2 => 
                           n60344, ZN => n12160);
   U3771 : OAI22_X1 port map( A1 => n60350, A2 => n61201, B1 => n4071, B2 => 
                           n15192, ZN => n12161);
   U3772 : OAI22_X1 port map( A1 => n60350, A2 => n61215, B1 => n4070, B2 => 
                           n15192, ZN => n12162);
   U3773 : OAI22_X1 port map( A1 => n60351, A2 => n61229, B1 => n4069, B2 => 
                           n15192, ZN => n12163);
   U3774 : OAI22_X1 port map( A1 => n60351, A2 => n61252, B1 => n4068, B2 => 
                           n15192, ZN => n12164);
   U3775 : OAI22_X1 port map( A1 => n60340, A2 => n61145, B1 => n4067, B2 => 
                           n60335, ZN => n12125);
   U3776 : OAI22_X1 port map( A1 => n60341, A2 => n61159, B1 => n4066, B2 => 
                           n60335, ZN => n12126);
   U3777 : OAI22_X1 port map( A1 => n60341, A2 => n61173, B1 => n4065, B2 => 
                           n60335, ZN => n12127);
   U3778 : OAI22_X1 port map( A1 => n60341, A2 => n61187, B1 => n4064, B2 => 
                           n60335, ZN => n12128);
   U3779 : OAI22_X1 port map( A1 => n60341, A2 => n61201, B1 => n4063, B2 => 
                           n15193, ZN => n12129);
   U3780 : OAI22_X1 port map( A1 => n60341, A2 => n61215, B1 => n4062, B2 => 
                           n15193, ZN => n12130);
   U3781 : OAI22_X1 port map( A1 => n60342, A2 => n61229, B1 => n4061, B2 => 
                           n15193, ZN => n12131);
   U3782 : OAI22_X1 port map( A1 => n60342, A2 => n61252, B1 => n4060, B2 => 
                           n15193, ZN => n12132);
   U3783 : OAI22_X1 port map( A1 => n60277, A2 => n61146, B1 => n4059, B2 => 
                           n60272, ZN => n11901);
   U3784 : OAI22_X1 port map( A1 => n60278, A2 => n61160, B1 => n4058, B2 => 
                           n60272, ZN => n11902);
   U3785 : OAI22_X1 port map( A1 => n60278, A2 => n61174, B1 => n4057, B2 => 
                           n60272, ZN => n11903);
   U3786 : OAI22_X1 port map( A1 => n60278, A2 => n61188, B1 => n4056, B2 => 
                           n60272, ZN => n11904);
   U3787 : OAI22_X1 port map( A1 => n60278, A2 => n61202, B1 => n4055, B2 => 
                           n15200, ZN => n11905);
   U3788 : OAI22_X1 port map( A1 => n60278, A2 => n61216, B1 => n4054, B2 => 
                           n15200, ZN => n11906);
   U3789 : OAI22_X1 port map( A1 => n60279, A2 => n61230, B1 => n4053, B2 => 
                           n15200, ZN => n11907);
   U3790 : OAI22_X1 port map( A1 => n60279, A2 => n61253, B1 => n4052, B2 => 
                           n15200, ZN => n11908);
   U3791 : OAI22_X1 port map( A1 => n60268, A2 => n61146, B1 => n4051, B2 => 
                           n60263, ZN => n11869);
   U3792 : OAI22_X1 port map( A1 => n60269, A2 => n61160, B1 => n4050, B2 => 
                           n60263, ZN => n11870);
   U3793 : OAI22_X1 port map( A1 => n60269, A2 => n61174, B1 => n4049, B2 => 
                           n60263, ZN => n11871);
   U3794 : OAI22_X1 port map( A1 => n60269, A2 => n61188, B1 => n4048, B2 => 
                           n60263, ZN => n11872);
   U3795 : OAI22_X1 port map( A1 => n60269, A2 => n61202, B1 => n4047, B2 => 
                           n15201, ZN => n11873);
   U3796 : OAI22_X1 port map( A1 => n60269, A2 => n61216, B1 => n4046, B2 => 
                           n15201, ZN => n11874);
   U3797 : OAI22_X1 port map( A1 => n60270, A2 => n61230, B1 => n4045, B2 => 
                           n15201, ZN => n11875);
   U3798 : OAI22_X1 port map( A1 => n60270, A2 => n61253, B1 => n4044, B2 => 
                           n15201, ZN => n11876);
   U3799 : OAI22_X1 port map( A1 => n60160, A2 => n61147, B1 => n4027, B2 => 
                           n60155, ZN => n11485);
   U3800 : OAI22_X1 port map( A1 => n60161, A2 => n61161, B1 => n4026, B2 => 
                           n60155, ZN => n11486);
   U3801 : OAI22_X1 port map( A1 => n60161, A2 => n61175, B1 => n4025, B2 => 
                           n60155, ZN => n11487);
   U3802 : OAI22_X1 port map( A1 => n60161, A2 => n61189, B1 => n4024, B2 => 
                           n60155, ZN => n11488);
   U3803 : OAI22_X1 port map( A1 => n60161, A2 => n61203, B1 => n4023, B2 => 
                           n15222, ZN => n11489);
   U3804 : OAI22_X1 port map( A1 => n60161, A2 => n61217, B1 => n4022, B2 => 
                           n15222, ZN => n11490);
   U3805 : OAI22_X1 port map( A1 => n60162, A2 => n61231, B1 => n4021, B2 => 
                           n15222, ZN => n11491);
   U3806 : OAI22_X1 port map( A1 => n60162, A2 => n61254, B1 => n4020, B2 => 
                           n15222, ZN => n11492);
   U3807 : OAI22_X1 port map( A1 => n60151, A2 => n61147, B1 => n4019, B2 => 
                           n60146, ZN => n11453);
   U3808 : OAI22_X1 port map( A1 => n60152, A2 => n61161, B1 => n4018, B2 => 
                           n60146, ZN => n11454);
   U3809 : OAI22_X1 port map( A1 => n60152, A2 => n61175, B1 => n4017, B2 => 
                           n60146, ZN => n11455);
   U3810 : OAI22_X1 port map( A1 => n60152, A2 => n61189, B1 => n4016, B2 => 
                           n60146, ZN => n11456);
   U3811 : OAI22_X1 port map( A1 => n60152, A2 => n61203, B1 => n4015, B2 => 
                           n15223, ZN => n11457);
   U3812 : OAI22_X1 port map( A1 => n60152, A2 => n61217, B1 => n4014, B2 => 
                           n15223, ZN => n11458);
   U3813 : OAI22_X1 port map( A1 => n60153, A2 => n61231, B1 => n4013, B2 => 
                           n15223, ZN => n11459);
   U3814 : OAI22_X1 port map( A1 => n60153, A2 => n61254, B1 => n4012, B2 => 
                           n15223, ZN => n11460);
   U3815 : OAI22_X1 port map( A1 => n60808, A2 => n61141, B1 => n4011, B2 => 
                           n60803, ZN => n13789);
   U3816 : OAI22_X1 port map( A1 => n60809, A2 => n61155, B1 => n4010, B2 => 
                           n60803, ZN => n13790);
   U3817 : OAI22_X1 port map( A1 => n60809, A2 => n61169, B1 => n4009, B2 => 
                           n60803, ZN => n13791);
   U3818 : OAI22_X1 port map( A1 => n60809, A2 => n61183, B1 => n4008, B2 => 
                           n60803, ZN => n13792);
   U3819 : OAI22_X1 port map( A1 => n60809, A2 => n61197, B1 => n4007, B2 => 
                           n15130, ZN => n13793);
   U3820 : OAI22_X1 port map( A1 => n60809, A2 => n61211, B1 => n4006, B2 => 
                           n15130, ZN => n13794);
   U3821 : OAI22_X1 port map( A1 => n60810, A2 => n61225, B1 => n4005, B2 => 
                           n15130, ZN => n13795);
   U3822 : OAI22_X1 port map( A1 => n60810, A2 => n61248, B1 => n4004, B2 => 
                           n15130, ZN => n13796);
   U3823 : OAI22_X1 port map( A1 => n60799, A2 => n61141, B1 => n4003, B2 => 
                           n60794, ZN => n13757);
   U3824 : OAI22_X1 port map( A1 => n60800, A2 => n61155, B1 => n4002, B2 => 
                           n60794, ZN => n13758);
   U3825 : OAI22_X1 port map( A1 => n60800, A2 => n61169, B1 => n4001, B2 => 
                           n60794, ZN => n13759);
   U3826 : OAI22_X1 port map( A1 => n60800, A2 => n61183, B1 => n4000, B2 => 
                           n60794, ZN => n13760);
   U3827 : OAI22_X1 port map( A1 => n60800, A2 => n61197, B1 => n3999, B2 => 
                           n15131, ZN => n13761);
   U3828 : OAI22_X1 port map( A1 => n60800, A2 => n61211, B1 => n3998, B2 => 
                           n15131, ZN => n13762);
   U3829 : OAI22_X1 port map( A1 => n60801, A2 => n61225, B1 => n3997, B2 => 
                           n15131, ZN => n13763);
   U3830 : OAI22_X1 port map( A1 => n60801, A2 => n61248, B1 => n3996, B2 => 
                           n15131, ZN => n13764);
   U3831 : OAI22_X1 port map( A1 => n60682, A2 => n61142, B1 => n3955, B2 => 
                           n60677, ZN => n13341);
   U3832 : OAI22_X1 port map( A1 => n60683, A2 => n61156, B1 => n3954, B2 => 
                           n60677, ZN => n13342);
   U3833 : OAI22_X1 port map( A1 => n60683, A2 => n61170, B1 => n3953, B2 => 
                           n60677, ZN => n13343);
   U3834 : OAI22_X1 port map( A1 => n60683, A2 => n61184, B1 => n3952, B2 => 
                           n60677, ZN => n13344);
   U3835 : OAI22_X1 port map( A1 => n60683, A2 => n61198, B1 => n3951, B2 => 
                           n15144, ZN => n13345);
   U3836 : OAI22_X1 port map( A1 => n60683, A2 => n61212, B1 => n3950, B2 => 
                           n15144, ZN => n13346);
   U3837 : OAI22_X1 port map( A1 => n60684, A2 => n61226, B1 => n3949, B2 => 
                           n15144, ZN => n13347);
   U3838 : OAI22_X1 port map( A1 => n60684, A2 => n61249, B1 => n3948, B2 => 
                           n15144, ZN => n13348);
   U3839 : OAI22_X1 port map( A1 => n60088, A2 => n61148, B1 => n1250, B2 => 
                           n60083, ZN => n11229);
   U3840 : OAI22_X1 port map( A1 => n60089, A2 => n61162, B1 => n1249, B2 => 
                           n60083, ZN => n11230);
   U3841 : OAI22_X1 port map( A1 => n60089, A2 => n61176, B1 => n1248, B2 => 
                           n60083, ZN => n11231);
   U3842 : OAI22_X1 port map( A1 => n60089, A2 => n61190, B1 => n1247, B2 => 
                           n60083, ZN => n11232);
   U3843 : OAI22_X1 port map( A1 => n60089, A2 => n61204, B1 => n1246, B2 => 
                           n15231, ZN => n11233);
   U3844 : OAI22_X1 port map( A1 => n60089, A2 => n61218, B1 => n1245, B2 => 
                           n15231, ZN => n11234);
   U3845 : OAI22_X1 port map( A1 => n60090, A2 => n61232, B1 => n1244, B2 => 
                           n15231, ZN => n11235);
   U3846 : OAI22_X1 port map( A1 => n60090, A2 => n61255, B1 => n1243, B2 => 
                           n15231, ZN => n11236);
   U3847 : OAI22_X1 port map( A1 => n60079, A2 => n61148, B1 => n1242, B2 => 
                           n60074, ZN => n11197);
   U3848 : OAI22_X1 port map( A1 => n60080, A2 => n61162, B1 => n1241, B2 => 
                           n60074, ZN => n11198);
   U3849 : OAI22_X1 port map( A1 => n60080, A2 => n61176, B1 => n1240, B2 => 
                           n60074, ZN => n11199);
   U3850 : OAI22_X1 port map( A1 => n60080, A2 => n61190, B1 => n1239, B2 => 
                           n60074, ZN => n11200);
   U3851 : OAI22_X1 port map( A1 => n60080, A2 => n61204, B1 => n1238, B2 => 
                           n15232, ZN => n11201);
   U3852 : OAI22_X1 port map( A1 => n60080, A2 => n61218, B1 => n1237, B2 => 
                           n15232, ZN => n11202);
   U3853 : OAI22_X1 port map( A1 => n60081, A2 => n61232, B1 => n1236, B2 => 
                           n15232, ZN => n11203);
   U3854 : OAI22_X1 port map( A1 => n60081, A2 => n61255, B1 => n1235, B2 => 
                           n15232, ZN => n11204);
   U3855 : OAI22_X1 port map( A1 => n60025, A2 => n61148, B1 => n1194, B2 => 
                           n60020, ZN => n11005);
   U3856 : OAI22_X1 port map( A1 => n60026, A2 => n61162, B1 => n1193, B2 => 
                           n60020, ZN => n11006);
   U3857 : OAI22_X1 port map( A1 => n60026, A2 => n61176, B1 => n1192, B2 => 
                           n60020, ZN => n11007);
   U3858 : OAI22_X1 port map( A1 => n60026, A2 => n61190, B1 => n1191, B2 => 
                           n60020, ZN => n11008);
   U3859 : OAI22_X1 port map( A1 => n60026, A2 => n61204, B1 => n1190, B2 => 
                           n15238, ZN => n11009);
   U3860 : OAI22_X1 port map( A1 => n60026, A2 => n61218, B1 => n1189, B2 => 
                           n15238, ZN => n11010);
   U3861 : OAI22_X1 port map( A1 => n60027, A2 => n61232, B1 => n1188, B2 => 
                           n15238, ZN => n11011);
   U3862 : OAI22_X1 port map( A1 => n60027, A2 => n61255, B1 => n1187, B2 => 
                           n15238, ZN => n11012);
   U3863 : OAI22_X1 port map( A1 => n60016, A2 => n61148, B1 => n1186, B2 => 
                           n60011, ZN => n10973);
   U3864 : OAI22_X1 port map( A1 => n60017, A2 => n61162, B1 => n1185, B2 => 
                           n60011, ZN => n10974);
   U3865 : OAI22_X1 port map( A1 => n60017, A2 => n61176, B1 => n1184, B2 => 
                           n60011, ZN => n10975);
   U3866 : OAI22_X1 port map( A1 => n60017, A2 => n61190, B1 => n1183, B2 => 
                           n60011, ZN => n10976);
   U3867 : OAI22_X1 port map( A1 => n60017, A2 => n61204, B1 => n1182, B2 => 
                           n15239, ZN => n10977);
   U3868 : OAI22_X1 port map( A1 => n60017, A2 => n61218, B1 => n1181, B2 => 
                           n15239, ZN => n10978);
   U3869 : OAI22_X1 port map( A1 => n60018, A2 => n61232, B1 => n1180, B2 => 
                           n15239, ZN => n10979);
   U3870 : OAI22_X1 port map( A1 => n60018, A2 => n61255, B1 => n1179, B2 => 
                           n15239, ZN => n10980);
   U3871 : OAI22_X1 port map( A1 => n60007, A2 => n61148, B1 => n1178, B2 => 
                           n60002, ZN => n10941);
   U3872 : OAI22_X1 port map( A1 => n60008, A2 => n61162, B1 => n1177, B2 => 
                           n60002, ZN => n10942);
   U3873 : OAI22_X1 port map( A1 => n60008, A2 => n61176, B1 => n1176, B2 => 
                           n60002, ZN => n10943);
   U3874 : OAI22_X1 port map( A1 => n60008, A2 => n61190, B1 => n1175, B2 => 
                           n60002, ZN => n10944);
   U3875 : OAI22_X1 port map( A1 => n60008, A2 => n61204, B1 => n1174, B2 => 
                           n15240, ZN => n10945);
   U3876 : OAI22_X1 port map( A1 => n60008, A2 => n61218, B1 => n1173, B2 => 
                           n15240, ZN => n10946);
   U3877 : OAI22_X1 port map( A1 => n60009, A2 => n61232, B1 => n1172, B2 => 
                           n15240, ZN => n10947);
   U3878 : OAI22_X1 port map( A1 => n60009, A2 => n61255, B1 => n1171, B2 => 
                           n15240, ZN => n10948);
   U3879 : OAI22_X1 port map( A1 => n59998, A2 => n61148, B1 => n1170, B2 => 
                           n59993, ZN => n10909);
   U3880 : OAI22_X1 port map( A1 => n59999, A2 => n61162, B1 => n1169, B2 => 
                           n59993, ZN => n10910);
   U3881 : OAI22_X1 port map( A1 => n59999, A2 => n61176, B1 => n1168, B2 => 
                           n59993, ZN => n10911);
   U3882 : OAI22_X1 port map( A1 => n59999, A2 => n61190, B1 => n1167, B2 => 
                           n59993, ZN => n10912);
   U3883 : OAI22_X1 port map( A1 => n59999, A2 => n61204, B1 => n1166, B2 => 
                           n15241, ZN => n10913);
   U3884 : OAI22_X1 port map( A1 => n59999, A2 => n61218, B1 => n1165, B2 => 
                           n15241, ZN => n10914);
   U3885 : OAI22_X1 port map( A1 => n60000, A2 => n61232, B1 => n1164, B2 => 
                           n15241, ZN => n10915);
   U3886 : OAI22_X1 port map( A1 => n60000, A2 => n61255, B1 => n1163, B2 => 
                           n15241, ZN => n10916);
   U3887 : OAI22_X1 port map( A1 => n59989, A2 => n61149, B1 => n1162, B2 => 
                           n59984, ZN => n10877);
   U3888 : OAI22_X1 port map( A1 => n59990, A2 => n61163, B1 => n1161, B2 => 
                           n59984, ZN => n10878);
   U3889 : OAI22_X1 port map( A1 => n59990, A2 => n61177, B1 => n1160, B2 => 
                           n59984, ZN => n10879);
   U3890 : OAI22_X1 port map( A1 => n59990, A2 => n61191, B1 => n1159, B2 => 
                           n59984, ZN => n10880);
   U3891 : OAI22_X1 port map( A1 => n59990, A2 => n61205, B1 => n1158, B2 => 
                           n15242, ZN => n10881);
   U3892 : OAI22_X1 port map( A1 => n59990, A2 => n61219, B1 => n1157, B2 => 
                           n15242, ZN => n10882);
   U3893 : OAI22_X1 port map( A1 => n59991, A2 => n61233, B1 => n1156, B2 => 
                           n15242, ZN => n10883);
   U3894 : OAI22_X1 port map( A1 => n59991, A2 => n61256, B1 => n1155, B2 => 
                           n15242, ZN => n10884);
   U3895 : OAI22_X1 port map( A1 => n59980, A2 => n61149, B1 => n1154, B2 => 
                           n59975, ZN => n10845);
   U3896 : OAI22_X1 port map( A1 => n59981, A2 => n61163, B1 => n1153, B2 => 
                           n59975, ZN => n10846);
   U3897 : OAI22_X1 port map( A1 => n59981, A2 => n61177, B1 => n1152, B2 => 
                           n59975, ZN => n10847);
   U3898 : OAI22_X1 port map( A1 => n59981, A2 => n61191, B1 => n1151, B2 => 
                           n59975, ZN => n10848);
   U3899 : OAI22_X1 port map( A1 => n59981, A2 => n61205, B1 => n1150, B2 => 
                           n15243, ZN => n10849);
   U3900 : OAI22_X1 port map( A1 => n59981, A2 => n61219, B1 => n1149, B2 => 
                           n15243, ZN => n10850);
   U3901 : OAI22_X1 port map( A1 => n59982, A2 => n61233, B1 => n1148, B2 => 
                           n15243, ZN => n10851);
   U3902 : OAI22_X1 port map( A1 => n59982, A2 => n61256, B1 => n1147, B2 => 
                           n15243, ZN => n10852);
   U3903 : OAI22_X1 port map( A1 => n59953, A2 => n61149, B1 => n1130, B2 => 
                           n59948, ZN => n10749);
   U3904 : OAI22_X1 port map( A1 => n59954, A2 => n61163, B1 => n1129, B2 => 
                           n59948, ZN => n10750);
   U3905 : OAI22_X1 port map( A1 => n59954, A2 => n61177, B1 => n1128, B2 => 
                           n59948, ZN => n10751);
   U3906 : OAI22_X1 port map( A1 => n59954, A2 => n61191, B1 => n1127, B2 => 
                           n59948, ZN => n10752);
   U3907 : OAI22_X1 port map( A1 => n59954, A2 => n61205, B1 => n1126, B2 => 
                           n15246, ZN => n10753);
   U3908 : OAI22_X1 port map( A1 => n59954, A2 => n61219, B1 => n1125, B2 => 
                           n15246, ZN => n10754);
   U3909 : OAI22_X1 port map( A1 => n59955, A2 => n61233, B1 => n1124, B2 => 
                           n15246, ZN => n10755);
   U3910 : OAI22_X1 port map( A1 => n59955, A2 => n61256, B1 => n1123, B2 => 
                           n15246, ZN => n10756);
   U3911 : OAI22_X1 port map( A1 => n59944, A2 => n61149, B1 => n1122, B2 => 
                           n59939, ZN => n10717);
   U3912 : OAI22_X1 port map( A1 => n59945, A2 => n61163, B1 => n1121, B2 => 
                           n59939, ZN => n10718);
   U3913 : OAI22_X1 port map( A1 => n59945, A2 => n61177, B1 => n1120, B2 => 
                           n59939, ZN => n10719);
   U3914 : OAI22_X1 port map( A1 => n59945, A2 => n61191, B1 => n1119, B2 => 
                           n59939, ZN => n10720);
   U3915 : OAI22_X1 port map( A1 => n59945, A2 => n61205, B1 => n1118, B2 => 
                           n15248, ZN => n10721);
   U3916 : OAI22_X1 port map( A1 => n59945, A2 => n61219, B1 => n1117, B2 => 
                           n15248, ZN => n10722);
   U3917 : OAI22_X1 port map( A1 => n59946, A2 => n61233, B1 => n1116, B2 => 
                           n15248, ZN => n10723);
   U3918 : OAI22_X1 port map( A1 => n59946, A2 => n61256, B1 => n1115, B2 => 
                           n15248, ZN => n10724);
   U3919 : OAI22_X1 port map( A1 => n59935, A2 => n61149, B1 => n1114, B2 => 
                           n59930, ZN => n10685);
   U3920 : OAI22_X1 port map( A1 => n59917, A2 => n61149, B1 => n1113, B2 => 
                           n59912, ZN => n10621);
   U3921 : OAI22_X1 port map( A1 => n59918, A2 => n61163, B1 => n1112, B2 => 
                           n59912, ZN => n10622);
   U3922 : OAI22_X1 port map( A1 => n59918, A2 => n61177, B1 => n1111, B2 => 
                           n59912, ZN => n10623);
   U3923 : OAI22_X1 port map( A1 => n59918, A2 => n61191, B1 => n1110, B2 => 
                           n59912, ZN => n10624);
   U3924 : OAI22_X1 port map( A1 => n59918, A2 => n61205, B1 => n1109, B2 => 
                           n15251, ZN => n10625);
   U3925 : OAI22_X1 port map( A1 => n59918, A2 => n61219, B1 => n1108, B2 => 
                           n15251, ZN => n10626);
   U3926 : OAI22_X1 port map( A1 => n59919, A2 => n61233, B1 => n1107, B2 => 
                           n15251, ZN => n10627);
   U3927 : OAI22_X1 port map( A1 => n59919, A2 => n61256, B1 => n1106, B2 => 
                           n15251, ZN => n10628);
   U3928 : OAI22_X1 port map( A1 => n59899, A2 => n61149, B1 => n1097, B2 => 
                           n59894, ZN => n10557);
   U3929 : OAI22_X1 port map( A1 => n59900, A2 => n61163, B1 => n1096, B2 => 
                           n59894, ZN => n10558);
   U3930 : OAI22_X1 port map( A1 => n59900, A2 => n61177, B1 => n1095, B2 => 
                           n59894, ZN => n10559);
   U3931 : OAI22_X1 port map( A1 => n59900, A2 => n61191, B1 => n1094, B2 => 
                           n59894, ZN => n10560);
   U3932 : OAI22_X1 port map( A1 => n59900, A2 => n61205, B1 => n1093, B2 => 
                           n15253, ZN => n10561);
   U3933 : OAI22_X1 port map( A1 => n59900, A2 => n61219, B1 => n1092, B2 => 
                           n15253, ZN => n10562);
   U3934 : OAI22_X1 port map( A1 => n59901, A2 => n61233, B1 => n1091, B2 => 
                           n15253, ZN => n10563);
   U3935 : OAI22_X1 port map( A1 => n59901, A2 => n61256, B1 => n1090, B2 => 
                           n15253, ZN => n10564);
   U3936 : OAI22_X1 port map( A1 => n59890, A2 => n61149, B1 => n1089, B2 => 
                           n59885, ZN => n10525);
   U3937 : OAI22_X1 port map( A1 => n59891, A2 => n61163, B1 => n1088, B2 => 
                           n59885, ZN => n10526);
   U3938 : OAI22_X1 port map( A1 => n59891, A2 => n61177, B1 => n1087, B2 => 
                           n59885, ZN => n10527);
   U3939 : OAI22_X1 port map( A1 => n59891, A2 => n61191, B1 => n1086, B2 => 
                           n59885, ZN => n10528);
   U3940 : OAI22_X1 port map( A1 => n59891, A2 => n61205, B1 => n1085, B2 => 
                           n15254, ZN => n10529);
   U3941 : OAI22_X1 port map( A1 => n59891, A2 => n61219, B1 => n1084, B2 => 
                           n15254, ZN => n10530);
   U3942 : OAI22_X1 port map( A1 => n59892, A2 => n61233, B1 => n1083, B2 => 
                           n15254, ZN => n10531);
   U3943 : OAI22_X1 port map( A1 => n59892, A2 => n61256, B1 => n1082, B2 => 
                           n15254, ZN => n10532);
   U3944 : OAI22_X1 port map( A1 => n59881, A2 => n61150, B1 => n1081, B2 => 
                           n59876, ZN => n10493);
   U3945 : OAI22_X1 port map( A1 => n59882, A2 => n61164, B1 => n1080, B2 => 
                           n59876, ZN => n10494);
   U3946 : OAI22_X1 port map( A1 => n59882, A2 => n61178, B1 => n1079, B2 => 
                           n59876, ZN => n10495);
   U3947 : OAI22_X1 port map( A1 => n59882, A2 => n61192, B1 => n1078, B2 => 
                           n59876, ZN => n10496);
   U3948 : OAI22_X1 port map( A1 => n59882, A2 => n61206, B1 => n1077, B2 => 
                           n15255, ZN => n10497);
   U3949 : OAI22_X1 port map( A1 => n59882, A2 => n61220, B1 => n1076, B2 => 
                           n15255, ZN => n10498);
   U3950 : OAI22_X1 port map( A1 => n59883, A2 => n61234, B1 => n1075, B2 => 
                           n15255, ZN => n10499);
   U3951 : OAI22_X1 port map( A1 => n59883, A2 => n61257, B1 => n1074, B2 => 
                           n15255, ZN => n10500);
   U3952 : OAI22_X1 port map( A1 => n59872, A2 => n61150, B1 => n1073, B2 => 
                           n59867, ZN => n10461);
   U3953 : OAI22_X1 port map( A1 => n59873, A2 => n61164, B1 => n1072, B2 => 
                           n59867, ZN => n10462);
   U3954 : OAI22_X1 port map( A1 => n59873, A2 => n61178, B1 => n1071, B2 => 
                           n59867, ZN => n10463);
   U3955 : OAI22_X1 port map( A1 => n59873, A2 => n61192, B1 => n1070, B2 => 
                           n59867, ZN => n10464);
   U3956 : OAI22_X1 port map( A1 => n59854, A2 => n61150, B1 => n1069, B2 => 
                           n59849, ZN => n10397);
   U3957 : OAI22_X1 port map( A1 => n59855, A2 => n61164, B1 => n1068, B2 => 
                           n59849, ZN => n10398);
   U3958 : OAI22_X1 port map( A1 => n59855, A2 => n61178, B1 => n1067, B2 => 
                           n59849, ZN => n10399);
   U3959 : OAI22_X1 port map( A1 => n59855, A2 => n61192, B1 => n1066, B2 => 
                           n59849, ZN => n10400);
   U3960 : OAI22_X1 port map( A1 => n59855, A2 => n61206, B1 => n1065, B2 => 
                           n15262, ZN => n10401);
   U3961 : OAI22_X1 port map( A1 => n59855, A2 => n61220, B1 => n1064, B2 => 
                           n15262, ZN => n10402);
   U3962 : OAI22_X1 port map( A1 => n59856, A2 => n61234, B1 => n1063, B2 => 
                           n15262, ZN => n10403);
   U3963 : OAI22_X1 port map( A1 => n59856, A2 => n61257, B1 => n1062, B2 => 
                           n15262, ZN => n10404);
   U3964 : OAI22_X1 port map( A1 => n59845, A2 => n61150, B1 => n1061, B2 => 
                           n59840, ZN => n10365);
   U3965 : OAI22_X1 port map( A1 => n59846, A2 => n61164, B1 => n1060, B2 => 
                           n59840, ZN => n10366);
   U3966 : OAI22_X1 port map( A1 => n59846, A2 => n61178, B1 => n1059, B2 => 
                           n59840, ZN => n10367);
   U3967 : OAI22_X1 port map( A1 => n59846, A2 => n61192, B1 => n1058, B2 => 
                           n59840, ZN => n10368);
   U3968 : OAI22_X1 port map( A1 => n59846, A2 => n61206, B1 => n1057, B2 => 
                           n15264, ZN => n10369);
   U3969 : OAI22_X1 port map( A1 => n59846, A2 => n61220, B1 => n1056, B2 => 
                           n15264, ZN => n10370);
   U3970 : OAI22_X1 port map( A1 => n59847, A2 => n61234, B1 => n1055, B2 => 
                           n15264, ZN => n10371);
   U3971 : OAI22_X1 port map( A1 => n59847, A2 => n61257, B1 => n1054, B2 => 
                           n15264, ZN => n10372);
   U3972 : OAI22_X1 port map( A1 => n60673, A2 => n61142, B1 => n1045, B2 => 
                           n60668, ZN => n13309);
   U3973 : OAI22_X1 port map( A1 => n60674, A2 => n61156, B1 => n1044, B2 => 
                           n60668, ZN => n13310);
   U3974 : OAI22_X1 port map( A1 => n60674, A2 => n61170, B1 => n1043, B2 => 
                           n60668, ZN => n13311);
   U3975 : OAI22_X1 port map( A1 => n60674, A2 => n61184, B1 => n1042, B2 => 
                           n60668, ZN => n13312);
   U3976 : OAI22_X1 port map( A1 => n60674, A2 => n61198, B1 => n1041, B2 => 
                           n15146, ZN => n13313);
   U3977 : OAI22_X1 port map( A1 => n60674, A2 => n61212, B1 => n1040, B2 => 
                           n15146, ZN => n13314);
   U3978 : OAI22_X1 port map( A1 => n60675, A2 => n61226, B1 => n1039, B2 => 
                           n15146, ZN => n13315);
   U3979 : OAI22_X1 port map( A1 => n60675, A2 => n61249, B1 => n1038, B2 => 
                           n15146, ZN => n13316);
   U3980 : OAI22_X1 port map( A1 => n60637, A2 => n61143, B1 => n1029, B2 => 
                           n60632, ZN => n13181);
   U3981 : OAI22_X1 port map( A1 => n60638, A2 => n61157, B1 => n1028, B2 => 
                           n60632, ZN => n13182);
   U3982 : OAI22_X1 port map( A1 => n60638, A2 => n61171, B1 => n1027, B2 => 
                           n60632, ZN => n13183);
   U3983 : OAI22_X1 port map( A1 => n60638, A2 => n61185, B1 => n1026, B2 => 
                           n60632, ZN => n13184);
   U3984 : OAI22_X1 port map( A1 => n60638, A2 => n61199, B1 => n1025, B2 => 
                           n15151, ZN => n13185);
   U3985 : OAI22_X1 port map( A1 => n60638, A2 => n61213, B1 => n1024, B2 => 
                           n15151, ZN => n13186);
   U3986 : OAI22_X1 port map( A1 => n60639, A2 => n61227, B1 => n1023, B2 => 
                           n15151, ZN => n13187);
   U3987 : OAI22_X1 port map( A1 => n60639, A2 => n61250, B1 => n1022, B2 => 
                           n15151, ZN => n13188);
   U3988 : OAI22_X1 port map( A1 => n60628, A2 => n61143, B1 => n1021, B2 => 
                           n60623, ZN => n13149);
   U3989 : OAI22_X1 port map( A1 => n60629, A2 => n61157, B1 => n1020, B2 => 
                           n60623, ZN => n13150);
   U3990 : OAI22_X1 port map( A1 => n60629, A2 => n61171, B1 => n1019, B2 => 
                           n60623, ZN => n13151);
   U3991 : OAI22_X1 port map( A1 => n60629, A2 => n61185, B1 => n1018, B2 => 
                           n60623, ZN => n13152);
   U3992 : OAI22_X1 port map( A1 => n60629, A2 => n61199, B1 => n1017, B2 => 
                           n15152, ZN => n13153);
   U3993 : OAI22_X1 port map( A1 => n60629, A2 => n61213, B1 => n1016, B2 => 
                           n15152, ZN => n13154);
   U3994 : OAI22_X1 port map( A1 => n60630, A2 => n61227, B1 => n1015, B2 => 
                           n15152, ZN => n13155);
   U3995 : OAI22_X1 port map( A1 => n60630, A2 => n61250, B1 => n1014, B2 => 
                           n15152, ZN => n13156);
   U3996 : OAI22_X1 port map( A1 => n60601, A2 => n61143, B1 => n1013, B2 => 
                           n60596, ZN => n13053);
   U3997 : OAI22_X1 port map( A1 => n60602, A2 => n61157, B1 => n1012, B2 => 
                           n60596, ZN => n13054);
   U3998 : OAI22_X1 port map( A1 => n60602, A2 => n61171, B1 => n1011, B2 => 
                           n60596, ZN => n13055);
   U3999 : OAI22_X1 port map( A1 => n60602, A2 => n61185, B1 => n1010, B2 => 
                           n60596, ZN => n13056);
   U4000 : OAI22_X1 port map( A1 => n60602, A2 => n61199, B1 => n1009, B2 => 
                           n15155, ZN => n13057);
   U4001 : OAI22_X1 port map( A1 => n60602, A2 => n61213, B1 => n1008, B2 => 
                           n15155, ZN => n13058);
   U4002 : OAI22_X1 port map( A1 => n60603, A2 => n61227, B1 => n1007, B2 => 
                           n15155, ZN => n13059);
   U4003 : OAI22_X1 port map( A1 => n60603, A2 => n61250, B1 => n1006, B2 => 
                           n15155, ZN => n13060);
   U4004 : OAI22_X1 port map( A1 => n60592, A2 => n61143, B1 => n1005, B2 => 
                           n60587, ZN => n13021);
   U4005 : OAI22_X1 port map( A1 => n60593, A2 => n61157, B1 => n1004, B2 => 
                           n60587, ZN => n13022);
   U4006 : OAI22_X1 port map( A1 => n60593, A2 => n61171, B1 => n1003, B2 => 
                           n60587, ZN => n13023);
   U4007 : OAI22_X1 port map( A1 => n60593, A2 => n61185, B1 => n1002, B2 => 
                           n60587, ZN => n13024);
   U4008 : OAI22_X1 port map( A1 => n60593, A2 => n61199, B1 => n1001, B2 => 
                           n15156, ZN => n13025);
   U4009 : OAI22_X1 port map( A1 => n60593, A2 => n61213, B1 => n1000, B2 => 
                           n15156, ZN => n13026);
   U4010 : OAI22_X1 port map( A1 => n60594, A2 => n61227, B1 => n995, B2 => 
                           n15156, ZN => n13027);
   U4011 : OAI22_X1 port map( A1 => n60594, A2 => n61250, B1 => n994, B2 => 
                           n15156, ZN => n13028);
   U4012 : OAI22_X1 port map( A1 => n60565, A2 => n61143, B1 => n993, B2 => 
                           n60560, ZN => n12925);
   U4013 : OAI22_X1 port map( A1 => n60566, A2 => n61157, B1 => n992, B2 => 
                           n60560, ZN => n12926);
   U4014 : OAI22_X1 port map( A1 => n60566, A2 => n61171, B1 => n991, B2 => 
                           n60560, ZN => n12927);
   U4015 : OAI22_X1 port map( A1 => n60566, A2 => n61185, B1 => n990, B2 => 
                           n60560, ZN => n12928);
   U4016 : OAI22_X1 port map( A1 => n60566, A2 => n61199, B1 => n989, B2 => 
                           n15159, ZN => n12929);
   U4017 : OAI22_X1 port map( A1 => n60566, A2 => n61213, B1 => n988, B2 => 
                           n15159, ZN => n12930);
   U4018 : OAI22_X1 port map( A1 => n60567, A2 => n61227, B1 => n987, B2 => 
                           n15159, ZN => n12931);
   U4019 : OAI22_X1 port map( A1 => n60567, A2 => n61250, B1 => n986, B2 => 
                           n15159, ZN => n12932);
   U4020 : OAI22_X1 port map( A1 => n60557, A2 => n61213, B1 => n985, B2 => 
                           n15160, ZN => n12898);
   U4021 : OAI22_X1 port map( A1 => n60558, A2 => n61227, B1 => n984, B2 => 
                           n15160, ZN => n12899);
   U4022 : OAI22_X1 port map( A1 => n60558, A2 => n61250, B1 => n983, B2 => 
                           n15160, ZN => n12900);
   U4023 : OAI22_X1 port map( A1 => n60529, A2 => n61144, B1 => n982, B2 => 
                           n60524, ZN => n12797);
   U4024 : OAI22_X1 port map( A1 => n60530, A2 => n61158, B1 => n981, B2 => 
                           n60524, ZN => n12798);
   U4025 : OAI22_X1 port map( A1 => n60530, A2 => n61172, B1 => n980, B2 => 
                           n60524, ZN => n12799);
   U4026 : OAI22_X1 port map( A1 => n60530, A2 => n61186, B1 => n979, B2 => 
                           n60524, ZN => n12800);
   U4027 : OAI22_X1 port map( A1 => n60530, A2 => n61200, B1 => n978, B2 => 
                           n15163, ZN => n12801);
   U4028 : OAI22_X1 port map( A1 => n60530, A2 => n61214, B1 => n977, B2 => 
                           n15163, ZN => n12802);
   U4029 : OAI22_X1 port map( A1 => n60531, A2 => n61228, B1 => n976, B2 => 
                           n15163, ZN => n12803);
   U4030 : OAI22_X1 port map( A1 => n60531, A2 => n61251, B1 => n975, B2 => 
                           n15163, ZN => n12804);
   U4031 : OAI22_X1 port map( A1 => n60520, A2 => n61144, B1 => n974, B2 => 
                           n60515, ZN => n12765);
   U4032 : OAI22_X1 port map( A1 => n60521, A2 => n61158, B1 => n973, B2 => 
                           n60515, ZN => n12766);
   U4033 : OAI22_X1 port map( A1 => n60521, A2 => n61172, B1 => n972, B2 => 
                           n60515, ZN => n12767);
   U4034 : OAI22_X1 port map( A1 => n60521, A2 => n61186, B1 => n815, B2 => 
                           n60515, ZN => n12768);
   U4035 : OAI22_X1 port map( A1 => n60521, A2 => n61200, B1 => n814, B2 => 
                           n15165, ZN => n12769);
   U4036 : OAI22_X1 port map( A1 => n60521, A2 => n61214, B1 => n813, B2 => 
                           n15165, ZN => n12770);
   U4037 : OAI22_X1 port map( A1 => n60522, A2 => n61228, B1 => n812, B2 => 
                           n15165, ZN => n12771);
   U4038 : OAI22_X1 port map( A1 => n60522, A2 => n61251, B1 => n811, B2 => 
                           n15165, ZN => n12772);
   U4039 : OAI22_X1 port map( A1 => n60502, A2 => n61144, B1 => n802, B2 => 
                           n60497, ZN => n12701);
   U4040 : OAI22_X1 port map( A1 => n60503, A2 => n61158, B1 => n801, B2 => 
                           n60497, ZN => n12702);
   U4041 : OAI22_X1 port map( A1 => n60503, A2 => n61172, B1 => n800, B2 => 
                           n60497, ZN => n12703);
   U4042 : OAI22_X1 port map( A1 => n60503, A2 => n61186, B1 => n799, B2 => 
                           n60497, ZN => n12704);
   U4043 : OAI22_X1 port map( A1 => n60503, A2 => n61200, B1 => n798, B2 => 
                           n15167, ZN => n12705);
   U4044 : OAI22_X1 port map( A1 => n60503, A2 => n61214, B1 => n797, B2 => 
                           n15167, ZN => n12706);
   U4045 : OAI22_X1 port map( A1 => n60504, A2 => n61228, B1 => n796, B2 => 
                           n15167, ZN => n12707);
   U4046 : OAI22_X1 port map( A1 => n60504, A2 => n61251, B1 => n795, B2 => 
                           n15167, ZN => n12708);
   U4047 : OAI22_X1 port map( A1 => n60493, A2 => n61144, B1 => n794, B2 => 
                           n60488, ZN => n12669);
   U4048 : OAI22_X1 port map( A1 => n60494, A2 => n61158, B1 => n793, B2 => 
                           n60488, ZN => n12670);
   U4049 : OAI22_X1 port map( A1 => n60494, A2 => n61172, B1 => n792, B2 => 
                           n60488, ZN => n12671);
   U4050 : OAI22_X1 port map( A1 => n60494, A2 => n61186, B1 => n791, B2 => 
                           n60488, ZN => n12672);
   U4051 : OAI22_X1 port map( A1 => n60494, A2 => n61200, B1 => n790, B2 => 
                           n15168, ZN => n12673);
   U4052 : OAI22_X1 port map( A1 => n60494, A2 => n61214, B1 => n789, B2 => 
                           n15168, ZN => n12674);
   U4053 : OAI22_X1 port map( A1 => n60495, A2 => n61228, B1 => n788, B2 => 
                           n15168, ZN => n12675);
   U4054 : OAI22_X1 port map( A1 => n60495, A2 => n61251, B1 => n787, B2 => 
                           n15168, ZN => n12676);
   U4055 : OAI22_X1 port map( A1 => n60448, A2 => n61144, B1 => n770, B2 => 
                           n60443, ZN => n12509);
   U4056 : OAI22_X1 port map( A1 => n60449, A2 => n61158, B1 => n769, B2 => 
                           n60443, ZN => n12510);
   U4057 : OAI22_X1 port map( A1 => n60449, A2 => n61172, B1 => n768, B2 => 
                           n60443, ZN => n12511);
   U4058 : OAI22_X1 port map( A1 => n60449, A2 => n61186, B1 => n767, B2 => 
                           n60443, ZN => n12512);
   U4059 : OAI22_X1 port map( A1 => n60449, A2 => n61200, B1 => n766, B2 => 
                           n15180, ZN => n12513);
   U4060 : OAI22_X1 port map( A1 => n60449, A2 => n61214, B1 => n765, B2 => 
                           n15180, ZN => n12514);
   U4061 : OAI22_X1 port map( A1 => n60450, A2 => n61228, B1 => n764, B2 => 
                           n15180, ZN => n12515);
   U4062 : OAI22_X1 port map( A1 => n60450, A2 => n61251, B1 => n763, B2 => 
                           n15180, ZN => n12516);
   U4063 : OAI22_X1 port map( A1 => n60439, A2 => n61144, B1 => n762, B2 => 
                           n60434, ZN => n12477);
   U4064 : OAI22_X1 port map( A1 => n60440, A2 => n61158, B1 => n761, B2 => 
                           n60434, ZN => n12478);
   U4065 : OAI22_X1 port map( A1 => n60440, A2 => n61172, B1 => n760, B2 => 
                           n60434, ZN => n12479);
   U4066 : OAI22_X1 port map( A1 => n60440, A2 => n61186, B1 => n567, B2 => 
                           n60434, ZN => n12480);
   U4067 : OAI22_X1 port map( A1 => n60440, A2 => n61200, B1 => n566, B2 => 
                           n15181, ZN => n12481);
   U4068 : OAI22_X1 port map( A1 => n60440, A2 => n61214, B1 => n565, B2 => 
                           n15181, ZN => n12482);
   U4069 : OAI22_X1 port map( A1 => n60441, A2 => n61228, B1 => n564, B2 => 
                           n15181, ZN => n12483);
   U4070 : OAI22_X1 port map( A1 => n60441, A2 => n61251, B1 => n563, B2 => 
                           n15181, ZN => n12484);
   U4071 : OAI22_X1 port map( A1 => n60430, A2 => n61144, B1 => n562, B2 => 
                           n60425, ZN => n12445);
   U4072 : OAI22_X1 port map( A1 => n60431, A2 => n61158, B1 => n561, B2 => 
                           n60425, ZN => n12446);
   U4073 : OAI22_X1 port map( A1 => n60431, A2 => n61172, B1 => n560, B2 => 
                           n60425, ZN => n12447);
   U4074 : OAI22_X1 port map( A1 => n60431, A2 => n61186, B1 => n499, B2 => 
                           n60425, ZN => n12448);
   U4075 : OAI22_X1 port map( A1 => n60431, A2 => n61200, B1 => n498, B2 => 
                           n15182, ZN => n12449);
   U4076 : OAI22_X1 port map( A1 => n60431, A2 => n61214, B1 => n497, B2 => 
                           n15182, ZN => n12450);
   U4077 : OAI22_X1 port map( A1 => n60432, A2 => n61228, B1 => n496, B2 => 
                           n15182, ZN => n12451);
   U4078 : OAI22_X1 port map( A1 => n60432, A2 => n61251, B1 => n495, B2 => 
                           n15182, ZN => n12452);
   U4079 : OAI22_X1 port map( A1 => n60421, A2 => n61145, B1 => n494, B2 => 
                           n60416, ZN => n12413);
   U4080 : OAI22_X1 port map( A1 => n60422, A2 => n61159, B1 => n493, B2 => 
                           n60416, ZN => n12414);
   U4081 : OAI22_X1 port map( A1 => n60422, A2 => n61173, B1 => n492, B2 => 
                           n60416, ZN => n12415);
   U4082 : OAI22_X1 port map( A1 => n60422, A2 => n61187, B1 => n491, B2 => 
                           n60416, ZN => n12416);
   U4083 : OAI22_X1 port map( A1 => n60422, A2 => n61201, B1 => n490, B2 => 
                           n15183, ZN => n12417);
   U4084 : OAI22_X1 port map( A1 => n60422, A2 => n61215, B1 => n489, B2 => 
                           n15183, ZN => n12418);
   U4085 : OAI22_X1 port map( A1 => n60423, A2 => n61229, B1 => n488, B2 => 
                           n15183, ZN => n12419);
   U4086 : OAI22_X1 port map( A1 => n60423, A2 => n61252, B1 => n487, B2 => 
                           n15183, ZN => n12420);
   U4087 : OAI22_X1 port map( A1 => n61241, A2 => n61140, B1 => n486, B2 => 
                           n61236, ZN => n14333);
   U4088 : OAI22_X1 port map( A1 => n61242, A2 => n61154, B1 => n485, B2 => 
                           n61236, ZN => n14334);
   U4089 : OAI22_X1 port map( A1 => n61242, A2 => n61168, B1 => n484, B2 => 
                           n61236, ZN => n14335);
   U4090 : OAI22_X1 port map( A1 => n61242, A2 => n61182, B1 => n483, B2 => 
                           n61236, ZN => n14336);
   U4091 : OAI22_X1 port map( A1 => n61242, A2 => n61196, B1 => n482, B2 => 
                           n15073, ZN => n14337);
   U4092 : OAI22_X1 port map( A1 => n61242, A2 => n61210, B1 => n481, B2 => 
                           n15073, ZN => n14338);
   U4093 : OAI22_X1 port map( A1 => n61243, A2 => n61224, B1 => n480, B2 => 
                           n15073, ZN => n14339);
   U4094 : OAI22_X1 port map( A1 => n61243, A2 => n61247, B1 => n479, B2 => 
                           n15073, ZN => n14340);
   U4095 : OAI22_X1 port map( A1 => n60952, A2 => n61140, B1 => n478, B2 => 
                           n60947, ZN => n14301);
   U4096 : OAI22_X1 port map( A1 => n60953, A2 => n61154, B1 => n477, B2 => 
                           n60947, ZN => n14302);
   U4097 : OAI22_X1 port map( A1 => n60953, A2 => n61168, B1 => n476, B2 => 
                           n60947, ZN => n14303);
   U4098 : OAI22_X1 port map( A1 => n60953, A2 => n61182, B1 => n473, B2 => 
                           n60947, ZN => n14304);
   U4099 : OAI22_X1 port map( A1 => n60953, A2 => n61196, B1 => n472, B2 => 
                           n15096, ZN => n14305);
   U4100 : OAI22_X1 port map( A1 => n60953, A2 => n61210, B1 => n471, B2 => 
                           n15096, ZN => n14306);
   U4101 : OAI22_X1 port map( A1 => n60954, A2 => n61224, B1 => n470, B2 => 
                           n15096, ZN => n14307);
   U4102 : OAI22_X1 port map( A1 => n60954, A2 => n61247, B1 => n469, B2 => 
                           n15096, ZN => n14308);
   U4103 : OAI22_X1 port map( A1 => n60907, A2 => n61140, B1 => n468, B2 => 
                           n60902, ZN => n14141);
   U4104 : OAI22_X1 port map( A1 => n60908, A2 => n61154, B1 => n467, B2 => 
                           n60902, ZN => n14142);
   U4105 : OAI22_X1 port map( A1 => n60908, A2 => n61168, B1 => n466, B2 => 
                           n60902, ZN => n14143);
   U4106 : OAI22_X1 port map( A1 => n60908, A2 => n61182, B1 => n465, B2 => 
                           n60902, ZN => n14144);
   U4107 : OAI22_X1 port map( A1 => n60908, A2 => n61196, B1 => n464, B2 => 
                           n15106, ZN => n14145);
   U4108 : OAI22_X1 port map( A1 => n60908, A2 => n61210, B1 => n463, B2 => 
                           n15106, ZN => n14146);
   U4109 : OAI22_X1 port map( A1 => n60909, A2 => n61224, B1 => n462, B2 => 
                           n15106, ZN => n14147);
   U4110 : OAI22_X1 port map( A1 => n60909, A2 => n61247, B1 => n461, B2 => 
                           n15106, ZN => n14148);
   U4111 : OAI22_X1 port map( A1 => n60385, A2 => n61145, B1 => n388, B2 => 
                           n60380, ZN => n12285);
   U4112 : OAI22_X1 port map( A1 => n60386, A2 => n61159, B1 => n371, B2 => 
                           n60380, ZN => n12286);
   U4113 : OAI22_X1 port map( A1 => n60386, A2 => n61173, B1 => n370, B2 => 
                           n60380, ZN => n12287);
   U4114 : OAI22_X1 port map( A1 => n60386, A2 => n61187, B1 => n369, B2 => 
                           n60380, ZN => n12288);
   U4115 : OAI22_X1 port map( A1 => n60386, A2 => n61201, B1 => n368, B2 => 
                           n15187, ZN => n12289);
   U4116 : OAI22_X1 port map( A1 => n60386, A2 => n61215, B1 => n367, B2 => 
                           n15187, ZN => n12290);
   U4117 : OAI22_X1 port map( A1 => n60387, A2 => n61229, B1 => n366, B2 => 
                           n15187, ZN => n12291);
   U4118 : OAI22_X1 port map( A1 => n60387, A2 => n61252, B1 => n365, B2 => 
                           n15187, ZN => n12292);
   U4119 : OAI22_X1 port map( A1 => n60313, A2 => n61146, B1 => n332, B2 => 
                           n60308, ZN => n12029);
   U4120 : OAI22_X1 port map( A1 => n60314, A2 => n61160, B1 => n331, B2 => 
                           n60308, ZN => n12030);
   U4121 : OAI22_X1 port map( A1 => n60314, A2 => n61174, B1 => n330, B2 => 
                           n60308, ZN => n12031);
   U4122 : OAI22_X1 port map( A1 => n60314, A2 => n61188, B1 => n329, B2 => 
                           n60308, ZN => n12032);
   U4123 : OAI22_X1 port map( A1 => n60314, A2 => n61202, B1 => n328, B2 => 
                           n15196, ZN => n12033);
   U4124 : OAI22_X1 port map( A1 => n60314, A2 => n61216, B1 => n327, B2 => 
                           n15196, ZN => n12034);
   U4125 : OAI22_X1 port map( A1 => n60315, A2 => n61230, B1 => n326, B2 => 
                           n15196, ZN => n12035);
   U4126 : OAI22_X1 port map( A1 => n60315, A2 => n61253, B1 => n325, B2 => 
                           n15196, ZN => n12036);
   U4127 : OAI22_X1 port map( A1 => n60304, A2 => n61146, B1 => n324, B2 => 
                           n60299, ZN => n11997);
   U4128 : OAI22_X1 port map( A1 => n60305, A2 => n61160, B1 => n323, B2 => 
                           n60299, ZN => n11998);
   U4129 : OAI22_X1 port map( A1 => n60305, A2 => n61174, B1 => n322, B2 => 
                           n60299, ZN => n11999);
   U4130 : OAI22_X1 port map( A1 => n60305, A2 => n61188, B1 => n321, B2 => 
                           n60299, ZN => n12000);
   U4131 : OAI22_X1 port map( A1 => n60305, A2 => n61202, B1 => n320, B2 => 
                           n15197, ZN => n12001);
   U4132 : OAI22_X1 port map( A1 => n60305, A2 => n61216, B1 => n319, B2 => 
                           n15197, ZN => n12002);
   U4133 : OAI22_X1 port map( A1 => n60306, A2 => n61230, B1 => n318, B2 => 
                           n15197, ZN => n12003);
   U4134 : OAI22_X1 port map( A1 => n60306, A2 => n61253, B1 => n317, B2 => 
                           n15197, ZN => n12004);
   U4135 : OAI22_X1 port map( A1 => n60259, A2 => n61146, B1 => n300, B2 => 
                           n60254, ZN => n11837);
   U4136 : OAI22_X1 port map( A1 => n60260, A2 => n61160, B1 => n299, B2 => 
                           n60254, ZN => n11838);
   U4137 : OAI22_X1 port map( A1 => n60260, A2 => n61174, B1 => n298, B2 => 
                           n60254, ZN => n11839);
   U4138 : OAI22_X1 port map( A1 => n60260, A2 => n61188, B1 => n297, B2 => 
                           n60254, ZN => n11840);
   U4139 : OAI22_X1 port map( A1 => n60260, A2 => n61202, B1 => n296, B2 => 
                           n15202, ZN => n11841);
   U4140 : OAI22_X1 port map( A1 => n60260, A2 => n61216, B1 => n295, B2 => 
                           n15202, ZN => n11842);
   U4141 : OAI22_X1 port map( A1 => n60261, A2 => n61230, B1 => n294, B2 => 
                           n15202, ZN => n11843);
   U4142 : OAI22_X1 port map( A1 => n60261, A2 => n61253, B1 => n293, B2 => 
                           n15202, ZN => n11844);
   U4143 : OAI22_X1 port map( A1 => n60241, A2 => n61146, B1 => n284, B2 => 
                           n60236, ZN => n11773);
   U4144 : OAI22_X1 port map( A1 => n60242, A2 => n61160, B1 => n283, B2 => 
                           n60236, ZN => n11774);
   U4145 : OAI22_X1 port map( A1 => n60242, A2 => n61174, B1 => n282, B2 => 
                           n60236, ZN => n11775);
   U4146 : OAI22_X1 port map( A1 => n60242, A2 => n61188, B1 => n281, B2 => 
                           n60236, ZN => n11776);
   U4147 : OAI22_X1 port map( A1 => n60242, A2 => n61202, B1 => n280, B2 => 
                           n15212, ZN => n11777);
   U4148 : OAI22_X1 port map( A1 => n60242, A2 => n61216, B1 => n279, B2 => 
                           n15212, ZN => n11778);
   U4149 : OAI22_X1 port map( A1 => n60243, A2 => n61230, B1 => n278, B2 => 
                           n15212, ZN => n11779);
   U4150 : OAI22_X1 port map( A1 => n60243, A2 => n61253, B1 => n277, B2 => 
                           n15212, ZN => n11780);
   U4151 : OAI22_X1 port map( A1 => n60232, A2 => n61146, B1 => n276, B2 => 
                           n60227, ZN => n11741);
   U4152 : OAI22_X1 port map( A1 => n60233, A2 => n61160, B1 => n275, B2 => 
                           n60227, ZN => n11742);
   U4153 : OAI22_X1 port map( A1 => n60233, A2 => n61174, B1 => n274, B2 => 
                           n60227, ZN => n11743);
   U4154 : OAI22_X1 port map( A1 => n60233, A2 => n61188, B1 => n273, B2 => 
                           n60227, ZN => n11744);
   U4155 : OAI22_X1 port map( A1 => n60233, A2 => n61202, B1 => n272, B2 => 
                           n15214, ZN => n11745);
   U4156 : OAI22_X1 port map( A1 => n60233, A2 => n61216, B1 => n271, B2 => 
                           n15214, ZN => n11746);
   U4157 : OAI22_X1 port map( A1 => n60234, A2 => n61230, B1 => n270, B2 => 
                           n15214, ZN => n11747);
   U4158 : OAI22_X1 port map( A1 => n60234, A2 => n61253, B1 => n269, B2 => 
                           n15214, ZN => n11748);
   U4159 : OAI22_X1 port map( A1 => n60205, A2 => n61147, B1 => n268, B2 => 
                           n60200, ZN => n11645);
   U4160 : OAI22_X1 port map( A1 => n60206, A2 => n61161, B1 => n267, B2 => 
                           n60200, ZN => n11646);
   U4161 : OAI22_X1 port map( A1 => n60206, A2 => n61175, B1 => n266, B2 => 
                           n60200, ZN => n11647);
   U4162 : OAI22_X1 port map( A1 => n60206, A2 => n61189, B1 => n265, B2 => 
                           n60200, ZN => n11648);
   U4163 : OAI22_X1 port map( A1 => n60206, A2 => n61203, B1 => n264, B2 => 
                           n15217, ZN => n11649);
   U4164 : OAI22_X1 port map( A1 => n60206, A2 => n61217, B1 => n263, B2 => 
                           n15217, ZN => n11650);
   U4165 : OAI22_X1 port map( A1 => n60207, A2 => n61231, B1 => n262, B2 => 
                           n15217, ZN => n11651);
   U4166 : OAI22_X1 port map( A1 => n60207, A2 => n61254, B1 => n261, B2 => 
                           n15217, ZN => n11652);
   U4167 : OAI22_X1 port map( A1 => n60196, A2 => n61147, B1 => n260, B2 => 
                           n60191, ZN => n11613);
   U4168 : OAI22_X1 port map( A1 => n60197, A2 => n61161, B1 => n259, B2 => 
                           n60191, ZN => n11614);
   U4169 : OAI22_X1 port map( A1 => n60197, A2 => n61175, B1 => n258, B2 => 
                           n60191, ZN => n11615);
   U4170 : OAI22_X1 port map( A1 => n60197, A2 => n61189, B1 => n257, B2 => 
                           n60191, ZN => n11616);
   U4171 : OAI22_X1 port map( A1 => n60197, A2 => n61203, B1 => n256, B2 => 
                           n15218, ZN => n11617);
   U4172 : OAI22_X1 port map( A1 => n60197, A2 => n61217, B1 => n255, B2 => 
                           n15218, ZN => n11618);
   U4173 : OAI22_X1 port map( A1 => n60198, A2 => n61231, B1 => n254, B2 => 
                           n15218, ZN => n11619);
   U4174 : OAI22_X1 port map( A1 => n60198, A2 => n61254, B1 => n253, B2 => 
                           n15218, ZN => n11620);
   U4175 : OAI22_X1 port map( A1 => n60187, A2 => n61147, B1 => n252, B2 => 
                           n60182, ZN => n11581);
   U4176 : OAI22_X1 port map( A1 => n60188, A2 => n61161, B1 => n251, B2 => 
                           n60182, ZN => n11582);
   U4177 : OAI22_X1 port map( A1 => n60188, A2 => n61175, B1 => n250, B2 => 
                           n60182, ZN => n11583);
   U4178 : OAI22_X1 port map( A1 => n60188, A2 => n61189, B1 => n249, B2 => 
                           n60182, ZN => n11584);
   U4179 : OAI22_X1 port map( A1 => n60188, A2 => n61203, B1 => n248, B2 => 
                           n15219, ZN => n11585);
   U4180 : OAI22_X1 port map( A1 => n60188, A2 => n61217, B1 => n247, B2 => 
                           n15219, ZN => n11586);
   U4181 : OAI22_X1 port map( A1 => n60189, A2 => n61231, B1 => n246, B2 => 
                           n15219, ZN => n11587);
   U4182 : OAI22_X1 port map( A1 => n60189, A2 => n61254, B1 => n245, B2 => 
                           n15219, ZN => n11588);
   U4183 : OAI22_X1 port map( A1 => n60124, A2 => n61147, B1 => n159, B2 => 
                           n60119, ZN => n11357);
   U4184 : OAI22_X1 port map( A1 => n60125, A2 => n61161, B1 => n158, B2 => 
                           n60119, ZN => n11358);
   U4185 : OAI22_X1 port map( A1 => n60125, A2 => n61175, B1 => n157, B2 => 
                           n60119, ZN => n11359);
   U4186 : OAI22_X1 port map( A1 => n60125, A2 => n61189, B1 => n156, B2 => 
                           n60119, ZN => n11360);
   U4187 : OAI22_X1 port map( A1 => n60125, A2 => n61203, B1 => n155, B2 => 
                           n15226, ZN => n11361);
   U4188 : OAI22_X1 port map( A1 => n60125, A2 => n61217, B1 => n154, B2 => 
                           n15226, ZN => n11362);
   U4189 : OAI22_X1 port map( A1 => n60126, A2 => n61231, B1 => n153, B2 => 
                           n15226, ZN => n11363);
   U4190 : OAI22_X1 port map( A1 => n60126, A2 => n61254, B1 => n152, B2 => 
                           n15226, ZN => n11364);
   U4191 : OAI22_X1 port map( A1 => n60115, A2 => n61147, B1 => n151, B2 => 
                           n60110, ZN => n11325);
   U4192 : OAI22_X1 port map( A1 => n60116, A2 => n61161, B1 => n150, B2 => 
                           n60110, ZN => n11326);
   U4193 : OAI22_X1 port map( A1 => n60116, A2 => n61175, B1 => n149, B2 => 
                           n60110, ZN => n11327);
   U4194 : OAI22_X1 port map( A1 => n60116, A2 => n61189, B1 => n148, B2 => 
                           n60110, ZN => n11328);
   U4195 : OAI22_X1 port map( A1 => n60116, A2 => n61203, B1 => n147, B2 => 
                           n15227, ZN => n11329);
   U4196 : OAI22_X1 port map( A1 => n60116, A2 => n61217, B1 => n146, B2 => 
                           n15227, ZN => n11330);
   U4197 : OAI22_X1 port map( A1 => n60117, A2 => n61231, B1 => n145, B2 => 
                           n15227, ZN => n11331);
   U4198 : OAI22_X1 port map( A1 => n60117, A2 => n61254, B1 => n144, B2 => 
                           n15227, ZN => n11332);
   U4199 : OAI22_X1 port map( A1 => n60736, A2 => n61142, B1 => n67, B2 => 
                           n60731, ZN => n13533);
   U4200 : OAI22_X1 port map( A1 => n60737, A2 => n61156, B1 => n66, B2 => 
                           n60731, ZN => n13534);
   U4201 : OAI22_X1 port map( A1 => n60737, A2 => n61170, B1 => n65, B2 => 
                           n60731, ZN => n13535);
   U4202 : OAI22_X1 port map( A1 => n60737, A2 => n61184, B1 => n64, B2 => 
                           n60731, ZN => n13536);
   U4203 : OAI22_X1 port map( A1 => n60737, A2 => n61198, B1 => n63, B2 => 
                           n15138, ZN => n13537);
   U4204 : OAI22_X1 port map( A1 => n60737, A2 => n61212, B1 => n62, B2 => 
                           n15138, ZN => n13538);
   U4205 : OAI22_X1 port map( A1 => n60738, A2 => n61226, B1 => n61, B2 => 
                           n15138, ZN => n13539);
   U4206 : OAI22_X1 port map( A1 => n60738, A2 => n61249, B1 => n60, B2 => 
                           n15138, ZN => n13540);
   U4207 : OAI22_X1 port map( A1 => n60727, A2 => n61142, B1 => n59, B2 => 
                           n60722, ZN => n13501);
   U4208 : OAI22_X1 port map( A1 => n60728, A2 => n61156, B1 => n58, B2 => 
                           n60722, ZN => n13502);
   U4209 : OAI22_X1 port map( A1 => n60728, A2 => n61170, B1 => n57, B2 => 
                           n60722, ZN => n13503);
   U4210 : OAI22_X1 port map( A1 => n60728, A2 => n61184, B1 => n56, B2 => 
                           n60722, ZN => n13504);
   U4211 : OAI22_X1 port map( A1 => n60728, A2 => n61198, B1 => n55, B2 => 
                           n15139, ZN => n13505);
   U4212 : OAI22_X1 port map( A1 => n60728, A2 => n61212, B1 => n54, B2 => 
                           n15139, ZN => n13506);
   U4213 : OAI22_X1 port map( A1 => n60729, A2 => n61226, B1 => n53, B2 => 
                           n15139, ZN => n13507);
   U4214 : OAI22_X1 port map( A1 => n60729, A2 => n61249, B1 => n52, B2 => 
                           n15139, ZN => n13508);
   U4215 : OAI22_X1 port map( A1 => n60700, A2 => n61142, B1 => n51, B2 => 
                           n60695, ZN => n13405);
   U4216 : OAI22_X1 port map( A1 => n60701, A2 => n61156, B1 => n50, B2 => 
                           n60695, ZN => n13406);
   U4217 : OAI22_X1 port map( A1 => n60701, A2 => n61170, B1 => n49, B2 => 
                           n60695, ZN => n13407);
   U4218 : OAI22_X1 port map( A1 => n60701, A2 => n61184, B1 => n48, B2 => 
                           n60695, ZN => n13408);
   U4219 : OAI22_X1 port map( A1 => n60701, A2 => n61198, B1 => n47, B2 => 
                           n15142, ZN => n13409);
   U4220 : OAI22_X1 port map( A1 => n60701, A2 => n61212, B1 => n46, B2 => 
                           n15142, ZN => n13410);
   U4221 : OAI22_X1 port map( A1 => n60702, A2 => n61226, B1 => n45, B2 => 
                           n15142, ZN => n13411);
   U4222 : OAI22_X1 port map( A1 => n60702, A2 => n61249, B1 => n44, B2 => 
                           n15142, ZN => n13412);
   U4223 : OAI22_X1 port map( A1 => n60691, A2 => n61142, B1 => n43, B2 => 
                           n60686, ZN => n13373);
   U4224 : OAI22_X1 port map( A1 => n60692, A2 => n61156, B1 => n42, B2 => 
                           n60686, ZN => n13374);
   U4225 : OAI22_X1 port map( A1 => n60692, A2 => n61170, B1 => n41, B2 => 
                           n60686, ZN => n13375);
   U4226 : OAI22_X1 port map( A1 => n60692, A2 => n61184, B1 => n40, B2 => 
                           n60686, ZN => n13376);
   U4227 : OAI22_X1 port map( A1 => n60692, A2 => n61198, B1 => n39, B2 => 
                           n15143, ZN => n13377);
   U4228 : OAI22_X1 port map( A1 => n60692, A2 => n61212, B1 => n38, B2 => 
                           n15143, ZN => n13378);
   U4229 : OAI22_X1 port map( A1 => n60693, A2 => n61226, B1 => n37, B2 => 
                           n15143, ZN => n13379);
   U4230 : OAI22_X1 port map( A1 => n60693, A2 => n61249, B1 => n36, B2 => 
                           n15143, ZN => n13380);
   U4231 : OAI22_X1 port map( A1 => n59800, A2 => n61150, B1 => n35, B2 => 
                           n59795, ZN => n10205);
   U4232 : OAI22_X1 port map( A1 => n59801, A2 => n61164, B1 => n34, B2 => 
                           n59795, ZN => n10206);
   U4233 : OAI22_X1 port map( A1 => n59801, A2 => n61178, B1 => n33, B2 => 
                           n59795, ZN => n10207);
   U4234 : OAI22_X1 port map( A1 => n59801, A2 => n61192, B1 => n32, B2 => 
                           n59795, ZN => n10208);
   U4235 : OAI22_X1 port map( A1 => n59801, A2 => n61206, B1 => n31, B2 => 
                           n15280, ZN => n10209);
   U4236 : OAI22_X1 port map( A1 => n59801, A2 => n61220, B1 => n30, B2 => 
                           n15280, ZN => n10210);
   U4237 : OAI22_X1 port map( A1 => n59802, A2 => n61234, B1 => n29, B2 => 
                           n15280, ZN => n10211);
   U4238 : OAI22_X1 port map( A1 => n59802, A2 => n61257, B1 => n28, B2 => 
                           n15280, ZN => n10212);
   U4239 : OAI22_X1 port map( A1 => n59791, A2 => n61150, B1 => n27, B2 => 
                           n59786, ZN => n10173);
   U4240 : OAI22_X1 port map( A1 => n59792, A2 => n61164, B1 => n26, B2 => 
                           n59786, ZN => n10174);
   U4241 : OAI22_X1 port map( A1 => n59792, A2 => n61178, B1 => n25, B2 => 
                           n59786, ZN => n10175);
   U4242 : OAI22_X1 port map( A1 => n59792, A2 => n61192, B1 => n24, B2 => 
                           n59786, ZN => n10176);
   U4243 : OAI22_X1 port map( A1 => n59792, A2 => n61206, B1 => n23, B2 => 
                           n15281, ZN => n10177);
   U4244 : OAI22_X1 port map( A1 => n59792, A2 => n61220, B1 => n22, B2 => 
                           n15281, ZN => n10178);
   U4245 : OAI22_X1 port map( A1 => n59793, A2 => n61234, B1 => n21, B2 => 
                           n15281, ZN => n10179);
   U4246 : OAI22_X1 port map( A1 => n59793, A2 => n61257, B1 => n20, B2 => 
                           n15281, ZN => n10180);
   U4247 : OAI22_X1 port map( A1 => n59782, A2 => n61150, B1 => n19, B2 => 
                           n59777, ZN => n10141);
   U4248 : OAI22_X1 port map( A1 => n59783, A2 => n61164, B1 => n18, B2 => 
                           n59777, ZN => n10142);
   U4249 : OAI22_X1 port map( A1 => n59783, A2 => n61178, B1 => n17, B2 => 
                           n59777, ZN => n10143);
   U4250 : OAI22_X1 port map( A1 => n59783, A2 => n61192, B1 => n16, B2 => 
                           n59777, ZN => n10144);
   U4251 : OAI22_X1 port map( A1 => n59783, A2 => n61206, B1 => n15, B2 => 
                           n15282, ZN => n10145);
   U4252 : OAI22_X1 port map( A1 => n59783, A2 => n61220, B1 => n14, B2 => 
                           n15282, ZN => n10146);
   U4253 : OAI22_X1 port map( A1 => n59784, A2 => n61234, B1 => n13, B2 => 
                           n15282, ZN => n10147);
   U4254 : OAI22_X1 port map( A1 => n59784, A2 => n61257, B1 => n12, B2 => 
                           n15282, ZN => n10148);
   U4255 : OAI22_X1 port map( A1 => n59773, A2 => n61151, B1 => n11, B2 => 
                           n59768, ZN => n10109);
   U4256 : OAI22_X1 port map( A1 => n59774, A2 => n61165, B1 => n10, B2 => 
                           n59768, ZN => n10110);
   U4257 : OAI22_X1 port map( A1 => n59774, A2 => n61179, B1 => n9, B2 => 
                           n59768, ZN => n10111);
   U4258 : OAI22_X1 port map( A1 => n59774, A2 => n61193, B1 => n8, B2 => 
                           n59768, ZN => n10112);
   U4259 : OAI22_X1 port map( A1 => n59774, A2 => n61207, B1 => n7, B2 => 
                           n15283, ZN => n10113);
   U4260 : OAI22_X1 port map( A1 => n59774, A2 => n61221, B1 => n6, B2 => 
                           n15283, ZN => n10114);
   U4261 : OAI22_X1 port map( A1 => n59775, A2 => n61235, B1 => n5, B2 => 
                           n15283, ZN => n10115);
   U4262 : OAI22_X1 port map( A1 => n59775, A2 => n61258, B1 => n4, B2 => 
                           n15283, ZN => n10116);
   U4263 : AOI22_X1 port map( A1 => n61906, A2 => n4364, B1 => n61904, B2 => 
                           n5010, ZN => n6738);
   U4264 : AOI22_X1 port map( A1 => n61906, A2 => n4363, B1 => n61904, B2 => 
                           n5009, ZN => n6663);
   U4265 : AOI22_X1 port map( A1 => n61906, A2 => n4362, B1 => n61904, B2 => 
                           n5008, ZN => n6588);
   U4266 : AOI22_X1 port map( A1 => n61906, A2 => n4361, B1 => n61904, B2 => 
                           n5007, ZN => n6513);
   U4267 : AOI22_X1 port map( A1 => n61906, A2 => n4360, B1 => n61904, B2 => 
                           n5006, ZN => n6438);
   U4268 : AOI22_X1 port map( A1 => n61906, A2 => n4359, B1 => n61903, B2 => 
                           n5005, ZN => n6363);
   U4269 : AOI22_X1 port map( A1 => n61906, A2 => n4358, B1 => n61903, B2 => 
                           n5004, ZN => n6288);
   U4270 : AOI22_X1 port map( A1 => n61906, A2 => n4357, B1 => n61903, B2 => 
                           n5003, ZN => n6213);
   U4271 : AOI22_X1 port map( A1 => n61906, A2 => n4356, B1 => n61903, B2 => 
                           n5002, ZN => n6138);
   U4272 : AOI22_X1 port map( A1 => n61907, A2 => n4369, B1 => n61904, B2 => 
                           n5015, ZN => n7113);
   U4273 : AOI22_X1 port map( A1 => n61907, A2 => n4368, B1 => n61904, B2 => 
                           n5014, ZN => n7038);
   U4274 : AOI22_X1 port map( A1 => n61906, A2 => n4366, B1 => n61904, B2 => 
                           n5012, ZN => n6888);
   U4275 : AOI22_X1 port map( A1 => n61906, A2 => n4365, B1 => n61904, B2 => 
                           n5011, ZN => n6813);
   U4276 : AOI22_X1 port map( A1 => n61907, A2 => n4371, B1 => n61904, B2 => 
                           n5017, ZN => n7263);
   U4277 : AOI22_X1 port map( A1 => n61906, A2 => n4378, B1 => n61905, B2 => 
                           n5025, ZN => n7882);
   U4278 : AOI22_X1 port map( A1 => n61907, A2 => n4377, B1 => n61905, B2 => 
                           n5024, ZN => n7788);
   U4279 : AOI22_X1 port map( A1 => n61907, A2 => n4376, B1 => n61905, B2 => 
                           n5023, ZN => n7713);
   U4280 : AOI22_X1 port map( A1 => n61907, A2 => n4375, B1 => n61905, B2 => 
                           n5022, ZN => n7638);
   U4281 : AOI22_X1 port map( A1 => n61907, A2 => n4374, B1 => n61905, B2 => 
                           n5020, ZN => n7488);
   U4282 : AOI22_X1 port map( A1 => n61907, A2 => n4373, B1 => n61905, B2 => 
                           n5019, ZN => n7413);
   U4283 : AOI22_X1 port map( A1 => n61907, A2 => n4372, B1 => n61904, B2 => 
                           n5018, ZN => n7338);
   U4284 : AOI22_X1 port map( A1 => n61907, A2 => n4370, B1 => n61904, B2 => 
                           n5016, ZN => n7188);
   U4285 : AOI22_X1 port map( A1 => n61544, A2 => n4945, B1 => n61542, B2 => 
                           n4921, ZN => n14393);
   U4286 : AOI22_X1 port map( A1 => n61646, A2 => n4639, B1 => n61644, B2 => 
                           n4447, ZN => n14377);
   U4287 : AOI22_X1 port map( A1 => n61544, A2 => n4944, B1 => n61542, B2 => 
                           n4920, ZN => n9902);
   U4288 : AOI22_X1 port map( A1 => n61646, A2 => n4638, B1 => n61644, B2 => 
                           n4446, ZN => n9886);
   U4289 : AOI22_X1 port map( A1 => n61544, A2 => n4943, B1 => n61542, B2 => 
                           n4919, ZN => n9827);
   U4290 : AOI22_X1 port map( A1 => n61646, A2 => n4637, B1 => n61644, B2 => 
                           n4445, ZN => n9811);
   U4291 : AOI22_X1 port map( A1 => n61544, A2 => n4942, B1 => n61542, B2 => 
                           n4918, ZN => n9688);
   U4292 : AOI22_X1 port map( A1 => n61646, A2 => n4636, B1 => n61644, B2 => 
                           n4444, ZN => n9672);
   U4293 : AOI22_X1 port map( A1 => n61545, A2 => n4941, B1 => n61542, B2 => 
                           n4917, ZN => n9597);
   U4294 : AOI22_X1 port map( A1 => n61647, A2 => n4635, B1 => n61644, B2 => 
                           n4443, ZN => n9581);
   U4295 : AOI22_X1 port map( A1 => n61545, A2 => n4940, B1 => n61542, B2 => 
                           n4916, ZN => n9522);
   U4296 : AOI22_X1 port map( A1 => n61647, A2 => n4634, B1 => n61644, B2 => 
                           n4442, ZN => n9506);
   U4297 : AOI22_X1 port map( A1 => n61545, A2 => n4939, B1 => n61542, B2 => 
                           n4915, ZN => n9447);
   U4298 : AOI22_X1 port map( A1 => n61647, A2 => n4633, B1 => n61644, B2 => 
                           n4441, ZN => n9431);
   U4299 : AOI22_X1 port map( A1 => n61545, A2 => n4938, B1 => n61542, B2 => 
                           n4914, ZN => n9372);
   U4300 : AOI22_X1 port map( A1 => n61647, A2 => n4632, B1 => n61644, B2 => 
                           n4440, ZN => n9356);
   U4301 : AOI22_X1 port map( A1 => n61545, A2 => n4937, B1 => n61542, B2 => 
                           n4913, ZN => n9233);
   U4302 : AOI22_X1 port map( A1 => n61647, A2 => n4631, B1 => n61644, B2 => 
                           n4439, ZN => n9217);
   U4303 : AOI22_X1 port map( A1 => n61545, A2 => n4936, B1 => n61542, B2 => 
                           n4912, ZN => n9158);
   U4304 : AOI22_X1 port map( A1 => n61647, A2 => n4630, B1 => n61644, B2 => 
                           n4438, ZN => n9142);
   U4305 : AOI22_X1 port map( A1 => n61545, A2 => n4935, B1 => n61542, B2 => 
                           n4911, ZN => n9083);
   U4306 : AOI22_X1 port map( A1 => n61647, A2 => n4629, B1 => n61644, B2 => 
                           n4437, ZN => n9067);
   U4307 : AOI22_X1 port map( A1 => n61545, A2 => n4934, B1 => n61542, B2 => 
                           n4910, ZN => n9008);
   U4308 : AOI22_X1 port map( A1 => n61647, A2 => n4628, B1 => n61644, B2 => 
                           n4436, ZN => n8992);
   U4309 : AOI22_X1 port map( A1 => n61545, A2 => n4933, B1 => n61541, B2 => 
                           n4909, ZN => n8933);
   U4310 : AOI22_X1 port map( A1 => n61647, A2 => n4627, B1 => n61643, B2 => 
                           n4435, ZN => n8917);
   U4311 : AOI22_X1 port map( A1 => n61545, A2 => n4932, B1 => n61541, B2 => 
                           n4908, ZN => n8858);
   U4312 : AOI22_X1 port map( A1 => n61647, A2 => n4626, B1 => n61643, B2 => 
                           n4434, ZN => n8842);
   U4313 : AOI22_X1 port map( A1 => n61545, A2 => n4931, B1 => n61541, B2 => 
                           n4907, ZN => n8783);
   U4314 : AOI22_X1 port map( A1 => n61647, A2 => n4625, B1 => n61643, B2 => 
                           n4433, ZN => n8767);
   U4315 : AOI22_X1 port map( A1 => n61545, A2 => n4930, B1 => n61541, B2 => 
                           n4906, ZN => n8708);
   U4316 : AOI22_X1 port map( A1 => n61647, A2 => n4624, B1 => n61643, B2 => 
                           n4432, ZN => n8692);
   U4317 : AOI22_X1 port map( A1 => n61544, A2 => n4953, B1 => n61543, B2 => 
                           n4929, ZN => n15011);
   U4318 : AOI22_X1 port map( A1 => n61646, A2 => n4647, B1 => n61645, B2 => 
                           n4455, ZN => n14982);
   U4319 : AOI22_X1 port map( A1 => n61544, A2 => n4952, B1 => n61543, B2 => 
                           n4928, ZN => n14918);
   U4320 : AOI22_X1 port map( A1 => n61646, A2 => n4646, B1 => n61645, B2 => 
                           n4454, ZN => n14902);
   U4321 : AOI22_X1 port map( A1 => n61544, A2 => n4951, B1 => n61543, B2 => 
                           n4927, ZN => n14843);
   U4322 : AOI22_X1 port map( A1 => n61646, A2 => n4645, B1 => n61645, B2 => 
                           n4453, ZN => n14827);
   U4323 : AOI22_X1 port map( A1 => n61544, A2 => n4950, B1 => n61543, B2 => 
                           n4926, ZN => n14768);
   U4324 : AOI22_X1 port map( A1 => n61646, A2 => n4644, B1 => n61645, B2 => 
                           n4452, ZN => n14752);
   U4325 : AOI22_X1 port map( A1 => n61544, A2 => n4949, B1 => n61543, B2 => 
                           n4925, ZN => n14693);
   U4326 : AOI22_X1 port map( A1 => n61646, A2 => n4643, B1 => n61645, B2 => 
                           n4451, ZN => n14677);
   U4327 : AOI22_X1 port map( A1 => n61544, A2 => n4948, B1 => n61543, B2 => 
                           n4924, ZN => n14618);
   U4328 : AOI22_X1 port map( A1 => n61646, A2 => n4642, B1 => n61645, B2 => 
                           n4450, ZN => n14602);
   U4329 : AOI22_X1 port map( A1 => n61544, A2 => n4947, B1 => n61543, B2 => 
                           n4923, ZN => n14543);
   U4330 : AOI22_X1 port map( A1 => n61646, A2 => n4641, B1 => n61645, B2 => 
                           n4449, ZN => n14527);
   U4331 : AOI22_X1 port map( A1 => n61544, A2 => n4946, B1 => n61543, B2 => 
                           n4922, ZN => n14468);
   U4332 : AOI22_X1 port map( A1 => n61646, A2 => n4640, B1 => n61645, B2 => 
                           n4448, ZN => n14452);
   U4333 : AOI22_X1 port map( A1 => n61907, A2 => n4367, B1 => n61904, B2 => 
                           n5013, ZN => n6963);
   U4334 : OAI22_X1 port map( A1 => n60543, A2 => n61968, B1 => n4857, B2 => 
                           n60542, ZN => n12837);
   U4335 : OAI22_X1 port map( A1 => n60543, A2 => n61982, B1 => n4856, B2 => 
                           n60542, ZN => n12838);
   U4336 : OAI22_X1 port map( A1 => n60543, A2 => n61996, B1 => n4855, B2 => 
                           n60542, ZN => n12839);
   U4337 : OAI22_X1 port map( A1 => n60543, A2 => n62010, B1 => n4854, B2 => 
                           n60542, ZN => n12840);
   U4338 : OAI22_X1 port map( A1 => n60543, A2 => n62024, B1 => n4853, B2 => 
                           n60542, ZN => n12841);
   U4339 : OAI22_X1 port map( A1 => n60544, A2 => n62038, B1 => n4852, B2 => 
                           n60542, ZN => n12842);
   U4340 : OAI22_X1 port map( A1 => n60544, A2 => n62052, B1 => n4851, B2 => 
                           n60542, ZN => n12843);
   U4341 : OAI22_X1 port map( A1 => n60544, A2 => n62066, B1 => n4850, B2 => 
                           n60542, ZN => n12844);
   U4342 : OAI22_X1 port map( A1 => n60544, A2 => n62080, B1 => n4849, B2 => 
                           n60542, ZN => n12845);
   U4343 : OAI22_X1 port map( A1 => n60544, A2 => n62094, B1 => n4848, B2 => 
                           n60542, ZN => n12846);
   U4344 : OAI22_X1 port map( A1 => n60545, A2 => n62108, B1 => n4847, B2 => 
                           n60542, ZN => n12847);
   U4345 : OAI22_X1 port map( A1 => n60545, A2 => n60961, B1 => n4846, B2 => 
                           n60542, ZN => n12848);
   U4346 : OAI22_X1 port map( A1 => n60545, A2 => n60975, B1 => n4845, B2 => 
                           n15161, ZN => n12849);
   U4347 : OAI22_X1 port map( A1 => n60545, A2 => n60989, B1 => n4844, B2 => 
                           n15161, ZN => n12850);
   U4348 : OAI22_X1 port map( A1 => n60545, A2 => n61003, B1 => n4843, B2 => 
                           n15161, ZN => n12851);
   U4349 : OAI22_X1 port map( A1 => n60546, A2 => n61017, B1 => n4842, B2 => 
                           n15161, ZN => n12852);
   U4350 : OAI22_X1 port map( A1 => n60546, A2 => n61031, B1 => n4841, B2 => 
                           n15161, ZN => n12853);
   U4351 : OAI22_X1 port map( A1 => n60546, A2 => n61045, B1 => n4840, B2 => 
                           n15161, ZN => n12854);
   U4352 : OAI22_X1 port map( A1 => n60546, A2 => n61059, B1 => n4839, B2 => 
                           n15161, ZN => n12855);
   U4353 : OAI22_X1 port map( A1 => n60546, A2 => n61073, B1 => n4838, B2 => 
                           n60542, ZN => n12856);
   U4354 : OAI22_X1 port map( A1 => n60547, A2 => n61087, B1 => n4837, B2 => 
                           n60542, ZN => n12857);
   U4355 : OAI22_X1 port map( A1 => n60547, A2 => n61101, B1 => n4836, B2 => 
                           n60542, ZN => n12858);
   U4356 : OAI22_X1 port map( A1 => n60547, A2 => n61115, B1 => n4835, B2 => 
                           n60542, ZN => n12859);
   U4357 : OAI22_X1 port map( A1 => n60547, A2 => n61129, B1 => n4834, B2 => 
                           n60542, ZN => n12860);
   U4358 : OAI22_X1 port map( A1 => n60536, A2 => n61003, B1 => n4833, B2 => 
                           n15162, ZN => n12819);
   U4359 : OAI22_X1 port map( A1 => n60537, A2 => n61017, B1 => n4832, B2 => 
                           n15162, ZN => n12820);
   U4360 : OAI22_X1 port map( A1 => n60537, A2 => n61031, B1 => n4831, B2 => 
                           n15162, ZN => n12821);
   U4361 : OAI22_X1 port map( A1 => n60537, A2 => n61045, B1 => n4830, B2 => 
                           n15162, ZN => n12822);
   U4362 : OAI22_X1 port map( A1 => n60537, A2 => n61059, B1 => n4829, B2 => 
                           n15162, ZN => n12823);
   U4363 : OAI22_X1 port map( A1 => n60537, A2 => n61073, B1 => n4828, B2 => 
                           n15162, ZN => n12824);
   U4364 : OAI22_X1 port map( A1 => n60538, A2 => n61087, B1 => n4827, B2 => 
                           n15162, ZN => n12825);
   U4365 : OAI22_X1 port map( A1 => n60538, A2 => n61101, B1 => n4826, B2 => 
                           n60533, ZN => n12826);
   U4366 : OAI22_X1 port map( A1 => n60538, A2 => n61115, B1 => n4825, B2 => 
                           n60533, ZN => n12827);
   U4367 : OAI22_X1 port map( A1 => n60538, A2 => n61129, B1 => n4824, B2 => 
                           n60533, ZN => n12828);
   U4368 : OAI22_X1 port map( A1 => n60498, A2 => n61969, B1 => n4785, B2 => 
                           n60497, ZN => n12677);
   U4369 : OAI22_X1 port map( A1 => n60498, A2 => n61983, B1 => n4784, B2 => 
                           n60497, ZN => n12678);
   U4370 : OAI22_X1 port map( A1 => n60498, A2 => n61997, B1 => n4783, B2 => 
                           n60497, ZN => n12679);
   U4371 : OAI22_X1 port map( A1 => n60498, A2 => n62011, B1 => n4782, B2 => 
                           n60497, ZN => n12680);
   U4372 : OAI22_X1 port map( A1 => n60498, A2 => n62025, B1 => n4781, B2 => 
                           n60497, ZN => n12681);
   U4373 : OAI22_X1 port map( A1 => n60499, A2 => n62039, B1 => n4780, B2 => 
                           n60497, ZN => n12682);
   U4374 : OAI22_X1 port map( A1 => n60499, A2 => n62053, B1 => n4779, B2 => 
                           n60497, ZN => n12683);
   U4375 : OAI22_X1 port map( A1 => n60499, A2 => n62067, B1 => n4778, B2 => 
                           n60497, ZN => n12684);
   U4376 : OAI22_X1 port map( A1 => n60499, A2 => n62081, B1 => n4777, B2 => 
                           n60497, ZN => n12685);
   U4377 : OAI22_X1 port map( A1 => n60499, A2 => n62095, B1 => n4776, B2 => 
                           n60497, ZN => n12686);
   U4378 : OAI22_X1 port map( A1 => n60500, A2 => n62109, B1 => n4775, B2 => 
                           n60497, ZN => n12687);
   U4379 : OAI22_X1 port map( A1 => n60500, A2 => n60962, B1 => n4774, B2 => 
                           n60497, ZN => n12688);
   U4380 : OAI22_X1 port map( A1 => n60500, A2 => n60976, B1 => n4773, B2 => 
                           n15167, ZN => n12689);
   U4381 : OAI22_X1 port map( A1 => n60500, A2 => n60990, B1 => n4772, B2 => 
                           n15167, ZN => n12690);
   U4382 : OAI22_X1 port map( A1 => n60500, A2 => n61004, B1 => n4771, B2 => 
                           n15167, ZN => n12691);
   U4383 : OAI22_X1 port map( A1 => n60501, A2 => n61018, B1 => n4770, B2 => 
                           n15167, ZN => n12692);
   U4384 : OAI22_X1 port map( A1 => n60501, A2 => n61032, B1 => n4769, B2 => 
                           n15167, ZN => n12693);
   U4385 : OAI22_X1 port map( A1 => n60501, A2 => n61046, B1 => n4768, B2 => 
                           n15167, ZN => n12694);
   U4386 : OAI22_X1 port map( A1 => n60501, A2 => n61060, B1 => n4767, B2 => 
                           n15167, ZN => n12695);
   U4387 : OAI22_X1 port map( A1 => n60501, A2 => n61074, B1 => n4766, B2 => 
                           n60497, ZN => n12696);
   U4388 : OAI22_X1 port map( A1 => n60502, A2 => n61088, B1 => n4765, B2 => 
                           n60497, ZN => n12697);
   U4389 : OAI22_X1 port map( A1 => n60502, A2 => n61102, B1 => n4764, B2 => 
                           n60497, ZN => n12698);
   U4390 : OAI22_X1 port map( A1 => n60502, A2 => n61116, B1 => n4763, B2 => 
                           n60497, ZN => n12699);
   U4391 : OAI22_X1 port map( A1 => n60502, A2 => n61130, B1 => n4762, B2 => 
                           n60497, ZN => n12700);
   U4392 : OAI22_X1 port map( A1 => n60489, A2 => n61969, B1 => n4761, B2 => 
                           n60488, ZN => n12645);
   U4393 : OAI22_X1 port map( A1 => n60489, A2 => n61983, B1 => n4760, B2 => 
                           n60488, ZN => n12646);
   U4394 : OAI22_X1 port map( A1 => n60489, A2 => n61997, B1 => n4759, B2 => 
                           n60488, ZN => n12647);
   U4395 : OAI22_X1 port map( A1 => n60489, A2 => n62011, B1 => n4758, B2 => 
                           n60488, ZN => n12648);
   U4396 : OAI22_X1 port map( A1 => n60489, A2 => n62025, B1 => n4757, B2 => 
                           n60488, ZN => n12649);
   U4397 : OAI22_X1 port map( A1 => n60490, A2 => n62039, B1 => n4756, B2 => 
                           n60488, ZN => n12650);
   U4398 : OAI22_X1 port map( A1 => n60490, A2 => n62053, B1 => n4755, B2 => 
                           n60488, ZN => n12651);
   U4399 : OAI22_X1 port map( A1 => n60490, A2 => n62067, B1 => n4754, B2 => 
                           n60488, ZN => n12652);
   U4400 : OAI22_X1 port map( A1 => n60490, A2 => n62081, B1 => n4753, B2 => 
                           n60488, ZN => n12653);
   U4401 : OAI22_X1 port map( A1 => n60490, A2 => n62095, B1 => n4752, B2 => 
                           n60488, ZN => n12654);
   U4402 : OAI22_X1 port map( A1 => n60491, A2 => n62109, B1 => n4751, B2 => 
                           n60488, ZN => n12655);
   U4403 : OAI22_X1 port map( A1 => n60491, A2 => n60962, B1 => n4750, B2 => 
                           n60488, ZN => n12656);
   U4404 : OAI22_X1 port map( A1 => n60491, A2 => n60976, B1 => n4749, B2 => 
                           n15168, ZN => n12657);
   U4405 : OAI22_X1 port map( A1 => n60491, A2 => n60990, B1 => n4748, B2 => 
                           n15168, ZN => n12658);
   U4406 : OAI22_X1 port map( A1 => n60491, A2 => n61004, B1 => n4747, B2 => 
                           n15168, ZN => n12659);
   U4407 : OAI22_X1 port map( A1 => n60492, A2 => n61018, B1 => n4746, B2 => 
                           n15168, ZN => n12660);
   U4408 : OAI22_X1 port map( A1 => n60492, A2 => n61032, B1 => n4745, B2 => 
                           n15168, ZN => n12661);
   U4409 : OAI22_X1 port map( A1 => n60492, A2 => n61046, B1 => n4744, B2 => 
                           n15168, ZN => n12662);
   U4410 : OAI22_X1 port map( A1 => n60492, A2 => n61060, B1 => n4743, B2 => 
                           n15168, ZN => n12663);
   U4411 : OAI22_X1 port map( A1 => n60492, A2 => n61074, B1 => n4742, B2 => 
                           n60488, ZN => n12664);
   U4412 : OAI22_X1 port map( A1 => n60493, A2 => n61088, B1 => n4741, B2 => 
                           n60488, ZN => n12665);
   U4413 : OAI22_X1 port map( A1 => n60493, A2 => n61102, B1 => n4740, B2 => 
                           n60488, ZN => n12666);
   U4414 : OAI22_X1 port map( A1 => n60493, A2 => n61116, B1 => n4739, B2 => 
                           n60488, ZN => n12667);
   U4415 : OAI22_X1 port map( A1 => n60493, A2 => n61130, B1 => n4738, B2 => 
                           n60488, ZN => n12668);
   U4416 : OAI22_X1 port map( A1 => n60426, A2 => n61969, B1 => n4737, B2 => 
                           n60425, ZN => n12421);
   U4417 : OAI22_X1 port map( A1 => n60426, A2 => n61983, B1 => n4736, B2 => 
                           n60425, ZN => n12422);
   U4418 : OAI22_X1 port map( A1 => n60426, A2 => n61997, B1 => n4735, B2 => 
                           n60425, ZN => n12423);
   U4419 : OAI22_X1 port map( A1 => n60426, A2 => n62011, B1 => n4734, B2 => 
                           n60425, ZN => n12424);
   U4420 : OAI22_X1 port map( A1 => n60426, A2 => n62025, B1 => n4733, B2 => 
                           n60425, ZN => n12425);
   U4421 : OAI22_X1 port map( A1 => n60427, A2 => n62039, B1 => n4732, B2 => 
                           n60425, ZN => n12426);
   U4422 : OAI22_X1 port map( A1 => n60427, A2 => n62053, B1 => n4731, B2 => 
                           n60425, ZN => n12427);
   U4423 : OAI22_X1 port map( A1 => n60427, A2 => n62067, B1 => n4730, B2 => 
                           n60425, ZN => n12428);
   U4424 : OAI22_X1 port map( A1 => n60427, A2 => n62081, B1 => n4729, B2 => 
                           n60425, ZN => n12429);
   U4425 : OAI22_X1 port map( A1 => n60427, A2 => n62095, B1 => n4728, B2 => 
                           n60425, ZN => n12430);
   U4426 : OAI22_X1 port map( A1 => n60428, A2 => n62109, B1 => n4727, B2 => 
                           n60425, ZN => n12431);
   U4427 : OAI22_X1 port map( A1 => n60428, A2 => n60962, B1 => n4726, B2 => 
                           n60425, ZN => n12432);
   U4428 : OAI22_X1 port map( A1 => n60428, A2 => n60976, B1 => n4725, B2 => 
                           n15182, ZN => n12433);
   U4429 : OAI22_X1 port map( A1 => n60428, A2 => n60990, B1 => n4724, B2 => 
                           n15182, ZN => n12434);
   U4430 : OAI22_X1 port map( A1 => n60428, A2 => n61004, B1 => n4723, B2 => 
                           n15182, ZN => n12435);
   U4431 : OAI22_X1 port map( A1 => n60429, A2 => n61018, B1 => n4722, B2 => 
                           n15182, ZN => n12436);
   U4432 : OAI22_X1 port map( A1 => n60429, A2 => n61032, B1 => n4721, B2 => 
                           n15182, ZN => n12437);
   U4433 : OAI22_X1 port map( A1 => n60429, A2 => n61046, B1 => n4720, B2 => 
                           n15182, ZN => n12438);
   U4434 : OAI22_X1 port map( A1 => n60429, A2 => n61060, B1 => n4719, B2 => 
                           n15182, ZN => n12439);
   U4435 : OAI22_X1 port map( A1 => n60429, A2 => n61074, B1 => n4718, B2 => 
                           n60425, ZN => n12440);
   U4436 : OAI22_X1 port map( A1 => n60430, A2 => n61088, B1 => n4717, B2 => 
                           n60425, ZN => n12441);
   U4437 : OAI22_X1 port map( A1 => n60430, A2 => n61102, B1 => n4716, B2 => 
                           n60425, ZN => n12442);
   U4438 : OAI22_X1 port map( A1 => n60430, A2 => n61116, B1 => n4715, B2 => 
                           n60425, ZN => n12443);
   U4439 : OAI22_X1 port map( A1 => n60430, A2 => n61130, B1 => n4714, B2 => 
                           n60425, ZN => n12444);
   U4440 : OAI22_X1 port map( A1 => n60921, A2 => n61965, B1 => n4695, B2 => 
                           n60920, ZN => n14181);
   U4441 : OAI22_X1 port map( A1 => n60921, A2 => n61979, B1 => n4694, B2 => 
                           n60920, ZN => n14182);
   U4442 : OAI22_X1 port map( A1 => n60921, A2 => n61993, B1 => n4693, B2 => 
                           n60920, ZN => n14183);
   U4443 : OAI22_X1 port map( A1 => n60921, A2 => n62007, B1 => n4692, B2 => 
                           n60920, ZN => n14184);
   U4444 : OAI22_X1 port map( A1 => n60921, A2 => n62021, B1 => n4691, B2 => 
                           n60920, ZN => n14185);
   U4445 : OAI22_X1 port map( A1 => n60922, A2 => n62035, B1 => n4690, B2 => 
                           n60920, ZN => n14186);
   U4446 : OAI22_X1 port map( A1 => n60922, A2 => n62049, B1 => n4689, B2 => 
                           n60920, ZN => n14187);
   U4447 : OAI22_X1 port map( A1 => n60922, A2 => n62063, B1 => n4688, B2 => 
                           n60920, ZN => n14188);
   U4448 : OAI22_X1 port map( A1 => n60922, A2 => n62077, B1 => n4687, B2 => 
                           n60920, ZN => n14189);
   U4449 : OAI22_X1 port map( A1 => n60922, A2 => n62091, B1 => n4686, B2 => 
                           n60920, ZN => n14190);
   U4450 : OAI22_X1 port map( A1 => n60923, A2 => n62105, B1 => n4685, B2 => 
                           n60920, ZN => n14191);
   U4451 : OAI22_X1 port map( A1 => n60923, A2 => n60958, B1 => n4684, B2 => 
                           n60920, ZN => n14192);
   U4452 : OAI22_X1 port map( A1 => n60923, A2 => n60972, B1 => n4683, B2 => 
                           n15102, ZN => n14193);
   U4453 : OAI22_X1 port map( A1 => n60923, A2 => n60986, B1 => n4682, B2 => 
                           n15102, ZN => n14194);
   U4454 : OAI22_X1 port map( A1 => n60923, A2 => n61000, B1 => n4681, B2 => 
                           n15102, ZN => n14195);
   U4455 : OAI22_X1 port map( A1 => n60924, A2 => n61014, B1 => n4680, B2 => 
                           n15102, ZN => n14196);
   U4456 : OAI22_X1 port map( A1 => n60924, A2 => n61028, B1 => n4679, B2 => 
                           n15102, ZN => n14197);
   U4457 : OAI22_X1 port map( A1 => n60924, A2 => n61042, B1 => n4678, B2 => 
                           n15102, ZN => n14198);
   U4458 : OAI22_X1 port map( A1 => n60924, A2 => n61056, B1 => n4677, B2 => 
                           n15102, ZN => n14199);
   U4459 : OAI22_X1 port map( A1 => n60924, A2 => n61070, B1 => n4676, B2 => 
                           n60920, ZN => n14200);
   U4460 : OAI22_X1 port map( A1 => n60925, A2 => n61084, B1 => n4675, B2 => 
                           n60920, ZN => n14201);
   U4461 : OAI22_X1 port map( A1 => n60925, A2 => n61098, B1 => n4674, B2 => 
                           n60920, ZN => n14202);
   U4462 : OAI22_X1 port map( A1 => n60925, A2 => n61112, B1 => n4673, B2 => 
                           n60920, ZN => n14203);
   U4463 : OAI22_X1 port map( A1 => n60925, A2 => n61126, B1 => n4672, B2 => 
                           n60920, ZN => n14204);
   U4464 : OAI22_X1 port map( A1 => n60912, A2 => n61965, B1 => n4671, B2 => 
                           n60911, ZN => n14149);
   U4465 : OAI22_X1 port map( A1 => n60912, A2 => n61979, B1 => n4670, B2 => 
                           n60911, ZN => n14150);
   U4466 : OAI22_X1 port map( A1 => n60912, A2 => n61993, B1 => n4669, B2 => 
                           n60911, ZN => n14151);
   U4467 : OAI22_X1 port map( A1 => n60912, A2 => n62007, B1 => n4668, B2 => 
                           n60911, ZN => n14152);
   U4468 : OAI22_X1 port map( A1 => n60912, A2 => n62021, B1 => n4667, B2 => 
                           n60911, ZN => n14153);
   U4469 : OAI22_X1 port map( A1 => n60913, A2 => n62035, B1 => n4666, B2 => 
                           n60911, ZN => n14154);
   U4470 : OAI22_X1 port map( A1 => n60913, A2 => n62049, B1 => n4665, B2 => 
                           n60911, ZN => n14155);
   U4471 : OAI22_X1 port map( A1 => n60913, A2 => n62063, B1 => n4664, B2 => 
                           n60911, ZN => n14156);
   U4472 : OAI22_X1 port map( A1 => n60913, A2 => n62077, B1 => n4663, B2 => 
                           n60911, ZN => n14157);
   U4473 : OAI22_X1 port map( A1 => n60913, A2 => n62091, B1 => n4662, B2 => 
                           n60911, ZN => n14158);
   U4474 : OAI22_X1 port map( A1 => n60914, A2 => n62105, B1 => n4661, B2 => 
                           n60911, ZN => n14159);
   U4475 : OAI22_X1 port map( A1 => n60914, A2 => n60958, B1 => n4660, B2 => 
                           n60911, ZN => n14160);
   U4476 : OAI22_X1 port map( A1 => n60914, A2 => n60972, B1 => n4659, B2 => 
                           n15104, ZN => n14161);
   U4477 : OAI22_X1 port map( A1 => n60914, A2 => n60986, B1 => n4658, B2 => 
                           n15104, ZN => n14162);
   U4478 : OAI22_X1 port map( A1 => n60914, A2 => n61000, B1 => n4657, B2 => 
                           n15104, ZN => n14163);
   U4479 : OAI22_X1 port map( A1 => n60915, A2 => n61014, B1 => n4656, B2 => 
                           n15104, ZN => n14164);
   U4480 : OAI22_X1 port map( A1 => n60915, A2 => n61028, B1 => n4655, B2 => 
                           n15104, ZN => n14165);
   U4481 : OAI22_X1 port map( A1 => n60915, A2 => n61042, B1 => n4654, B2 => 
                           n15104, ZN => n14166);
   U4482 : OAI22_X1 port map( A1 => n60915, A2 => n61056, B1 => n4653, B2 => 
                           n15104, ZN => n14167);
   U4483 : OAI22_X1 port map( A1 => n60915, A2 => n61070, B1 => n4652, B2 => 
                           n60911, ZN => n14168);
   U4484 : OAI22_X1 port map( A1 => n60916, A2 => n61084, B1 => n4651, B2 => 
                           n60911, ZN => n14169);
   U4485 : OAI22_X1 port map( A1 => n60916, A2 => n61098, B1 => n4650, B2 => 
                           n60911, ZN => n14170);
   U4486 : OAI22_X1 port map( A1 => n60916, A2 => n61112, B1 => n4649, B2 => 
                           n60911, ZN => n14171);
   U4487 : OAI22_X1 port map( A1 => n60916, A2 => n61126, B1 => n4648, B2 => 
                           n60911, ZN => n14172);
   U4488 : OAI22_X1 port map( A1 => n60885, A2 => n61965, B1 => n4623, B2 => 
                           n60884, ZN => n14053);
   U4489 : OAI22_X1 port map( A1 => n60885, A2 => n61979, B1 => n4622, B2 => 
                           n60884, ZN => n14054);
   U4490 : OAI22_X1 port map( A1 => n60885, A2 => n61993, B1 => n4621, B2 => 
                           n60884, ZN => n14055);
   U4491 : OAI22_X1 port map( A1 => n60885, A2 => n62007, B1 => n4620, B2 => 
                           n60884, ZN => n14056);
   U4492 : OAI22_X1 port map( A1 => n60885, A2 => n62021, B1 => n4619, B2 => 
                           n60884, ZN => n14057);
   U4493 : OAI22_X1 port map( A1 => n60886, A2 => n62035, B1 => n4618, B2 => 
                           n60884, ZN => n14058);
   U4494 : OAI22_X1 port map( A1 => n60886, A2 => n62049, B1 => n4617, B2 => 
                           n60884, ZN => n14059);
   U4495 : OAI22_X1 port map( A1 => n60886, A2 => n62063, B1 => n4616, B2 => 
                           n60884, ZN => n14060);
   U4496 : OAI22_X1 port map( A1 => n60886, A2 => n62077, B1 => n4615, B2 => 
                           n60884, ZN => n14061);
   U4497 : OAI22_X1 port map( A1 => n60886, A2 => n62091, B1 => n4614, B2 => 
                           n60884, ZN => n14062);
   U4498 : OAI22_X1 port map( A1 => n60887, A2 => n62105, B1 => n4613, B2 => 
                           n60884, ZN => n14063);
   U4499 : OAI22_X1 port map( A1 => n60887, A2 => n60958, B1 => n4612, B2 => 
                           n60884, ZN => n14064);
   U4500 : OAI22_X1 port map( A1 => n60887, A2 => n60972, B1 => n4611, B2 => 
                           n15110, ZN => n14065);
   U4501 : OAI22_X1 port map( A1 => n60887, A2 => n60986, B1 => n4610, B2 => 
                           n15110, ZN => n14066);
   U4502 : OAI22_X1 port map( A1 => n60887, A2 => n61000, B1 => n4609, B2 => 
                           n15110, ZN => n14067);
   U4503 : OAI22_X1 port map( A1 => n60888, A2 => n61014, B1 => n4608, B2 => 
                           n15110, ZN => n14068);
   U4504 : OAI22_X1 port map( A1 => n60888, A2 => n61028, B1 => n4607, B2 => 
                           n15110, ZN => n14069);
   U4505 : OAI22_X1 port map( A1 => n60888, A2 => n61042, B1 => n4606, B2 => 
                           n15110, ZN => n14070);
   U4506 : OAI22_X1 port map( A1 => n60888, A2 => n61056, B1 => n4605, B2 => 
                           n15110, ZN => n14071);
   U4507 : OAI22_X1 port map( A1 => n60888, A2 => n61070, B1 => n4604, B2 => 
                           n60884, ZN => n14072);
   U4508 : OAI22_X1 port map( A1 => n60889, A2 => n61084, B1 => n4603, B2 => 
                           n60884, ZN => n14073);
   U4509 : OAI22_X1 port map( A1 => n60889, A2 => n61098, B1 => n4602, B2 => 
                           n60884, ZN => n14074);
   U4510 : OAI22_X1 port map( A1 => n60889, A2 => n61112, B1 => n4601, B2 => 
                           n60884, ZN => n14075);
   U4511 : OAI22_X1 port map( A1 => n60889, A2 => n61126, B1 => n4600, B2 => 
                           n60884, ZN => n14076);
   U4512 : OAI22_X1 port map( A1 => n60876, A2 => n61965, B1 => n4599, B2 => 
                           n60875, ZN => n14021);
   U4513 : OAI22_X1 port map( A1 => n60876, A2 => n61979, B1 => n4598, B2 => 
                           n60875, ZN => n14022);
   U4514 : OAI22_X1 port map( A1 => n60876, A2 => n61993, B1 => n4597, B2 => 
                           n60875, ZN => n14023);
   U4515 : OAI22_X1 port map( A1 => n60876, A2 => n62007, B1 => n4596, B2 => 
                           n60875, ZN => n14024);
   U4516 : OAI22_X1 port map( A1 => n60876, A2 => n62021, B1 => n4595, B2 => 
                           n60875, ZN => n14025);
   U4517 : OAI22_X1 port map( A1 => n60877, A2 => n62035, B1 => n4594, B2 => 
                           n60875, ZN => n14026);
   U4518 : OAI22_X1 port map( A1 => n60877, A2 => n62049, B1 => n4593, B2 => 
                           n60875, ZN => n14027);
   U4519 : OAI22_X1 port map( A1 => n60877, A2 => n62063, B1 => n4592, B2 => 
                           n60875, ZN => n14028);
   U4520 : OAI22_X1 port map( A1 => n60877, A2 => n62077, B1 => n4591, B2 => 
                           n60875, ZN => n14029);
   U4521 : OAI22_X1 port map( A1 => n60877, A2 => n62091, B1 => n4590, B2 => 
                           n60875, ZN => n14030);
   U4522 : OAI22_X1 port map( A1 => n60878, A2 => n62105, B1 => n4589, B2 => 
                           n60875, ZN => n14031);
   U4523 : OAI22_X1 port map( A1 => n60878, A2 => n60958, B1 => n4588, B2 => 
                           n60875, ZN => n14032);
   U4524 : OAI22_X1 port map( A1 => n60878, A2 => n60972, B1 => n4587, B2 => 
                           n15112, ZN => n14033);
   U4525 : OAI22_X1 port map( A1 => n60878, A2 => n60986, B1 => n4586, B2 => 
                           n15112, ZN => n14034);
   U4526 : OAI22_X1 port map( A1 => n60878, A2 => n61000, B1 => n4585, B2 => 
                           n15112, ZN => n14035);
   U4527 : OAI22_X1 port map( A1 => n60879, A2 => n61014, B1 => n4584, B2 => 
                           n15112, ZN => n14036);
   U4528 : OAI22_X1 port map( A1 => n60879, A2 => n61028, B1 => n4583, B2 => 
                           n15112, ZN => n14037);
   U4529 : OAI22_X1 port map( A1 => n60879, A2 => n61042, B1 => n4582, B2 => 
                           n15112, ZN => n14038);
   U4530 : OAI22_X1 port map( A1 => n60879, A2 => n61056, B1 => n4581, B2 => 
                           n15112, ZN => n14039);
   U4531 : OAI22_X1 port map( A1 => n60879, A2 => n61070, B1 => n4580, B2 => 
                           n60875, ZN => n14040);
   U4532 : OAI22_X1 port map( A1 => n60880, A2 => n61084, B1 => n4579, B2 => 
                           n60875, ZN => n14041);
   U4533 : OAI22_X1 port map( A1 => n60880, A2 => n61098, B1 => n4578, B2 => 
                           n60875, ZN => n14042);
   U4534 : OAI22_X1 port map( A1 => n60880, A2 => n61112, B1 => n4577, B2 => 
                           n60875, ZN => n14043);
   U4535 : OAI22_X1 port map( A1 => n60880, A2 => n61126, B1 => n4576, B2 => 
                           n60875, ZN => n14044);
   U4536 : OAI22_X1 port map( A1 => n60849, A2 => n61966, B1 => n4551, B2 => 
                           n60848, ZN => n13925);
   U4537 : OAI22_X1 port map( A1 => n60849, A2 => n61980, B1 => n4550, B2 => 
                           n60848, ZN => n13926);
   U4538 : OAI22_X1 port map( A1 => n60849, A2 => n61994, B1 => n4549, B2 => 
                           n60848, ZN => n13927);
   U4539 : OAI22_X1 port map( A1 => n60849, A2 => n62008, B1 => n4548, B2 => 
                           n60848, ZN => n13928);
   U4540 : OAI22_X1 port map( A1 => n60849, A2 => n62022, B1 => n4547, B2 => 
                           n60848, ZN => n13929);
   U4541 : OAI22_X1 port map( A1 => n60850, A2 => n62036, B1 => n4546, B2 => 
                           n60848, ZN => n13930);
   U4542 : OAI22_X1 port map( A1 => n60850, A2 => n62050, B1 => n4545, B2 => 
                           n60848, ZN => n13931);
   U4543 : OAI22_X1 port map( A1 => n60850, A2 => n62064, B1 => n4544, B2 => 
                           n60848, ZN => n13932);
   U4544 : OAI22_X1 port map( A1 => n60850, A2 => n62078, B1 => n4543, B2 => 
                           n60848, ZN => n13933);
   U4545 : OAI22_X1 port map( A1 => n60850, A2 => n62092, B1 => n4542, B2 => 
                           n60848, ZN => n13934);
   U4546 : OAI22_X1 port map( A1 => n60851, A2 => n62106, B1 => n4541, B2 => 
                           n60848, ZN => n13935);
   U4547 : OAI22_X1 port map( A1 => n60851, A2 => n60959, B1 => n4540, B2 => 
                           n60848, ZN => n13936);
   U4548 : OAI22_X1 port map( A1 => n60851, A2 => n60973, B1 => n4539, B2 => 
                           n15118, ZN => n13937);
   U4549 : OAI22_X1 port map( A1 => n60851, A2 => n60987, B1 => n4538, B2 => 
                           n15118, ZN => n13938);
   U4550 : OAI22_X1 port map( A1 => n60851, A2 => n61001, B1 => n4537, B2 => 
                           n15118, ZN => n13939);
   U4551 : OAI22_X1 port map( A1 => n60852, A2 => n61015, B1 => n4536, B2 => 
                           n15118, ZN => n13940);
   U4552 : OAI22_X1 port map( A1 => n60852, A2 => n61029, B1 => n4535, B2 => 
                           n15118, ZN => n13941);
   U4553 : OAI22_X1 port map( A1 => n60852, A2 => n61043, B1 => n4534, B2 => 
                           n15118, ZN => n13942);
   U4554 : OAI22_X1 port map( A1 => n60852, A2 => n61057, B1 => n4533, B2 => 
                           n15118, ZN => n13943);
   U4555 : OAI22_X1 port map( A1 => n60852, A2 => n61071, B1 => n4532, B2 => 
                           n60848, ZN => n13944);
   U4556 : OAI22_X1 port map( A1 => n60853, A2 => n61085, B1 => n4531, B2 => 
                           n60848, ZN => n13945);
   U4557 : OAI22_X1 port map( A1 => n60853, A2 => n61099, B1 => n4530, B2 => 
                           n60848, ZN => n13946);
   U4558 : OAI22_X1 port map( A1 => n60853, A2 => n61113, B1 => n4529, B2 => 
                           n60848, ZN => n13947);
   U4559 : OAI22_X1 port map( A1 => n60853, A2 => n61127, B1 => n4528, B2 => 
                           n60848, ZN => n13948);
   U4560 : OAI22_X1 port map( A1 => n60840, A2 => n61966, B1 => n4527, B2 => 
                           n60839, ZN => n13893);
   U4561 : OAI22_X1 port map( A1 => n60840, A2 => n61980, B1 => n4526, B2 => 
                           n60839, ZN => n13894);
   U4562 : OAI22_X1 port map( A1 => n60840, A2 => n61994, B1 => n4525, B2 => 
                           n60839, ZN => n13895);
   U4563 : OAI22_X1 port map( A1 => n60840, A2 => n62008, B1 => n4524, B2 => 
                           n60839, ZN => n13896);
   U4564 : OAI22_X1 port map( A1 => n60840, A2 => n62022, B1 => n4523, B2 => 
                           n60839, ZN => n13897);
   U4565 : OAI22_X1 port map( A1 => n60841, A2 => n62036, B1 => n4522, B2 => 
                           n60839, ZN => n13898);
   U4566 : OAI22_X1 port map( A1 => n60841, A2 => n62050, B1 => n4521, B2 => 
                           n60839, ZN => n13899);
   U4567 : OAI22_X1 port map( A1 => n60841, A2 => n62064, B1 => n4520, B2 => 
                           n60839, ZN => n13900);
   U4568 : OAI22_X1 port map( A1 => n60841, A2 => n62078, B1 => n4519, B2 => 
                           n60839, ZN => n13901);
   U4569 : OAI22_X1 port map( A1 => n60841, A2 => n62092, B1 => n4518, B2 => 
                           n60839, ZN => n13902);
   U4570 : OAI22_X1 port map( A1 => n60842, A2 => n62106, B1 => n4517, B2 => 
                           n60839, ZN => n13903);
   U4571 : OAI22_X1 port map( A1 => n60842, A2 => n60959, B1 => n4516, B2 => 
                           n60839, ZN => n13904);
   U4572 : OAI22_X1 port map( A1 => n60842, A2 => n60973, B1 => n4515, B2 => 
                           n15120, ZN => n13905);
   U4573 : OAI22_X1 port map( A1 => n60842, A2 => n60987, B1 => n4514, B2 => 
                           n15120, ZN => n13906);
   U4574 : OAI22_X1 port map( A1 => n60842, A2 => n61001, B1 => n4513, B2 => 
                           n15120, ZN => n13907);
   U4575 : OAI22_X1 port map( A1 => n60843, A2 => n61015, B1 => n4512, B2 => 
                           n15120, ZN => n13908);
   U4576 : OAI22_X1 port map( A1 => n60843, A2 => n61029, B1 => n4511, B2 => 
                           n15120, ZN => n13909);
   U4577 : OAI22_X1 port map( A1 => n60843, A2 => n61043, B1 => n4510, B2 => 
                           n15120, ZN => n13910);
   U4578 : OAI22_X1 port map( A1 => n60843, A2 => n61057, B1 => n4509, B2 => 
                           n15120, ZN => n13911);
   U4579 : OAI22_X1 port map( A1 => n60843, A2 => n61071, B1 => n4508, B2 => 
                           n60839, ZN => n13912);
   U4580 : OAI22_X1 port map( A1 => n60844, A2 => n61085, B1 => n4507, B2 => 
                           n60839, ZN => n13913);
   U4581 : OAI22_X1 port map( A1 => n60844, A2 => n61099, B1 => n4506, B2 => 
                           n60839, ZN => n13914);
   U4582 : OAI22_X1 port map( A1 => n60844, A2 => n61113, B1 => n4505, B2 => 
                           n60839, ZN => n13915);
   U4583 : OAI22_X1 port map( A1 => n60844, A2 => n61127, B1 => n4504, B2 => 
                           n60839, ZN => n13916);
   U4584 : OAI22_X1 port map( A1 => n60102, A2 => n61972, B1 => n4407, B2 => 
                           n60101, ZN => n11269);
   U4585 : OAI22_X1 port map( A1 => n60102, A2 => n61986, B1 => n4406, B2 => 
                           n60101, ZN => n11270);
   U4586 : OAI22_X1 port map( A1 => n60102, A2 => n62000, B1 => n4405, B2 => 
                           n60101, ZN => n11271);
   U4587 : OAI22_X1 port map( A1 => n60102, A2 => n62014, B1 => n4404, B2 => 
                           n60101, ZN => n11272);
   U4588 : OAI22_X1 port map( A1 => n60102, A2 => n62028, B1 => n4403, B2 => 
                           n60101, ZN => n11273);
   U4589 : OAI22_X1 port map( A1 => n60093, A2 => n61973, B1 => n3918, B2 => 
                           n60092, ZN => n11237);
   U4590 : OAI22_X1 port map( A1 => n60093, A2 => n61987, B1 => n3917, B2 => 
                           n60092, ZN => n11238);
   U4591 : OAI22_X1 port map( A1 => n60093, A2 => n62001, B1 => n3916, B2 => 
                           n60092, ZN => n11239);
   U4592 : OAI22_X1 port map( A1 => n60093, A2 => n62015, B1 => n3915, B2 => 
                           n60092, ZN => n11240);
   U4593 : OAI22_X1 port map( A1 => n60093, A2 => n62029, B1 => n3914, B2 => 
                           n60092, ZN => n11241);
   U4594 : OAI22_X1 port map( A1 => n60094, A2 => n62043, B1 => n3913, B2 => 
                           n60092, ZN => n11242);
   U4595 : OAI22_X1 port map( A1 => n60094, A2 => n62057, B1 => n3912, B2 => 
                           n60092, ZN => n11243);
   U4596 : OAI22_X1 port map( A1 => n60094, A2 => n62071, B1 => n3911, B2 => 
                           n60092, ZN => n11244);
   U4597 : OAI22_X1 port map( A1 => n60094, A2 => n62085, B1 => n3910, B2 => 
                           n60092, ZN => n11245);
   U4598 : OAI22_X1 port map( A1 => n60094, A2 => n62099, B1 => n3909, B2 => 
                           n60092, ZN => n11246);
   U4599 : OAI22_X1 port map( A1 => n60095, A2 => n62113, B1 => n3908, B2 => 
                           n60092, ZN => n11247);
   U4600 : OAI22_X1 port map( A1 => n60095, A2 => n60966, B1 => n3907, B2 => 
                           n60092, ZN => n11248);
   U4601 : OAI22_X1 port map( A1 => n60095, A2 => n60980, B1 => n3906, B2 => 
                           n15229, ZN => n11249);
   U4602 : OAI22_X1 port map( A1 => n60095, A2 => n60994, B1 => n3905, B2 => 
                           n15229, ZN => n11250);
   U4603 : OAI22_X1 port map( A1 => n60095, A2 => n61008, B1 => n3904, B2 => 
                           n15229, ZN => n11251);
   U4604 : OAI22_X1 port map( A1 => n60096, A2 => n61022, B1 => n3903, B2 => 
                           n15229, ZN => n11252);
   U4605 : OAI22_X1 port map( A1 => n60096, A2 => n61036, B1 => n3902, B2 => 
                           n15229, ZN => n11253);
   U4606 : OAI22_X1 port map( A1 => n60096, A2 => n61050, B1 => n3901, B2 => 
                           n15229, ZN => n11254);
   U4607 : OAI22_X1 port map( A1 => n60096, A2 => n61064, B1 => n3900, B2 => 
                           n15229, ZN => n11255);
   U4608 : OAI22_X1 port map( A1 => n60096, A2 => n61078, B1 => n3899, B2 => 
                           n60092, ZN => n11256);
   U4609 : OAI22_X1 port map( A1 => n60097, A2 => n61092, B1 => n3898, B2 => 
                           n60092, ZN => n11257);
   U4610 : OAI22_X1 port map( A1 => n60097, A2 => n61106, B1 => n3897, B2 => 
                           n60092, ZN => n11258);
   U4611 : OAI22_X1 port map( A1 => n60097, A2 => n61120, B1 => n3896, B2 => 
                           n60092, ZN => n11259);
   U4612 : OAI22_X1 port map( A1 => n60097, A2 => n61134, B1 => n3895, B2 => 
                           n60092, ZN => n11260);
   U4613 : OAI22_X1 port map( A1 => n60084, A2 => n61973, B1 => n3894, B2 => 
                           n60083, ZN => n11205);
   U4614 : OAI22_X1 port map( A1 => n60084, A2 => n61987, B1 => n3893, B2 => 
                           n60083, ZN => n11206);
   U4615 : OAI22_X1 port map( A1 => n60084, A2 => n62001, B1 => n3892, B2 => 
                           n60083, ZN => n11207);
   U4616 : OAI22_X1 port map( A1 => n60084, A2 => n62015, B1 => n3891, B2 => 
                           n60083, ZN => n11208);
   U4617 : OAI22_X1 port map( A1 => n60084, A2 => n62029, B1 => n3890, B2 => 
                           n60083, ZN => n11209);
   U4618 : OAI22_X1 port map( A1 => n60085, A2 => n62043, B1 => n3889, B2 => 
                           n60083, ZN => n11210);
   U4619 : OAI22_X1 port map( A1 => n60085, A2 => n62057, B1 => n3888, B2 => 
                           n60083, ZN => n11211);
   U4620 : OAI22_X1 port map( A1 => n60085, A2 => n62071, B1 => n3887, B2 => 
                           n60083, ZN => n11212);
   U4621 : OAI22_X1 port map( A1 => n60085, A2 => n62085, B1 => n3886, B2 => 
                           n60083, ZN => n11213);
   U4622 : OAI22_X1 port map( A1 => n60085, A2 => n62099, B1 => n3885, B2 => 
                           n60083, ZN => n11214);
   U4623 : OAI22_X1 port map( A1 => n60086, A2 => n62113, B1 => n3884, B2 => 
                           n60083, ZN => n11215);
   U4624 : OAI22_X1 port map( A1 => n60086, A2 => n60966, B1 => n3883, B2 => 
                           n60083, ZN => n11216);
   U4625 : OAI22_X1 port map( A1 => n60086, A2 => n60980, B1 => n3882, B2 => 
                           n15231, ZN => n11217);
   U4626 : OAI22_X1 port map( A1 => n60086, A2 => n60994, B1 => n3881, B2 => 
                           n15231, ZN => n11218);
   U4627 : OAI22_X1 port map( A1 => n60086, A2 => n61008, B1 => n3880, B2 => 
                           n15231, ZN => n11219);
   U4628 : OAI22_X1 port map( A1 => n60087, A2 => n61022, B1 => n3879, B2 => 
                           n15231, ZN => n11220);
   U4629 : OAI22_X1 port map( A1 => n60087, A2 => n61036, B1 => n3878, B2 => 
                           n15231, ZN => n11221);
   U4630 : OAI22_X1 port map( A1 => n60087, A2 => n61050, B1 => n3877, B2 => 
                           n15231, ZN => n11222);
   U4631 : OAI22_X1 port map( A1 => n60087, A2 => n61064, B1 => n3876, B2 => 
                           n15231, ZN => n11223);
   U4632 : OAI22_X1 port map( A1 => n60087, A2 => n61078, B1 => n3875, B2 => 
                           n60083, ZN => n11224);
   U4633 : OAI22_X1 port map( A1 => n60088, A2 => n61092, B1 => n3874, B2 => 
                           n60083, ZN => n11225);
   U4634 : OAI22_X1 port map( A1 => n60088, A2 => n61106, B1 => n3873, B2 => 
                           n60083, ZN => n11226);
   U4635 : OAI22_X1 port map( A1 => n60088, A2 => n61120, B1 => n3872, B2 => 
                           n60083, ZN => n11227);
   U4636 : OAI22_X1 port map( A1 => n60088, A2 => n61134, B1 => n3871, B2 => 
                           n60083, ZN => n11228);
   U4637 : OAI22_X1 port map( A1 => n60075, A2 => n61973, B1 => n3870, B2 => 
                           n60074, ZN => n11173);
   U4638 : OAI22_X1 port map( A1 => n60075, A2 => n61987, B1 => n3869, B2 => 
                           n60074, ZN => n11174);
   U4639 : OAI22_X1 port map( A1 => n60075, A2 => n62001, B1 => n3868, B2 => 
                           n60074, ZN => n11175);
   U4640 : OAI22_X1 port map( A1 => n60075, A2 => n62015, B1 => n3867, B2 => 
                           n60074, ZN => n11176);
   U4641 : OAI22_X1 port map( A1 => n60075, A2 => n62029, B1 => n3866, B2 => 
                           n60074, ZN => n11177);
   U4642 : OAI22_X1 port map( A1 => n60076, A2 => n62043, B1 => n3865, B2 => 
                           n60074, ZN => n11178);
   U4643 : OAI22_X1 port map( A1 => n60076, A2 => n62057, B1 => n3864, B2 => 
                           n60074, ZN => n11179);
   U4644 : OAI22_X1 port map( A1 => n60076, A2 => n62071, B1 => n3863, B2 => 
                           n60074, ZN => n11180);
   U4645 : OAI22_X1 port map( A1 => n60076, A2 => n62085, B1 => n3862, B2 => 
                           n60074, ZN => n11181);
   U4646 : OAI22_X1 port map( A1 => n60076, A2 => n62099, B1 => n3861, B2 => 
                           n60074, ZN => n11182);
   U4647 : OAI22_X1 port map( A1 => n60077, A2 => n62113, B1 => n3860, B2 => 
                           n60074, ZN => n11183);
   U4648 : OAI22_X1 port map( A1 => n60077, A2 => n60966, B1 => n3859, B2 => 
                           n60074, ZN => n11184);
   U4649 : OAI22_X1 port map( A1 => n60077, A2 => n60980, B1 => n3858, B2 => 
                           n15232, ZN => n11185);
   U4650 : OAI22_X1 port map( A1 => n60077, A2 => n60994, B1 => n3857, B2 => 
                           n15232, ZN => n11186);
   U4651 : OAI22_X1 port map( A1 => n60077, A2 => n61008, B1 => n3856, B2 => 
                           n15232, ZN => n11187);
   U4652 : OAI22_X1 port map( A1 => n60078, A2 => n61022, B1 => n3855, B2 => 
                           n15232, ZN => n11188);
   U4653 : OAI22_X1 port map( A1 => n60078, A2 => n61036, B1 => n3854, B2 => 
                           n15232, ZN => n11189);
   U4654 : OAI22_X1 port map( A1 => n60078, A2 => n61050, B1 => n3853, B2 => 
                           n15232, ZN => n11190);
   U4655 : OAI22_X1 port map( A1 => n60078, A2 => n61064, B1 => n3852, B2 => 
                           n15232, ZN => n11191);
   U4656 : OAI22_X1 port map( A1 => n60078, A2 => n61078, B1 => n3851, B2 => 
                           n60074, ZN => n11192);
   U4657 : OAI22_X1 port map( A1 => n60079, A2 => n61092, B1 => n3850, B2 => 
                           n60074, ZN => n11193);
   U4658 : OAI22_X1 port map( A1 => n60079, A2 => n61106, B1 => n3849, B2 => 
                           n60074, ZN => n11194);
   U4659 : OAI22_X1 port map( A1 => n60079, A2 => n61120, B1 => n3848, B2 => 
                           n60074, ZN => n11195);
   U4660 : OAI22_X1 port map( A1 => n60079, A2 => n61134, B1 => n3847, B2 => 
                           n60074, ZN => n11196);
   U4661 : OAI22_X1 port map( A1 => n60057, A2 => n61973, B1 => n3822, B2 => 
                           n60056, ZN => n11109);
   U4662 : OAI22_X1 port map( A1 => n60057, A2 => n61987, B1 => n3821, B2 => 
                           n60056, ZN => n11110);
   U4663 : OAI22_X1 port map( A1 => n60057, A2 => n62001, B1 => n3820, B2 => 
                           n60056, ZN => n11111);
   U4664 : OAI22_X1 port map( A1 => n60057, A2 => n62015, B1 => n3819, B2 => 
                           n60056, ZN => n11112);
   U4665 : OAI22_X1 port map( A1 => n60057, A2 => n62029, B1 => n3818, B2 => 
                           n60056, ZN => n11113);
   U4666 : OAI22_X1 port map( A1 => n60058, A2 => n62043, B1 => n3817, B2 => 
                           n60056, ZN => n11114);
   U4667 : OAI22_X1 port map( A1 => n60058, A2 => n62057, B1 => n3816, B2 => 
                           n60056, ZN => n11115);
   U4668 : OAI22_X1 port map( A1 => n60058, A2 => n62071, B1 => n3815, B2 => 
                           n60056, ZN => n11116);
   U4669 : OAI22_X1 port map( A1 => n60058, A2 => n62085, B1 => n3814, B2 => 
                           n60056, ZN => n11117);
   U4670 : OAI22_X1 port map( A1 => n60058, A2 => n62099, B1 => n3813, B2 => 
                           n60056, ZN => n11118);
   U4671 : OAI22_X1 port map( A1 => n60059, A2 => n62113, B1 => n3812, B2 => 
                           n60056, ZN => n11119);
   U4672 : OAI22_X1 port map( A1 => n60059, A2 => n60966, B1 => n3811, B2 => 
                           n60056, ZN => n11120);
   U4673 : OAI22_X1 port map( A1 => n60059, A2 => n60980, B1 => n3810, B2 => 
                           n15234, ZN => n11121);
   U4674 : OAI22_X1 port map( A1 => n60059, A2 => n60994, B1 => n3809, B2 => 
                           n15234, ZN => n11122);
   U4675 : OAI22_X1 port map( A1 => n60059, A2 => n61008, B1 => n3808, B2 => 
                           n15234, ZN => n11123);
   U4676 : OAI22_X1 port map( A1 => n60060, A2 => n61022, B1 => n3807, B2 => 
                           n15234, ZN => n11124);
   U4677 : OAI22_X1 port map( A1 => n60060, A2 => n61036, B1 => n3806, B2 => 
                           n15234, ZN => n11125);
   U4678 : OAI22_X1 port map( A1 => n60060, A2 => n61050, B1 => n3805, B2 => 
                           n15234, ZN => n11126);
   U4679 : OAI22_X1 port map( A1 => n60060, A2 => n61064, B1 => n3804, B2 => 
                           n15234, ZN => n11127);
   U4680 : OAI22_X1 port map( A1 => n60060, A2 => n61078, B1 => n3803, B2 => 
                           n60056, ZN => n11128);
   U4681 : OAI22_X1 port map( A1 => n60061, A2 => n61092, B1 => n3802, B2 => 
                           n60056, ZN => n11129);
   U4682 : OAI22_X1 port map( A1 => n60061, A2 => n61106, B1 => n3801, B2 => 
                           n60056, ZN => n11130);
   U4683 : OAI22_X1 port map( A1 => n60061, A2 => n61120, B1 => n3800, B2 => 
                           n60056, ZN => n11131);
   U4684 : OAI22_X1 port map( A1 => n60061, A2 => n61134, B1 => n3799, B2 => 
                           n60056, ZN => n11132);
   U4685 : OAI22_X1 port map( A1 => n60021, A2 => n61973, B1 => n3726, B2 => 
                           n60020, ZN => n10981);
   U4686 : OAI22_X1 port map( A1 => n60021, A2 => n61987, B1 => n3725, B2 => 
                           n60020, ZN => n10982);
   U4687 : OAI22_X1 port map( A1 => n60021, A2 => n62001, B1 => n3724, B2 => 
                           n60020, ZN => n10983);
   U4688 : OAI22_X1 port map( A1 => n60021, A2 => n62015, B1 => n3723, B2 => 
                           n60020, ZN => n10984);
   U4689 : OAI22_X1 port map( A1 => n60021, A2 => n62029, B1 => n3722, B2 => 
                           n60020, ZN => n10985);
   U4690 : OAI22_X1 port map( A1 => n60022, A2 => n62043, B1 => n3721, B2 => 
                           n60020, ZN => n10986);
   U4691 : OAI22_X1 port map( A1 => n60022, A2 => n62057, B1 => n3720, B2 => 
                           n60020, ZN => n10987);
   U4692 : OAI22_X1 port map( A1 => n60022, A2 => n62071, B1 => n3719, B2 => 
                           n60020, ZN => n10988);
   U4693 : OAI22_X1 port map( A1 => n60022, A2 => n62085, B1 => n3718, B2 => 
                           n60020, ZN => n10989);
   U4694 : OAI22_X1 port map( A1 => n60022, A2 => n62099, B1 => n3717, B2 => 
                           n60020, ZN => n10990);
   U4695 : OAI22_X1 port map( A1 => n60023, A2 => n62113, B1 => n3716, B2 => 
                           n60020, ZN => n10991);
   U4696 : OAI22_X1 port map( A1 => n60023, A2 => n60966, B1 => n3715, B2 => 
                           n60020, ZN => n10992);
   U4697 : OAI22_X1 port map( A1 => n60023, A2 => n60980, B1 => n3714, B2 => 
                           n15238, ZN => n10993);
   U4698 : OAI22_X1 port map( A1 => n60023, A2 => n60994, B1 => n3713, B2 => 
                           n15238, ZN => n10994);
   U4699 : OAI22_X1 port map( A1 => n60023, A2 => n61008, B1 => n3712, B2 => 
                           n15238, ZN => n10995);
   U4700 : OAI22_X1 port map( A1 => n60024, A2 => n61022, B1 => n3711, B2 => 
                           n15238, ZN => n10996);
   U4701 : OAI22_X1 port map( A1 => n60024, A2 => n61036, B1 => n3710, B2 => 
                           n15238, ZN => n10997);
   U4702 : OAI22_X1 port map( A1 => n60024, A2 => n61050, B1 => n3709, B2 => 
                           n15238, ZN => n10998);
   U4703 : OAI22_X1 port map( A1 => n60024, A2 => n61064, B1 => n3708, B2 => 
                           n15238, ZN => n10999);
   U4704 : OAI22_X1 port map( A1 => n60024, A2 => n61078, B1 => n3707, B2 => 
                           n60020, ZN => n11000);
   U4705 : OAI22_X1 port map( A1 => n60025, A2 => n61092, B1 => n3706, B2 => 
                           n60020, ZN => n11001);
   U4706 : OAI22_X1 port map( A1 => n60025, A2 => n61106, B1 => n3705, B2 => 
                           n60020, ZN => n11002);
   U4707 : OAI22_X1 port map( A1 => n60025, A2 => n61120, B1 => n3704, B2 => 
                           n60020, ZN => n11003);
   U4708 : OAI22_X1 port map( A1 => n60025, A2 => n61134, B1 => n3703, B2 => 
                           n60020, ZN => n11004);
   U4709 : OAI22_X1 port map( A1 => n60012, A2 => n61973, B1 => n3702, B2 => 
                           n60011, ZN => n10949);
   U4710 : OAI22_X1 port map( A1 => n60012, A2 => n61987, B1 => n3701, B2 => 
                           n60011, ZN => n10950);
   U4711 : OAI22_X1 port map( A1 => n60012, A2 => n62001, B1 => n3700, B2 => 
                           n60011, ZN => n10951);
   U4712 : OAI22_X1 port map( A1 => n60012, A2 => n62015, B1 => n3699, B2 => 
                           n60011, ZN => n10952);
   U4713 : OAI22_X1 port map( A1 => n60012, A2 => n62029, B1 => n3698, B2 => 
                           n60011, ZN => n10953);
   U4714 : OAI22_X1 port map( A1 => n60013, A2 => n62043, B1 => n3697, B2 => 
                           n60011, ZN => n10954);
   U4715 : OAI22_X1 port map( A1 => n60013, A2 => n62057, B1 => n3696, B2 => 
                           n60011, ZN => n10955);
   U4716 : OAI22_X1 port map( A1 => n60013, A2 => n62071, B1 => n3695, B2 => 
                           n60011, ZN => n10956);
   U4717 : OAI22_X1 port map( A1 => n60013, A2 => n62085, B1 => n3694, B2 => 
                           n60011, ZN => n10957);
   U4718 : OAI22_X1 port map( A1 => n60013, A2 => n62099, B1 => n3693, B2 => 
                           n60011, ZN => n10958);
   U4719 : OAI22_X1 port map( A1 => n60014, A2 => n62113, B1 => n3692, B2 => 
                           n60011, ZN => n10959);
   U4720 : OAI22_X1 port map( A1 => n60014, A2 => n60966, B1 => n3691, B2 => 
                           n60011, ZN => n10960);
   U4721 : OAI22_X1 port map( A1 => n60014, A2 => n60980, B1 => n3690, B2 => 
                           n15239, ZN => n10961);
   U4722 : OAI22_X1 port map( A1 => n60014, A2 => n60994, B1 => n3689, B2 => 
                           n15239, ZN => n10962);
   U4723 : OAI22_X1 port map( A1 => n60014, A2 => n61008, B1 => n3688, B2 => 
                           n15239, ZN => n10963);
   U4724 : OAI22_X1 port map( A1 => n60015, A2 => n61022, B1 => n3687, B2 => 
                           n15239, ZN => n10964);
   U4725 : OAI22_X1 port map( A1 => n60015, A2 => n61036, B1 => n3686, B2 => 
                           n15239, ZN => n10965);
   U4726 : OAI22_X1 port map( A1 => n60015, A2 => n61050, B1 => n3685, B2 => 
                           n15239, ZN => n10966);
   U4727 : OAI22_X1 port map( A1 => n60015, A2 => n61064, B1 => n3684, B2 => 
                           n15239, ZN => n10967);
   U4728 : OAI22_X1 port map( A1 => n60015, A2 => n61078, B1 => n3683, B2 => 
                           n60011, ZN => n10968);
   U4729 : OAI22_X1 port map( A1 => n60016, A2 => n61092, B1 => n3682, B2 => 
                           n60011, ZN => n10969);
   U4730 : OAI22_X1 port map( A1 => n60016, A2 => n61106, B1 => n3681, B2 => 
                           n60011, ZN => n10970);
   U4731 : OAI22_X1 port map( A1 => n60016, A2 => n61120, B1 => n3680, B2 => 
                           n60011, ZN => n10971);
   U4732 : OAI22_X1 port map( A1 => n60016, A2 => n61134, B1 => n3679, B2 => 
                           n60011, ZN => n10972);
   U4733 : OAI22_X1 port map( A1 => n59949, A2 => n61974, B1 => n3596, B2 => 
                           n59948, ZN => n10725);
   U4734 : OAI22_X1 port map( A1 => n59949, A2 => n61988, B1 => n3595, B2 => 
                           n59948, ZN => n10726);
   U4735 : OAI22_X1 port map( A1 => n59949, A2 => n62002, B1 => n3594, B2 => 
                           n59948, ZN => n10727);
   U4736 : OAI22_X1 port map( A1 => n59949, A2 => n62016, B1 => n3593, B2 => 
                           n59948, ZN => n10728);
   U4737 : OAI22_X1 port map( A1 => n59949, A2 => n62030, B1 => n3592, B2 => 
                           n59948, ZN => n10729);
   U4738 : OAI22_X1 port map( A1 => n59950, A2 => n62044, B1 => n3591, B2 => 
                           n59948, ZN => n10730);
   U4739 : OAI22_X1 port map( A1 => n59950, A2 => n62058, B1 => n3590, B2 => 
                           n59948, ZN => n10731);
   U4740 : OAI22_X1 port map( A1 => n59950, A2 => n62072, B1 => n3589, B2 => 
                           n59948, ZN => n10732);
   U4741 : OAI22_X1 port map( A1 => n59950, A2 => n62086, B1 => n3588, B2 => 
                           n59948, ZN => n10733);
   U4742 : OAI22_X1 port map( A1 => n59950, A2 => n62100, B1 => n3587, B2 => 
                           n59948, ZN => n10734);
   U4743 : OAI22_X1 port map( A1 => n59951, A2 => n62114, B1 => n3586, B2 => 
                           n59948, ZN => n10735);
   U4744 : OAI22_X1 port map( A1 => n59951, A2 => n60967, B1 => n3585, B2 => 
                           n59948, ZN => n10736);
   U4745 : OAI22_X1 port map( A1 => n59951, A2 => n60981, B1 => n3584, B2 => 
                           n15246, ZN => n10737);
   U4746 : OAI22_X1 port map( A1 => n59951, A2 => n60995, B1 => n3583, B2 => 
                           n15246, ZN => n10738);
   U4747 : OAI22_X1 port map( A1 => n59951, A2 => n61009, B1 => n3582, B2 => 
                           n15246, ZN => n10739);
   U4748 : OAI22_X1 port map( A1 => n59952, A2 => n61023, B1 => n3581, B2 => 
                           n15246, ZN => n10740);
   U4749 : OAI22_X1 port map( A1 => n59952, A2 => n61037, B1 => n3580, B2 => 
                           n15246, ZN => n10741);
   U4750 : OAI22_X1 port map( A1 => n59952, A2 => n61051, B1 => n3579, B2 => 
                           n15246, ZN => n10742);
   U4751 : OAI22_X1 port map( A1 => n59952, A2 => n61065, B1 => n3578, B2 => 
                           n15246, ZN => n10743);
   U4752 : OAI22_X1 port map( A1 => n59952, A2 => n61079, B1 => n3577, B2 => 
                           n59948, ZN => n10744);
   U4753 : OAI22_X1 port map( A1 => n59953, A2 => n61093, B1 => n3576, B2 => 
                           n59948, ZN => n10745);
   U4754 : OAI22_X1 port map( A1 => n59953, A2 => n61107, B1 => n3575, B2 => 
                           n59948, ZN => n10746);
   U4755 : OAI22_X1 port map( A1 => n59953, A2 => n61121, B1 => n3574, B2 => 
                           n59948, ZN => n10747);
   U4756 : OAI22_X1 port map( A1 => n59953, A2 => n61135, B1 => n3573, B2 => 
                           n59948, ZN => n10748);
   U4757 : OAI22_X1 port map( A1 => n59940, A2 => n61974, B1 => n3572, B2 => 
                           n59939, ZN => n10693);
   U4758 : OAI22_X1 port map( A1 => n59940, A2 => n61988, B1 => n3571, B2 => 
                           n59939, ZN => n10694);
   U4759 : OAI22_X1 port map( A1 => n59940, A2 => n62002, B1 => n3570, B2 => 
                           n59939, ZN => n10695);
   U4760 : OAI22_X1 port map( A1 => n59940, A2 => n62016, B1 => n3569, B2 => 
                           n59939, ZN => n10696);
   U4761 : OAI22_X1 port map( A1 => n59940, A2 => n62030, B1 => n3568, B2 => 
                           n59939, ZN => n10697);
   U4762 : OAI22_X1 port map( A1 => n59941, A2 => n62044, B1 => n3567, B2 => 
                           n59939, ZN => n10698);
   U4763 : OAI22_X1 port map( A1 => n59941, A2 => n62058, B1 => n3566, B2 => 
                           n59939, ZN => n10699);
   U4764 : OAI22_X1 port map( A1 => n59941, A2 => n62072, B1 => n3565, B2 => 
                           n59939, ZN => n10700);
   U4765 : OAI22_X1 port map( A1 => n59941, A2 => n62086, B1 => n3564, B2 => 
                           n59939, ZN => n10701);
   U4766 : OAI22_X1 port map( A1 => n59941, A2 => n62100, B1 => n3563, B2 => 
                           n59939, ZN => n10702);
   U4767 : OAI22_X1 port map( A1 => n59942, A2 => n62114, B1 => n3562, B2 => 
                           n59939, ZN => n10703);
   U4768 : OAI22_X1 port map( A1 => n59942, A2 => n60967, B1 => n3561, B2 => 
                           n59939, ZN => n10704);
   U4769 : OAI22_X1 port map( A1 => n59942, A2 => n60981, B1 => n3560, B2 => 
                           n15248, ZN => n10705);
   U4770 : OAI22_X1 port map( A1 => n59942, A2 => n60995, B1 => n3559, B2 => 
                           n15248, ZN => n10706);
   U4771 : OAI22_X1 port map( A1 => n59942, A2 => n61009, B1 => n3558, B2 => 
                           n15248, ZN => n10707);
   U4772 : OAI22_X1 port map( A1 => n59943, A2 => n61023, B1 => n3557, B2 => 
                           n15248, ZN => n10708);
   U4773 : OAI22_X1 port map( A1 => n59943, A2 => n61037, B1 => n3556, B2 => 
                           n15248, ZN => n10709);
   U4774 : OAI22_X1 port map( A1 => n59943, A2 => n61051, B1 => n3555, B2 => 
                           n15248, ZN => n10710);
   U4775 : OAI22_X1 port map( A1 => n59943, A2 => n61065, B1 => n3554, B2 => 
                           n15248, ZN => n10711);
   U4776 : OAI22_X1 port map( A1 => n59943, A2 => n61079, B1 => n3553, B2 => 
                           n59939, ZN => n10712);
   U4777 : OAI22_X1 port map( A1 => n59944, A2 => n61093, B1 => n3552, B2 => 
                           n59939, ZN => n10713);
   U4778 : OAI22_X1 port map( A1 => n59944, A2 => n61107, B1 => n3551, B2 => 
                           n59939, ZN => n10714);
   U4779 : OAI22_X1 port map( A1 => n59944, A2 => n61121, B1 => n3550, B2 => 
                           n59939, ZN => n10715);
   U4780 : OAI22_X1 port map( A1 => n59944, A2 => n61135, B1 => n3549, B2 => 
                           n59939, ZN => n10716);
   U4781 : OAI22_X1 port map( A1 => n59931, A2 => n61974, B1 => n3548, B2 => 
                           n59930, ZN => n10661);
   U4782 : OAI22_X1 port map( A1 => n59931, A2 => n61988, B1 => n3547, B2 => 
                           n59930, ZN => n10662);
   U4783 : OAI22_X1 port map( A1 => n59931, A2 => n62002, B1 => n3546, B2 => 
                           n59930, ZN => n10663);
   U4784 : OAI22_X1 port map( A1 => n59931, A2 => n62016, B1 => n3545, B2 => 
                           n59930, ZN => n10664);
   U4785 : OAI22_X1 port map( A1 => n59931, A2 => n62030, B1 => n3544, B2 => 
                           n59930, ZN => n10665);
   U4786 : OAI22_X1 port map( A1 => n59932, A2 => n62044, B1 => n3543, B2 => 
                           n59930, ZN => n10666);
   U4787 : OAI22_X1 port map( A1 => n59932, A2 => n62058, B1 => n3542, B2 => 
                           n59930, ZN => n10667);
   U4788 : OAI22_X1 port map( A1 => n59932, A2 => n62072, B1 => n3541, B2 => 
                           n59930, ZN => n10668);
   U4789 : OAI22_X1 port map( A1 => n59932, A2 => n62086, B1 => n3540, B2 => 
                           n59930, ZN => n10669);
   U4790 : OAI22_X1 port map( A1 => n59932, A2 => n62100, B1 => n3539, B2 => 
                           n59930, ZN => n10670);
   U4791 : OAI22_X1 port map( A1 => n59933, A2 => n62114, B1 => n3538, B2 => 
                           n59930, ZN => n10671);
   U4792 : OAI22_X1 port map( A1 => n59933, A2 => n60967, B1 => n3537, B2 => 
                           n59930, ZN => n10672);
   U4793 : OAI22_X1 port map( A1 => n59933, A2 => n60981, B1 => n3536, B2 => 
                           n15249, ZN => n10673);
   U4794 : OAI22_X1 port map( A1 => n59933, A2 => n60995, B1 => n3535, B2 => 
                           n15249, ZN => n10674);
   U4795 : OAI22_X1 port map( A1 => n59933, A2 => n61009, B1 => n3534, B2 => 
                           n15249, ZN => n10675);
   U4796 : OAI22_X1 port map( A1 => n59934, A2 => n61023, B1 => n3533, B2 => 
                           n15249, ZN => n10676);
   U4797 : OAI22_X1 port map( A1 => n59934, A2 => n61037, B1 => n3532, B2 => 
                           n15249, ZN => n10677);
   U4798 : OAI22_X1 port map( A1 => n59934, A2 => n61051, B1 => n3531, B2 => 
                           n15249, ZN => n10678);
   U4799 : OAI22_X1 port map( A1 => n59934, A2 => n61065, B1 => n3530, B2 => 
                           n15249, ZN => n10679);
   U4800 : OAI22_X1 port map( A1 => n59934, A2 => n61079, B1 => n3529, B2 => 
                           n59930, ZN => n10680);
   U4801 : OAI22_X1 port map( A1 => n59935, A2 => n61093, B1 => n3528, B2 => 
                           n59930, ZN => n10681);
   U4802 : OAI22_X1 port map( A1 => n59935, A2 => n61107, B1 => n3527, B2 => 
                           n59930, ZN => n10682);
   U4803 : OAI22_X1 port map( A1 => n59935, A2 => n61121, B1 => n3526, B2 => 
                           n59930, ZN => n10683);
   U4804 : OAI22_X1 port map( A1 => n59935, A2 => n61135, B1 => n3525, B2 => 
                           n59930, ZN => n10684);
   U4805 : OAI22_X1 port map( A1 => n59922, A2 => n61974, B1 => n3524, B2 => 
                           n59921, ZN => n10629);
   U4806 : OAI22_X1 port map( A1 => n59922, A2 => n61988, B1 => n3523, B2 => 
                           n59921, ZN => n10630);
   U4807 : OAI22_X1 port map( A1 => n59922, A2 => n62002, B1 => n3522, B2 => 
                           n59921, ZN => n10631);
   U4808 : OAI22_X1 port map( A1 => n59922, A2 => n62016, B1 => n3521, B2 => 
                           n59921, ZN => n10632);
   U4809 : OAI22_X1 port map( A1 => n59922, A2 => n62030, B1 => n3520, B2 => 
                           n59921, ZN => n10633);
   U4810 : OAI22_X1 port map( A1 => n59923, A2 => n62044, B1 => n3519, B2 => 
                           n59921, ZN => n10634);
   U4811 : OAI22_X1 port map( A1 => n59923, A2 => n62058, B1 => n3518, B2 => 
                           n59921, ZN => n10635);
   U4812 : OAI22_X1 port map( A1 => n59923, A2 => n62072, B1 => n3517, B2 => 
                           n59921, ZN => n10636);
   U4813 : OAI22_X1 port map( A1 => n59923, A2 => n62086, B1 => n3516, B2 => 
                           n59921, ZN => n10637);
   U4814 : OAI22_X1 port map( A1 => n59923, A2 => n62100, B1 => n3515, B2 => 
                           n59921, ZN => n10638);
   U4815 : OAI22_X1 port map( A1 => n59924, A2 => n62114, B1 => n3514, B2 => 
                           n59921, ZN => n10639);
   U4816 : OAI22_X1 port map( A1 => n59924, A2 => n60967, B1 => n3513, B2 => 
                           n59921, ZN => n10640);
   U4817 : OAI22_X1 port map( A1 => n59924, A2 => n60981, B1 => n3512, B2 => 
                           n15250, ZN => n10641);
   U4818 : OAI22_X1 port map( A1 => n59924, A2 => n60995, B1 => n3511, B2 => 
                           n15250, ZN => n10642);
   U4819 : OAI22_X1 port map( A1 => n59924, A2 => n61009, B1 => n3510, B2 => 
                           n15250, ZN => n10643);
   U4820 : OAI22_X1 port map( A1 => n59925, A2 => n61023, B1 => n3509, B2 => 
                           n15250, ZN => n10644);
   U4821 : OAI22_X1 port map( A1 => n59925, A2 => n61037, B1 => n3508, B2 => 
                           n15250, ZN => n10645);
   U4822 : OAI22_X1 port map( A1 => n59925, A2 => n61051, B1 => n3507, B2 => 
                           n15250, ZN => n10646);
   U4823 : OAI22_X1 port map( A1 => n59925, A2 => n61065, B1 => n3506, B2 => 
                           n15250, ZN => n10647);
   U4824 : OAI22_X1 port map( A1 => n59925, A2 => n61079, B1 => n3505, B2 => 
                           n59921, ZN => n10648);
   U4825 : OAI22_X1 port map( A1 => n59926, A2 => n61093, B1 => n3504, B2 => 
                           n59921, ZN => n10649);
   U4826 : OAI22_X1 port map( A1 => n59926, A2 => n61107, B1 => n3503, B2 => 
                           n59921, ZN => n10650);
   U4827 : OAI22_X1 port map( A1 => n59926, A2 => n61121, B1 => n3502, B2 => 
                           n59921, ZN => n10651);
   U4828 : OAI22_X1 port map( A1 => n59926, A2 => n61135, B1 => n3501, B2 => 
                           n59921, ZN => n10652);
   U4829 : OAI22_X1 port map( A1 => n59868, A2 => n61975, B1 => n3380, B2 => 
                           n59867, ZN => n10437);
   U4830 : OAI22_X1 port map( A1 => n59868, A2 => n61989, B1 => n3379, B2 => 
                           n59867, ZN => n10438);
   U4831 : OAI22_X1 port map( A1 => n59868, A2 => n62003, B1 => n3378, B2 => 
                           n59867, ZN => n10439);
   U4832 : OAI22_X1 port map( A1 => n59868, A2 => n62017, B1 => n3377, B2 => 
                           n59867, ZN => n10440);
   U4833 : OAI22_X1 port map( A1 => n59868, A2 => n62031, B1 => n3376, B2 => 
                           n59867, ZN => n10441);
   U4834 : OAI22_X1 port map( A1 => n59869, A2 => n62045, B1 => n3375, B2 => 
                           n59867, ZN => n10442);
   U4835 : OAI22_X1 port map( A1 => n59869, A2 => n62059, B1 => n3374, B2 => 
                           n59867, ZN => n10443);
   U4836 : OAI22_X1 port map( A1 => n59869, A2 => n62073, B1 => n3373, B2 => 
                           n59867, ZN => n10444);
   U4837 : OAI22_X1 port map( A1 => n59869, A2 => n62087, B1 => n3372, B2 => 
                           n59867, ZN => n10445);
   U4838 : OAI22_X1 port map( A1 => n59869, A2 => n62101, B1 => n3371, B2 => 
                           n59867, ZN => n10446);
   U4839 : OAI22_X1 port map( A1 => n59870, A2 => n62115, B1 => n3370, B2 => 
                           n59867, ZN => n10447);
   U4840 : OAI22_X1 port map( A1 => n59870, A2 => n60968, B1 => n3369, B2 => 
                           n59867, ZN => n10448);
   U4841 : OAI22_X1 port map( A1 => n59870, A2 => n60982, B1 => n3368, B2 => 
                           n15258, ZN => n10449);
   U4842 : OAI22_X1 port map( A1 => n59870, A2 => n60996, B1 => n3367, B2 => 
                           n15258, ZN => n10450);
   U4843 : OAI22_X1 port map( A1 => n59870, A2 => n61010, B1 => n3366, B2 => 
                           n15258, ZN => n10451);
   U4844 : OAI22_X1 port map( A1 => n59871, A2 => n61024, B1 => n3365, B2 => 
                           n15258, ZN => n10452);
   U4845 : OAI22_X1 port map( A1 => n59871, A2 => n61038, B1 => n3364, B2 => 
                           n15258, ZN => n10453);
   U4846 : OAI22_X1 port map( A1 => n59871, A2 => n61052, B1 => n3363, B2 => 
                           n15258, ZN => n10454);
   U4847 : OAI22_X1 port map( A1 => n59871, A2 => n61066, B1 => n3362, B2 => 
                           n15258, ZN => n10455);
   U4848 : OAI22_X1 port map( A1 => n59871, A2 => n61080, B1 => n3361, B2 => 
                           n59867, ZN => n10456);
   U4849 : OAI22_X1 port map( A1 => n59872, A2 => n61094, B1 => n3360, B2 => 
                           n59867, ZN => n10457);
   U4850 : OAI22_X1 port map( A1 => n59872, A2 => n61108, B1 => n3359, B2 => 
                           n59867, ZN => n10458);
   U4851 : OAI22_X1 port map( A1 => n59872, A2 => n61122, B1 => n3358, B2 => 
                           n59867, ZN => n10459);
   U4852 : OAI22_X1 port map( A1 => n59872, A2 => n61136, B1 => n3357, B2 => 
                           n59867, ZN => n10460);
   U4853 : OAI22_X1 port map( A1 => n59859, A2 => n61975, B1 => n3356, B2 => 
                           n59858, ZN => n10405);
   U4854 : OAI22_X1 port map( A1 => n59859, A2 => n61989, B1 => n3355, B2 => 
                           n59858, ZN => n10406);
   U4855 : OAI22_X1 port map( A1 => n59859, A2 => n62003, B1 => n3354, B2 => 
                           n59858, ZN => n10407);
   U4856 : OAI22_X1 port map( A1 => n59859, A2 => n62017, B1 => n3353, B2 => 
                           n59858, ZN => n10408);
   U4857 : OAI22_X1 port map( A1 => n59859, A2 => n62031, B1 => n3352, B2 => 
                           n59858, ZN => n10409);
   U4858 : OAI22_X1 port map( A1 => n59860, A2 => n62045, B1 => n3351, B2 => 
                           n59858, ZN => n10410);
   U4859 : OAI22_X1 port map( A1 => n59860, A2 => n62059, B1 => n3350, B2 => 
                           n59858, ZN => n10411);
   U4860 : OAI22_X1 port map( A1 => n59860, A2 => n62073, B1 => n3349, B2 => 
                           n59858, ZN => n10412);
   U4861 : OAI22_X1 port map( A1 => n59860, A2 => n62087, B1 => n3348, B2 => 
                           n59858, ZN => n10413);
   U4862 : OAI22_X1 port map( A1 => n59860, A2 => n62101, B1 => n3347, B2 => 
                           n59858, ZN => n10414);
   U4863 : OAI22_X1 port map( A1 => n59861, A2 => n62115, B1 => n3346, B2 => 
                           n59858, ZN => n10415);
   U4864 : OAI22_X1 port map( A1 => n59861, A2 => n60968, B1 => n3345, B2 => 
                           n59858, ZN => n10416);
   U4865 : OAI22_X1 port map( A1 => n59861, A2 => n60982, B1 => n3344, B2 => 
                           n15260, ZN => n10417);
   U4866 : OAI22_X1 port map( A1 => n59861, A2 => n60996, B1 => n3343, B2 => 
                           n15260, ZN => n10418);
   U4867 : OAI22_X1 port map( A1 => n59861, A2 => n61010, B1 => n3342, B2 => 
                           n15260, ZN => n10419);
   U4868 : OAI22_X1 port map( A1 => n59862, A2 => n61024, B1 => n3341, B2 => 
                           n15260, ZN => n10420);
   U4869 : OAI22_X1 port map( A1 => n59862, A2 => n61038, B1 => n3340, B2 => 
                           n15260, ZN => n10421);
   U4870 : OAI22_X1 port map( A1 => n59862, A2 => n61052, B1 => n3339, B2 => 
                           n15260, ZN => n10422);
   U4871 : OAI22_X1 port map( A1 => n59862, A2 => n61066, B1 => n3338, B2 => 
                           n15260, ZN => n10423);
   U4872 : OAI22_X1 port map( A1 => n59862, A2 => n61080, B1 => n3337, B2 => 
                           n59858, ZN => n10424);
   U4873 : OAI22_X1 port map( A1 => n59863, A2 => n61094, B1 => n3336, B2 => 
                           n59858, ZN => n10425);
   U4874 : OAI22_X1 port map( A1 => n59863, A2 => n61108, B1 => n3335, B2 => 
                           n59858, ZN => n10426);
   U4875 : OAI22_X1 port map( A1 => n59863, A2 => n61122, B1 => n3334, B2 => 
                           n59858, ZN => n10427);
   U4876 : OAI22_X1 port map( A1 => n59863, A2 => n61136, B1 => n3333, B2 => 
                           n59858, ZN => n10428);
   U4877 : OAI22_X1 port map( A1 => n59850, A2 => n61975, B1 => n3332, B2 => 
                           n59849, ZN => n10373);
   U4878 : OAI22_X1 port map( A1 => n59850, A2 => n61989, B1 => n3331, B2 => 
                           n59849, ZN => n10374);
   U4879 : OAI22_X1 port map( A1 => n59850, A2 => n62003, B1 => n3330, B2 => 
                           n59849, ZN => n10375);
   U4880 : OAI22_X1 port map( A1 => n59850, A2 => n62017, B1 => n3329, B2 => 
                           n59849, ZN => n10376);
   U4881 : OAI22_X1 port map( A1 => n59850, A2 => n62031, B1 => n3328, B2 => 
                           n59849, ZN => n10377);
   U4882 : OAI22_X1 port map( A1 => n59851, A2 => n62045, B1 => n3327, B2 => 
                           n59849, ZN => n10378);
   U4883 : OAI22_X1 port map( A1 => n59851, A2 => n62059, B1 => n3326, B2 => 
                           n59849, ZN => n10379);
   U4884 : OAI22_X1 port map( A1 => n59851, A2 => n62073, B1 => n3325, B2 => 
                           n59849, ZN => n10380);
   U4885 : OAI22_X1 port map( A1 => n59851, A2 => n62087, B1 => n3324, B2 => 
                           n59849, ZN => n10381);
   U4886 : OAI22_X1 port map( A1 => n59851, A2 => n62101, B1 => n3323, B2 => 
                           n59849, ZN => n10382);
   U4887 : OAI22_X1 port map( A1 => n59852, A2 => n62115, B1 => n3322, B2 => 
                           n59849, ZN => n10383);
   U4888 : OAI22_X1 port map( A1 => n59852, A2 => n60968, B1 => n3321, B2 => 
                           n59849, ZN => n10384);
   U4889 : OAI22_X1 port map( A1 => n59852, A2 => n60982, B1 => n3320, B2 => 
                           n15262, ZN => n10385);
   U4890 : OAI22_X1 port map( A1 => n59852, A2 => n60996, B1 => n3319, B2 => 
                           n15262, ZN => n10386);
   U4891 : OAI22_X1 port map( A1 => n59852, A2 => n61010, B1 => n3318, B2 => 
                           n15262, ZN => n10387);
   U4892 : OAI22_X1 port map( A1 => n59853, A2 => n61024, B1 => n3317, B2 => 
                           n15262, ZN => n10388);
   U4893 : OAI22_X1 port map( A1 => n59853, A2 => n61038, B1 => n3316, B2 => 
                           n15262, ZN => n10389);
   U4894 : OAI22_X1 port map( A1 => n59853, A2 => n61052, B1 => n3315, B2 => 
                           n15262, ZN => n10390);
   U4895 : OAI22_X1 port map( A1 => n59853, A2 => n61066, B1 => n3314, B2 => 
                           n15262, ZN => n10391);
   U4896 : OAI22_X1 port map( A1 => n59853, A2 => n61080, B1 => n3313, B2 => 
                           n59849, ZN => n10392);
   U4897 : OAI22_X1 port map( A1 => n59854, A2 => n61094, B1 => n3312, B2 => 
                           n59849, ZN => n10393);
   U4898 : OAI22_X1 port map( A1 => n59854, A2 => n61108, B1 => n3311, B2 => 
                           n59849, ZN => n10394);
   U4899 : OAI22_X1 port map( A1 => n59854, A2 => n61122, B1 => n3310, B2 => 
                           n59849, ZN => n10395);
   U4900 : OAI22_X1 port map( A1 => n59854, A2 => n61136, B1 => n3309, B2 => 
                           n59849, ZN => n10396);
   U4901 : OAI22_X1 port map( A1 => n59841, A2 => n61975, B1 => n3308, B2 => 
                           n59840, ZN => n10341);
   U4902 : OAI22_X1 port map( A1 => n59841, A2 => n61989, B1 => n3307, B2 => 
                           n59840, ZN => n10342);
   U4903 : OAI22_X1 port map( A1 => n59841, A2 => n62003, B1 => n3306, B2 => 
                           n59840, ZN => n10343);
   U4904 : OAI22_X1 port map( A1 => n59841, A2 => n62017, B1 => n3305, B2 => 
                           n59840, ZN => n10344);
   U4905 : OAI22_X1 port map( A1 => n59841, A2 => n62031, B1 => n3304, B2 => 
                           n59840, ZN => n10345);
   U4906 : OAI22_X1 port map( A1 => n59842, A2 => n62045, B1 => n3303, B2 => 
                           n59840, ZN => n10346);
   U4907 : OAI22_X1 port map( A1 => n59842, A2 => n62059, B1 => n3302, B2 => 
                           n59840, ZN => n10347);
   U4908 : OAI22_X1 port map( A1 => n59842, A2 => n62073, B1 => n3301, B2 => 
                           n59840, ZN => n10348);
   U4909 : OAI22_X1 port map( A1 => n59842, A2 => n62087, B1 => n3300, B2 => 
                           n59840, ZN => n10349);
   U4910 : OAI22_X1 port map( A1 => n59842, A2 => n62101, B1 => n3299, B2 => 
                           n59840, ZN => n10350);
   U4911 : OAI22_X1 port map( A1 => n59843, A2 => n62115, B1 => n3298, B2 => 
                           n59840, ZN => n10351);
   U4912 : OAI22_X1 port map( A1 => n59843, A2 => n60968, B1 => n3297, B2 => 
                           n59840, ZN => n10352);
   U4913 : OAI22_X1 port map( A1 => n59843, A2 => n60982, B1 => n3296, B2 => 
                           n15264, ZN => n10353);
   U4914 : OAI22_X1 port map( A1 => n59843, A2 => n60996, B1 => n3295, B2 => 
                           n15264, ZN => n10354);
   U4915 : OAI22_X1 port map( A1 => n59843, A2 => n61010, B1 => n3294, B2 => 
                           n15264, ZN => n10355);
   U4916 : OAI22_X1 port map( A1 => n59844, A2 => n61024, B1 => n3293, B2 => 
                           n15264, ZN => n10356);
   U4917 : OAI22_X1 port map( A1 => n59844, A2 => n61038, B1 => n3292, B2 => 
                           n15264, ZN => n10357);
   U4918 : OAI22_X1 port map( A1 => n59844, A2 => n61052, B1 => n3291, B2 => 
                           n15264, ZN => n10358);
   U4919 : OAI22_X1 port map( A1 => n59844, A2 => n61066, B1 => n3290, B2 => 
                           n15264, ZN => n10359);
   U4920 : OAI22_X1 port map( A1 => n59844, A2 => n61080, B1 => n3289, B2 => 
                           n59840, ZN => n10360);
   U4921 : OAI22_X1 port map( A1 => n59845, A2 => n61094, B1 => n3288, B2 => 
                           n59840, ZN => n10361);
   U4922 : OAI22_X1 port map( A1 => n59845, A2 => n61108, B1 => n3287, B2 => 
                           n59840, ZN => n10362);
   U4923 : OAI22_X1 port map( A1 => n59845, A2 => n61122, B1 => n3286, B2 => 
                           n59840, ZN => n10363);
   U4924 : OAI22_X1 port map( A1 => n59845, A2 => n61136, B1 => n3285, B2 => 
                           n59840, ZN => n10364);
   U4925 : OAI22_X1 port map( A1 => n60597, A2 => n61968, B1 => n3256, B2 => 
                           n60596, ZN => n13029);
   U4926 : OAI22_X1 port map( A1 => n60597, A2 => n61982, B1 => n3255, B2 => 
                           n60596, ZN => n13030);
   U4927 : OAI22_X1 port map( A1 => n60597, A2 => n61996, B1 => n3254, B2 => 
                           n60596, ZN => n13031);
   U4928 : OAI22_X1 port map( A1 => n60597, A2 => n62010, B1 => n3253, B2 => 
                           n60596, ZN => n13032);
   U4929 : OAI22_X1 port map( A1 => n60597, A2 => n62024, B1 => n3252, B2 => 
                           n60596, ZN => n13033);
   U4930 : OAI22_X1 port map( A1 => n60598, A2 => n62038, B1 => n3251, B2 => 
                           n60596, ZN => n13034);
   U4931 : OAI22_X1 port map( A1 => n60598, A2 => n62052, B1 => n3250, B2 => 
                           n60596, ZN => n13035);
   U4932 : OAI22_X1 port map( A1 => n60598, A2 => n62066, B1 => n3249, B2 => 
                           n60596, ZN => n13036);
   U4933 : OAI22_X1 port map( A1 => n60598, A2 => n62080, B1 => n3248, B2 => 
                           n60596, ZN => n13037);
   U4934 : OAI22_X1 port map( A1 => n60598, A2 => n62094, B1 => n3247, B2 => 
                           n60596, ZN => n13038);
   U4935 : OAI22_X1 port map( A1 => n60599, A2 => n62108, B1 => n3246, B2 => 
                           n60596, ZN => n13039);
   U4936 : OAI22_X1 port map( A1 => n60599, A2 => n60961, B1 => n3245, B2 => 
                           n60596, ZN => n13040);
   U4937 : OAI22_X1 port map( A1 => n60599, A2 => n60975, B1 => n3244, B2 => 
                           n15155, ZN => n13041);
   U4938 : OAI22_X1 port map( A1 => n60599, A2 => n60989, B1 => n3243, B2 => 
                           n15155, ZN => n13042);
   U4939 : OAI22_X1 port map( A1 => n60599, A2 => n61003, B1 => n3242, B2 => 
                           n15155, ZN => n13043);
   U4940 : OAI22_X1 port map( A1 => n60600, A2 => n61017, B1 => n3241, B2 => 
                           n15155, ZN => n13044);
   U4941 : OAI22_X1 port map( A1 => n60600, A2 => n61031, B1 => n3240, B2 => 
                           n15155, ZN => n13045);
   U4942 : OAI22_X1 port map( A1 => n60600, A2 => n61045, B1 => n3239, B2 => 
                           n15155, ZN => n13046);
   U4943 : OAI22_X1 port map( A1 => n60600, A2 => n61059, B1 => n3238, B2 => 
                           n15155, ZN => n13047);
   U4944 : OAI22_X1 port map( A1 => n60600, A2 => n61073, B1 => n3237, B2 => 
                           n60596, ZN => n13048);
   U4945 : OAI22_X1 port map( A1 => n60601, A2 => n61087, B1 => n3236, B2 => 
                           n60596, ZN => n13049);
   U4946 : OAI22_X1 port map( A1 => n60601, A2 => n61101, B1 => n3235, B2 => 
                           n60596, ZN => n13050);
   U4947 : OAI22_X1 port map( A1 => n60601, A2 => n61115, B1 => n3234, B2 => 
                           n60596, ZN => n13051);
   U4948 : OAI22_X1 port map( A1 => n60601, A2 => n61129, B1 => n3233, B2 => 
                           n60596, ZN => n13052);
   U4949 : OAI22_X1 port map( A1 => n60588, A2 => n61968, B1 => n3232, B2 => 
                           n60587, ZN => n12997);
   U4950 : OAI22_X1 port map( A1 => n60588, A2 => n61982, B1 => n3231, B2 => 
                           n60587, ZN => n12998);
   U4951 : OAI22_X1 port map( A1 => n60588, A2 => n61996, B1 => n3230, B2 => 
                           n60587, ZN => n12999);
   U4952 : OAI22_X1 port map( A1 => n60588, A2 => n62010, B1 => n3229, B2 => 
                           n60587, ZN => n13000);
   U4953 : OAI22_X1 port map( A1 => n60588, A2 => n62024, B1 => n3228, B2 => 
                           n60587, ZN => n13001);
   U4954 : OAI22_X1 port map( A1 => n60589, A2 => n62038, B1 => n3227, B2 => 
                           n60587, ZN => n13002);
   U4955 : OAI22_X1 port map( A1 => n60589, A2 => n62052, B1 => n3226, B2 => 
                           n60587, ZN => n13003);
   U4956 : OAI22_X1 port map( A1 => n60589, A2 => n62066, B1 => n3225, B2 => 
                           n60587, ZN => n13004);
   U4957 : OAI22_X1 port map( A1 => n60589, A2 => n62080, B1 => n3224, B2 => 
                           n60587, ZN => n13005);
   U4958 : OAI22_X1 port map( A1 => n60589, A2 => n62094, B1 => n3223, B2 => 
                           n60587, ZN => n13006);
   U4959 : OAI22_X1 port map( A1 => n60590, A2 => n62108, B1 => n3222, B2 => 
                           n60587, ZN => n13007);
   U4960 : OAI22_X1 port map( A1 => n60590, A2 => n60961, B1 => n3221, B2 => 
                           n60587, ZN => n13008);
   U4961 : OAI22_X1 port map( A1 => n60590, A2 => n60975, B1 => n3220, B2 => 
                           n15156, ZN => n13009);
   U4962 : OAI22_X1 port map( A1 => n60590, A2 => n60989, B1 => n3219, B2 => 
                           n15156, ZN => n13010);
   U4963 : OAI22_X1 port map( A1 => n60590, A2 => n61003, B1 => n3218, B2 => 
                           n15156, ZN => n13011);
   U4964 : OAI22_X1 port map( A1 => n60591, A2 => n61017, B1 => n3217, B2 => 
                           n15156, ZN => n13012);
   U4965 : OAI22_X1 port map( A1 => n60591, A2 => n61031, B1 => n3216, B2 => 
                           n15156, ZN => n13013);
   U4966 : OAI22_X1 port map( A1 => n60591, A2 => n61045, B1 => n3215, B2 => 
                           n15156, ZN => n13014);
   U4967 : OAI22_X1 port map( A1 => n60591, A2 => n61059, B1 => n3214, B2 => 
                           n15156, ZN => n13015);
   U4968 : OAI22_X1 port map( A1 => n60591, A2 => n61073, B1 => n3213, B2 => 
                           n60587, ZN => n13016);
   U4969 : OAI22_X1 port map( A1 => n60592, A2 => n61087, B1 => n3212, B2 => 
                           n60587, ZN => n13017);
   U4970 : OAI22_X1 port map( A1 => n60592, A2 => n61101, B1 => n3211, B2 => 
                           n60587, ZN => n13018);
   U4971 : OAI22_X1 port map( A1 => n60592, A2 => n61115, B1 => n3210, B2 => 
                           n60587, ZN => n13019);
   U4972 : OAI22_X1 port map( A1 => n60592, A2 => n61129, B1 => n3209, B2 => 
                           n60587, ZN => n13020);
   U4973 : OAI22_X1 port map( A1 => n60561, A2 => n61968, B1 => n3208, B2 => 
                           n60560, ZN => n12901);
   U4974 : OAI22_X1 port map( A1 => n60561, A2 => n61982, B1 => n3207, B2 => 
                           n60560, ZN => n12902);
   U4975 : OAI22_X1 port map( A1 => n60561, A2 => n61996, B1 => n3206, B2 => 
                           n60560, ZN => n12903);
   U4976 : OAI22_X1 port map( A1 => n60561, A2 => n62010, B1 => n3205, B2 => 
                           n60560, ZN => n12904);
   U4977 : OAI22_X1 port map( A1 => n60561, A2 => n62024, B1 => n3204, B2 => 
                           n60560, ZN => n12905);
   U4978 : OAI22_X1 port map( A1 => n60562, A2 => n62038, B1 => n3203, B2 => 
                           n60560, ZN => n12906);
   U4979 : OAI22_X1 port map( A1 => n60562, A2 => n62052, B1 => n3202, B2 => 
                           n60560, ZN => n12907);
   U4980 : OAI22_X1 port map( A1 => n60562, A2 => n62066, B1 => n3201, B2 => 
                           n60560, ZN => n12908);
   U4981 : OAI22_X1 port map( A1 => n60562, A2 => n62080, B1 => n3200, B2 => 
                           n60560, ZN => n12909);
   U4982 : OAI22_X1 port map( A1 => n60562, A2 => n62094, B1 => n3199, B2 => 
                           n60560, ZN => n12910);
   U4983 : OAI22_X1 port map( A1 => n60552, A2 => n61968, B1 => n3198, B2 => 
                           n60551, ZN => n12869);
   U4984 : OAI22_X1 port map( A1 => n60552, A2 => n61982, B1 => n3197, B2 => 
                           n60551, ZN => n12870);
   U4985 : OAI22_X1 port map( A1 => n60552, A2 => n61996, B1 => n3196, B2 => 
                           n60551, ZN => n12871);
   U4986 : OAI22_X1 port map( A1 => n60552, A2 => n62010, B1 => n3195, B2 => 
                           n60551, ZN => n12872);
   U4987 : OAI22_X1 port map( A1 => n60552, A2 => n62024, B1 => n3194, B2 => 
                           n60551, ZN => n12873);
   U4988 : OAI22_X1 port map( A1 => n60553, A2 => n62038, B1 => n3193, B2 => 
                           n60551, ZN => n12874);
   U4989 : OAI22_X1 port map( A1 => n60553, A2 => n62052, B1 => n3192, B2 => 
                           n60551, ZN => n12875);
   U4990 : OAI22_X1 port map( A1 => n60553, A2 => n62066, B1 => n3191, B2 => 
                           n60551, ZN => n12876);
   U4991 : OAI22_X1 port map( A1 => n60553, A2 => n62080, B1 => n3190, B2 => 
                           n60551, ZN => n12877);
   U4992 : OAI22_X1 port map( A1 => n60553, A2 => n62094, B1 => n3189, B2 => 
                           n60551, ZN => n12878);
   U4993 : OAI22_X1 port map( A1 => n60554, A2 => n62108, B1 => n3188, B2 => 
                           n60551, ZN => n12879);
   U4994 : OAI22_X1 port map( A1 => n60554, A2 => n60961, B1 => n3187, B2 => 
                           n60551, ZN => n12880);
   U4995 : OAI22_X1 port map( A1 => n60554, A2 => n60975, B1 => n3186, B2 => 
                           n15160, ZN => n12881);
   U4996 : OAI22_X1 port map( A1 => n60554, A2 => n60989, B1 => n3185, B2 => 
                           n15160, ZN => n12882);
   U4997 : OAI22_X1 port map( A1 => n60554, A2 => n61003, B1 => n3184, B2 => 
                           n15160, ZN => n12883);
   U4998 : OAI22_X1 port map( A1 => n60555, A2 => n61017, B1 => n3183, B2 => 
                           n15160, ZN => n12884);
   U4999 : OAI22_X1 port map( A1 => n60555, A2 => n61031, B1 => n3182, B2 => 
                           n15160, ZN => n12885);
   U5000 : OAI22_X1 port map( A1 => n60555, A2 => n61045, B1 => n3181, B2 => 
                           n15160, ZN => n12886);
   U5001 : OAI22_X1 port map( A1 => n60555, A2 => n61059, B1 => n3180, B2 => 
                           n15160, ZN => n12887);
   U5002 : OAI22_X1 port map( A1 => n60555, A2 => n61073, B1 => n3179, B2 => 
                           n60551, ZN => n12888);
   U5003 : OAI22_X1 port map( A1 => n60556, A2 => n61087, B1 => n3178, B2 => 
                           n60551, ZN => n12889);
   U5004 : OAI22_X1 port map( A1 => n60556, A2 => n61101, B1 => n3177, B2 => 
                           n60551, ZN => n12890);
   U5005 : OAI22_X1 port map( A1 => n60556, A2 => n61115, B1 => n3176, B2 => 
                           n60551, ZN => n12891);
   U5006 : OAI22_X1 port map( A1 => n60556, A2 => n61129, B1 => n3175, B2 => 
                           n60551, ZN => n12892);
   U5007 : OAI22_X1 port map( A1 => n60534, A2 => n61968, B1 => n3174, B2 => 
                           n60533, ZN => n12805);
   U5008 : OAI22_X1 port map( A1 => n60534, A2 => n61982, B1 => n3173, B2 => 
                           n60533, ZN => n12806);
   U5009 : OAI22_X1 port map( A1 => n60534, A2 => n61996, B1 => n3172, B2 => 
                           n60533, ZN => n12807);
   U5010 : OAI22_X1 port map( A1 => n60534, A2 => n62010, B1 => n3171, B2 => 
                           n60533, ZN => n12808);
   U5011 : OAI22_X1 port map( A1 => n60534, A2 => n62024, B1 => n3170, B2 => 
                           n60533, ZN => n12809);
   U5012 : OAI22_X1 port map( A1 => n60535, A2 => n62038, B1 => n3169, B2 => 
                           n60533, ZN => n12810);
   U5013 : OAI22_X1 port map( A1 => n60535, A2 => n62052, B1 => n3168, B2 => 
                           n60533, ZN => n12811);
   U5014 : OAI22_X1 port map( A1 => n60535, A2 => n62066, B1 => n3167, B2 => 
                           n60533, ZN => n12812);
   U5015 : OAI22_X1 port map( A1 => n60535, A2 => n62080, B1 => n3166, B2 => 
                           n60533, ZN => n12813);
   U5016 : OAI22_X1 port map( A1 => n60535, A2 => n62094, B1 => n3165, B2 => 
                           n60533, ZN => n12814);
   U5017 : OAI22_X1 port map( A1 => n60536, A2 => n62108, B1 => n3164, B2 => 
                           n60533, ZN => n12815);
   U5018 : OAI22_X1 port map( A1 => n60536, A2 => n60961, B1 => n3163, B2 => 
                           n60533, ZN => n12816);
   U5019 : OAI22_X1 port map( A1 => n60536, A2 => n60975, B1 => n3162, B2 => 
                           n60533, ZN => n12817);
   U5020 : OAI22_X1 port map( A1 => n60536, A2 => n60989, B1 => n3161, B2 => 
                           n60533, ZN => n12818);
   U5021 : OAI22_X1 port map( A1 => n60525, A2 => n61968, B1 => n3160, B2 => 
                           n60524, ZN => n12773);
   U5022 : OAI22_X1 port map( A1 => n60525, A2 => n61982, B1 => n3159, B2 => 
                           n60524, ZN => n12774);
   U5023 : OAI22_X1 port map( A1 => n60525, A2 => n61996, B1 => n3158, B2 => 
                           n60524, ZN => n12775);
   U5024 : OAI22_X1 port map( A1 => n60525, A2 => n62010, B1 => n3157, B2 => 
                           n60524, ZN => n12776);
   U5025 : OAI22_X1 port map( A1 => n60525, A2 => n62024, B1 => n3156, B2 => 
                           n60524, ZN => n12777);
   U5026 : OAI22_X1 port map( A1 => n60526, A2 => n62038, B1 => n3155, B2 => 
                           n60524, ZN => n12778);
   U5027 : OAI22_X1 port map( A1 => n60526, A2 => n62052, B1 => n3154, B2 => 
                           n60524, ZN => n12779);
   U5028 : OAI22_X1 port map( A1 => n60526, A2 => n62066, B1 => n3153, B2 => 
                           n60524, ZN => n12780);
   U5029 : OAI22_X1 port map( A1 => n60526, A2 => n62080, B1 => n3152, B2 => 
                           n60524, ZN => n12781);
   U5030 : OAI22_X1 port map( A1 => n60526, A2 => n62094, B1 => n3151, B2 => 
                           n60524, ZN => n12782);
   U5031 : OAI22_X1 port map( A1 => n60507, A2 => n61969, B1 => n3150, B2 => 
                           n60506, ZN => n12709);
   U5032 : OAI22_X1 port map( A1 => n60507, A2 => n61983, B1 => n3149, B2 => 
                           n60506, ZN => n12710);
   U5033 : OAI22_X1 port map( A1 => n60507, A2 => n61997, B1 => n3148, B2 => 
                           n60506, ZN => n12711);
   U5034 : OAI22_X1 port map( A1 => n60507, A2 => n62011, B1 => n3147, B2 => 
                           n60506, ZN => n12712);
   U5035 : OAI22_X1 port map( A1 => n60507, A2 => n62025, B1 => n3146, B2 => 
                           n60506, ZN => n12713);
   U5036 : OAI22_X1 port map( A1 => n60508, A2 => n62039, B1 => n3145, B2 => 
                           n60506, ZN => n12714);
   U5037 : OAI22_X1 port map( A1 => n60508, A2 => n62053, B1 => n3144, B2 => 
                           n60506, ZN => n12715);
   U5038 : OAI22_X1 port map( A1 => n60508, A2 => n62067, B1 => n3143, B2 => 
                           n60506, ZN => n12716);
   U5039 : OAI22_X1 port map( A1 => n60508, A2 => n62081, B1 => n3142, B2 => 
                           n60506, ZN => n12717);
   U5040 : OAI22_X1 port map( A1 => n60508, A2 => n62095, B1 => n3141, B2 => 
                           n60506, ZN => n12718);
   U5041 : OAI22_X1 port map( A1 => n60509, A2 => n62109, B1 => n3140, B2 => 
                           n60506, ZN => n12719);
   U5042 : OAI22_X1 port map( A1 => n60509, A2 => n60962, B1 => n3139, B2 => 
                           n60506, ZN => n12720);
   U5043 : OAI22_X1 port map( A1 => n60509, A2 => n60976, B1 => n3138, B2 => 
                           n15166, ZN => n12721);
   U5044 : OAI22_X1 port map( A1 => n60509, A2 => n60990, B1 => n3137, B2 => 
                           n15166, ZN => n12722);
   U5045 : OAI22_X1 port map( A1 => n60509, A2 => n61004, B1 => n3136, B2 => 
                           n15166, ZN => n12723);
   U5046 : OAI22_X1 port map( A1 => n60510, A2 => n61018, B1 => n3135, B2 => 
                           n15166, ZN => n12724);
   U5047 : OAI22_X1 port map( A1 => n60510, A2 => n61032, B1 => n3134, B2 => 
                           n15166, ZN => n12725);
   U5048 : OAI22_X1 port map( A1 => n60510, A2 => n61046, B1 => n3133, B2 => 
                           n15166, ZN => n12726);
   U5049 : OAI22_X1 port map( A1 => n60510, A2 => n61060, B1 => n3132, B2 => 
                           n15166, ZN => n12727);
   U5050 : OAI22_X1 port map( A1 => n60510, A2 => n61074, B1 => n3131, B2 => 
                           n60506, ZN => n12728);
   U5051 : OAI22_X1 port map( A1 => n60511, A2 => n61088, B1 => n3130, B2 => 
                           n60506, ZN => n12729);
   U5052 : OAI22_X1 port map( A1 => n60511, A2 => n61102, B1 => n3129, B2 => 
                           n60506, ZN => n12730);
   U5053 : OAI22_X1 port map( A1 => n60511, A2 => n61116, B1 => n3128, B2 => 
                           n60506, ZN => n12731);
   U5054 : OAI22_X1 port map( A1 => n60511, A2 => n61130, B1 => n3127, B2 => 
                           n60506, ZN => n12732);
   U5055 : OAI22_X1 port map( A1 => n60462, A2 => n61969, B1 => n3054, B2 => 
                           n60461, ZN => n12549);
   U5056 : OAI22_X1 port map( A1 => n60462, A2 => n61983, B1 => n3053, B2 => 
                           n60461, ZN => n12550);
   U5057 : OAI22_X1 port map( A1 => n60462, A2 => n61997, B1 => n3052, B2 => 
                           n60461, ZN => n12551);
   U5058 : OAI22_X1 port map( A1 => n60462, A2 => n62011, B1 => n3051, B2 => 
                           n60461, ZN => n12552);
   U5059 : OAI22_X1 port map( A1 => n60462, A2 => n62025, B1 => n3050, B2 => 
                           n60461, ZN => n12553);
   U5060 : OAI22_X1 port map( A1 => n60463, A2 => n62039, B1 => n3049, B2 => 
                           n60461, ZN => n12554);
   U5061 : OAI22_X1 port map( A1 => n60463, A2 => n62053, B1 => n3048, B2 => 
                           n60461, ZN => n12555);
   U5062 : OAI22_X1 port map( A1 => n60463, A2 => n62067, B1 => n3047, B2 => 
                           n60461, ZN => n12556);
   U5063 : OAI22_X1 port map( A1 => n60463, A2 => n62081, B1 => n3046, B2 => 
                           n60461, ZN => n12557);
   U5064 : OAI22_X1 port map( A1 => n60463, A2 => n62095, B1 => n3045, B2 => 
                           n60461, ZN => n12558);
   U5065 : OAI22_X1 port map( A1 => n60464, A2 => n62109, B1 => n3044, B2 => 
                           n60461, ZN => n12559);
   U5066 : OAI22_X1 port map( A1 => n60464, A2 => n60962, B1 => n3043, B2 => 
                           n60461, ZN => n12560);
   U5067 : OAI22_X1 port map( A1 => n60464, A2 => n60976, B1 => n3042, B2 => 
                           n15178, ZN => n12561);
   U5068 : OAI22_X1 port map( A1 => n60464, A2 => n60990, B1 => n3041, B2 => 
                           n15178, ZN => n12562);
   U5069 : OAI22_X1 port map( A1 => n60464, A2 => n61004, B1 => n3040, B2 => 
                           n15178, ZN => n12563);
   U5070 : OAI22_X1 port map( A1 => n60465, A2 => n61018, B1 => n3039, B2 => 
                           n15178, ZN => n12564);
   U5071 : OAI22_X1 port map( A1 => n60465, A2 => n61032, B1 => n3038, B2 => 
                           n15178, ZN => n12565);
   U5072 : OAI22_X1 port map( A1 => n60465, A2 => n61046, B1 => n3037, B2 => 
                           n15178, ZN => n12566);
   U5073 : OAI22_X1 port map( A1 => n60465, A2 => n61060, B1 => n3036, B2 => 
                           n15178, ZN => n12567);
   U5074 : OAI22_X1 port map( A1 => n60465, A2 => n61074, B1 => n3035, B2 => 
                           n60461, ZN => n12568);
   U5075 : OAI22_X1 port map( A1 => n60466, A2 => n61088, B1 => n3034, B2 => 
                           n60461, ZN => n12569);
   U5076 : OAI22_X1 port map( A1 => n60466, A2 => n61102, B1 => n3033, B2 => 
                           n60461, ZN => n12570);
   U5077 : OAI22_X1 port map( A1 => n60466, A2 => n61116, B1 => n3032, B2 => 
                           n60461, ZN => n12571);
   U5078 : OAI22_X1 port map( A1 => n60466, A2 => n61130, B1 => n3031, B2 => 
                           n60461, ZN => n12572);
   U5079 : OAI22_X1 port map( A1 => n60444, A2 => n61969, B1 => n2958, B2 => 
                           n60443, ZN => n12485);
   U5080 : OAI22_X1 port map( A1 => n60444, A2 => n61983, B1 => n2957, B2 => 
                           n60443, ZN => n12486);
   U5081 : OAI22_X1 port map( A1 => n60444, A2 => n61997, B1 => n2956, B2 => 
                           n60443, ZN => n12487);
   U5082 : OAI22_X1 port map( A1 => n60444, A2 => n62011, B1 => n2955, B2 => 
                           n60443, ZN => n12488);
   U5083 : OAI22_X1 port map( A1 => n60444, A2 => n62025, B1 => n2954, B2 => 
                           n60443, ZN => n12489);
   U5084 : OAI22_X1 port map( A1 => n60445, A2 => n62039, B1 => n2953, B2 => 
                           n60443, ZN => n12490);
   U5085 : OAI22_X1 port map( A1 => n60445, A2 => n62053, B1 => n2952, B2 => 
                           n60443, ZN => n12491);
   U5086 : OAI22_X1 port map( A1 => n60445, A2 => n62067, B1 => n2951, B2 => 
                           n60443, ZN => n12492);
   U5087 : OAI22_X1 port map( A1 => n60445, A2 => n62081, B1 => n2950, B2 => 
                           n60443, ZN => n12493);
   U5088 : OAI22_X1 port map( A1 => n60445, A2 => n62095, B1 => n2949, B2 => 
                           n60443, ZN => n12494);
   U5089 : OAI22_X1 port map( A1 => n60446, A2 => n62109, B1 => n2948, B2 => 
                           n60443, ZN => n12495);
   U5090 : OAI22_X1 port map( A1 => n60446, A2 => n60962, B1 => n2947, B2 => 
                           n60443, ZN => n12496);
   U5091 : OAI22_X1 port map( A1 => n60446, A2 => n60976, B1 => n2946, B2 => 
                           n15180, ZN => n12497);
   U5092 : OAI22_X1 port map( A1 => n60446, A2 => n60990, B1 => n2945, B2 => 
                           n15180, ZN => n12498);
   U5093 : OAI22_X1 port map( A1 => n60446, A2 => n61004, B1 => n2944, B2 => 
                           n15180, ZN => n12499);
   U5094 : OAI22_X1 port map( A1 => n60447, A2 => n61018, B1 => n2943, B2 => 
                           n15180, ZN => n12500);
   U5095 : OAI22_X1 port map( A1 => n60447, A2 => n61032, B1 => n2942, B2 => 
                           n15180, ZN => n12501);
   U5096 : OAI22_X1 port map( A1 => n60447, A2 => n61046, B1 => n2941, B2 => 
                           n15180, ZN => n12502);
   U5097 : OAI22_X1 port map( A1 => n60447, A2 => n61060, B1 => n2940, B2 => 
                           n15180, ZN => n12503);
   U5098 : OAI22_X1 port map( A1 => n60447, A2 => n61074, B1 => n2939, B2 => 
                           n60443, ZN => n12504);
   U5099 : OAI22_X1 port map( A1 => n60448, A2 => n61088, B1 => n2938, B2 => 
                           n60443, ZN => n12505);
   U5100 : OAI22_X1 port map( A1 => n60448, A2 => n61102, B1 => n2937, B2 => 
                           n60443, ZN => n12506);
   U5101 : OAI22_X1 port map( A1 => n60448, A2 => n61116, B1 => n2936, B2 => 
                           n60443, ZN => n12507);
   U5102 : OAI22_X1 port map( A1 => n60448, A2 => n61130, B1 => n2935, B2 => 
                           n60443, ZN => n12508);
   U5103 : OAI22_X1 port map( A1 => n60435, A2 => n61969, B1 => n2934, B2 => 
                           n60434, ZN => n12453);
   U5104 : OAI22_X1 port map( A1 => n60435, A2 => n61983, B1 => n2933, B2 => 
                           n60434, ZN => n12454);
   U5105 : OAI22_X1 port map( A1 => n60435, A2 => n61997, B1 => n2932, B2 => 
                           n60434, ZN => n12455);
   U5106 : OAI22_X1 port map( A1 => n60435, A2 => n62011, B1 => n2931, B2 => 
                           n60434, ZN => n12456);
   U5107 : OAI22_X1 port map( A1 => n60435, A2 => n62025, B1 => n2930, B2 => 
                           n60434, ZN => n12457);
   U5108 : OAI22_X1 port map( A1 => n60436, A2 => n62039, B1 => n2929, B2 => 
                           n60434, ZN => n12458);
   U5109 : OAI22_X1 port map( A1 => n60436, A2 => n62053, B1 => n2928, B2 => 
                           n60434, ZN => n12459);
   U5110 : OAI22_X1 port map( A1 => n60436, A2 => n62067, B1 => n2927, B2 => 
                           n60434, ZN => n12460);
   U5111 : OAI22_X1 port map( A1 => n60436, A2 => n62081, B1 => n2926, B2 => 
                           n60434, ZN => n12461);
   U5112 : OAI22_X1 port map( A1 => n60436, A2 => n62095, B1 => n2925, B2 => 
                           n60434, ZN => n12462);
   U5113 : OAI22_X1 port map( A1 => n60437, A2 => n62109, B1 => n2908, B2 => 
                           n60434, ZN => n12463);
   U5114 : OAI22_X1 port map( A1 => n60437, A2 => n60962, B1 => n2907, B2 => 
                           n60434, ZN => n12464);
   U5115 : OAI22_X1 port map( A1 => n60437, A2 => n60976, B1 => n2886, B2 => 
                           n15181, ZN => n12465);
   U5116 : OAI22_X1 port map( A1 => n60437, A2 => n60990, B1 => n2885, B2 => 
                           n15181, ZN => n12466);
   U5117 : OAI22_X1 port map( A1 => n60437, A2 => n61004, B1 => n2884, B2 => 
                           n15181, ZN => n12467);
   U5118 : OAI22_X1 port map( A1 => n60438, A2 => n61018, B1 => n2883, B2 => 
                           n15181, ZN => n12468);
   U5119 : OAI22_X1 port map( A1 => n60438, A2 => n61032, B1 => n2882, B2 => 
                           n15181, ZN => n12469);
   U5120 : OAI22_X1 port map( A1 => n60438, A2 => n61046, B1 => n2881, B2 => 
                           n15181, ZN => n12470);
   U5121 : OAI22_X1 port map( A1 => n60438, A2 => n61060, B1 => n2880, B2 => 
                           n15181, ZN => n12471);
   U5122 : OAI22_X1 port map( A1 => n60438, A2 => n61074, B1 => n2879, B2 => 
                           n60434, ZN => n12472);
   U5123 : OAI22_X1 port map( A1 => n60439, A2 => n61088, B1 => n2878, B2 => 
                           n60434, ZN => n12473);
   U5124 : OAI22_X1 port map( A1 => n60439, A2 => n61102, B1 => n2877, B2 => 
                           n60434, ZN => n12474);
   U5125 : OAI22_X1 port map( A1 => n60439, A2 => n61116, B1 => n2876, B2 => 
                           n60434, ZN => n12475);
   U5126 : OAI22_X1 port map( A1 => n60439, A2 => n61130, B1 => n2875, B2 => 
                           n60434, ZN => n12476);
   U5127 : OAI22_X1 port map( A1 => n60408, A2 => n61970, B1 => n2874, B2 => 
                           n60407, ZN => n12357);
   U5128 : OAI22_X1 port map( A1 => n60408, A2 => n61984, B1 => n2873, B2 => 
                           n60407, ZN => n12358);
   U5129 : OAI22_X1 port map( A1 => n60408, A2 => n61998, B1 => n2872, B2 => 
                           n60407, ZN => n12359);
   U5130 : OAI22_X1 port map( A1 => n60408, A2 => n62012, B1 => n2871, B2 => 
                           n60407, ZN => n12360);
   U5131 : OAI22_X1 port map( A1 => n60408, A2 => n62026, B1 => n2870, B2 => 
                           n60407, ZN => n12361);
   U5132 : OAI22_X1 port map( A1 => n60409, A2 => n62040, B1 => n2869, B2 => 
                           n60407, ZN => n12362);
   U5133 : OAI22_X1 port map( A1 => n60409, A2 => n62054, B1 => n2868, B2 => 
                           n60407, ZN => n12363);
   U5134 : OAI22_X1 port map( A1 => n60409, A2 => n62068, B1 => n2867, B2 => 
                           n60407, ZN => n12364);
   U5135 : OAI22_X1 port map( A1 => n60409, A2 => n62082, B1 => n2866, B2 => 
                           n60407, ZN => n12365);
   U5136 : OAI22_X1 port map( A1 => n60409, A2 => n62096, B1 => n2865, B2 => 
                           n60407, ZN => n12366);
   U5137 : OAI22_X1 port map( A1 => n60410, A2 => n62110, B1 => n2864, B2 => 
                           n60407, ZN => n12367);
   U5138 : OAI22_X1 port map( A1 => n60410, A2 => n60963, B1 => n2863, B2 => 
                           n60407, ZN => n12368);
   U5139 : OAI22_X1 port map( A1 => n60410, A2 => n60977, B1 => n2862, B2 => 
                           n15184, ZN => n12369);
   U5140 : OAI22_X1 port map( A1 => n60410, A2 => n60991, B1 => n2861, B2 => 
                           n15184, ZN => n12370);
   U5141 : OAI22_X1 port map( A1 => n60410, A2 => n61005, B1 => n2860, B2 => 
                           n15184, ZN => n12371);
   U5142 : OAI22_X1 port map( A1 => n60411, A2 => n61019, B1 => n2859, B2 => 
                           n15184, ZN => n12372);
   U5143 : OAI22_X1 port map( A1 => n60411, A2 => n61033, B1 => n2858, B2 => 
                           n15184, ZN => n12373);
   U5144 : OAI22_X1 port map( A1 => n60411, A2 => n61047, B1 => n2857, B2 => 
                           n15184, ZN => n12374);
   U5145 : OAI22_X1 port map( A1 => n60411, A2 => n61061, B1 => n2856, B2 => 
                           n15184, ZN => n12375);
   U5146 : OAI22_X1 port map( A1 => n60411, A2 => n61075, B1 => n2855, B2 => 
                           n60407, ZN => n12376);
   U5147 : OAI22_X1 port map( A1 => n60412, A2 => n61089, B1 => n2854, B2 => 
                           n60407, ZN => n12377);
   U5148 : OAI22_X1 port map( A1 => n60412, A2 => n61103, B1 => n2853, B2 => 
                           n60407, ZN => n12378);
   U5149 : OAI22_X1 port map( A1 => n60412, A2 => n61117, B1 => n2852, B2 => 
                           n60407, ZN => n12379);
   U5150 : OAI22_X1 port map( A1 => n60412, A2 => n61131, B1 => n2851, B2 => 
                           n60407, ZN => n12380);
   U5151 : OAI22_X1 port map( A1 => n60399, A2 => n61970, B1 => n2850, B2 => 
                           n60398, ZN => n12325);
   U5152 : OAI22_X1 port map( A1 => n60399, A2 => n61984, B1 => n2849, B2 => 
                           n60398, ZN => n12326);
   U5153 : OAI22_X1 port map( A1 => n60399, A2 => n61998, B1 => n2848, B2 => 
                           n60398, ZN => n12327);
   U5154 : OAI22_X1 port map( A1 => n60399, A2 => n62012, B1 => n2847, B2 => 
                           n60398, ZN => n12328);
   U5155 : OAI22_X1 port map( A1 => n60399, A2 => n62026, B1 => n2846, B2 => 
                           n60398, ZN => n12329);
   U5156 : OAI22_X1 port map( A1 => n60400, A2 => n62040, B1 => n2845, B2 => 
                           n60398, ZN => n12330);
   U5157 : OAI22_X1 port map( A1 => n60400, A2 => n62054, B1 => n2844, B2 => 
                           n60398, ZN => n12331);
   U5158 : OAI22_X1 port map( A1 => n60400, A2 => n62068, B1 => n2843, B2 => 
                           n60398, ZN => n12332);
   U5159 : OAI22_X1 port map( A1 => n60400, A2 => n62082, B1 => n2842, B2 => 
                           n60398, ZN => n12333);
   U5160 : OAI22_X1 port map( A1 => n60400, A2 => n62096, B1 => n2841, B2 => 
                           n60398, ZN => n12334);
   U5161 : OAI22_X1 port map( A1 => n60401, A2 => n62110, B1 => n2840, B2 => 
                           n60398, ZN => n12335);
   U5162 : OAI22_X1 port map( A1 => n60401, A2 => n60963, B1 => n2839, B2 => 
                           n60398, ZN => n12336);
   U5163 : OAI22_X1 port map( A1 => n60401, A2 => n60977, B1 => n2790, B2 => 
                           n15185, ZN => n12337);
   U5164 : OAI22_X1 port map( A1 => n60401, A2 => n60991, B1 => n2789, B2 => 
                           n15185, ZN => n12338);
   U5165 : OAI22_X1 port map( A1 => n60401, A2 => n61005, B1 => n2788, B2 => 
                           n15185, ZN => n12339);
   U5166 : OAI22_X1 port map( A1 => n60402, A2 => n61019, B1 => n2787, B2 => 
                           n15185, ZN => n12340);
   U5167 : OAI22_X1 port map( A1 => n60402, A2 => n61033, B1 => n2786, B2 => 
                           n15185, ZN => n12341);
   U5168 : OAI22_X1 port map( A1 => n60402, A2 => n61047, B1 => n2785, B2 => 
                           n15185, ZN => n12342);
   U5169 : OAI22_X1 port map( A1 => n60402, A2 => n61061, B1 => n2784, B2 => 
                           n15185, ZN => n12343);
   U5170 : OAI22_X1 port map( A1 => n60402, A2 => n61075, B1 => n2783, B2 => 
                           n60398, ZN => n12344);
   U5171 : OAI22_X1 port map( A1 => n60403, A2 => n61089, B1 => n2782, B2 => 
                           n60398, ZN => n12345);
   U5172 : OAI22_X1 port map( A1 => n60403, A2 => n61103, B1 => n2781, B2 => 
                           n60398, ZN => n12346);
   U5173 : OAI22_X1 port map( A1 => n60403, A2 => n61117, B1 => n2780, B2 => 
                           n60398, ZN => n12347);
   U5174 : OAI22_X1 port map( A1 => n60403, A2 => n61131, B1 => n2779, B2 => 
                           n60398, ZN => n12348);
   U5175 : OAI22_X1 port map( A1 => n60939, A2 => n61965, B1 => n2778, B2 => 
                           n60938, ZN => n14245);
   U5176 : OAI22_X1 port map( A1 => n60939, A2 => n61979, B1 => n2777, B2 => 
                           n60938, ZN => n14246);
   U5177 : OAI22_X1 port map( A1 => n60939, A2 => n61993, B1 => n2776, B2 => 
                           n60938, ZN => n14247);
   U5178 : OAI22_X1 port map( A1 => n60939, A2 => n62007, B1 => n2775, B2 => 
                           n60938, ZN => n14248);
   U5179 : OAI22_X1 port map( A1 => n60939, A2 => n62021, B1 => n2774, B2 => 
                           n60938, ZN => n14249);
   U5180 : OAI22_X1 port map( A1 => n60940, A2 => n62035, B1 => n2773, B2 => 
                           n60938, ZN => n14250);
   U5181 : OAI22_X1 port map( A1 => n60940, A2 => n62049, B1 => n2772, B2 => 
                           n60938, ZN => n14251);
   U5182 : OAI22_X1 port map( A1 => n60940, A2 => n62063, B1 => n2771, B2 => 
                           n60938, ZN => n14252);
   U5183 : OAI22_X1 port map( A1 => n60940, A2 => n62077, B1 => n2770, B2 => 
                           n60938, ZN => n14253);
   U5184 : OAI22_X1 port map( A1 => n60930, A2 => n62007, B1 => n2769, B2 => 
                           n15100, ZN => n14216);
   U5185 : OAI22_X1 port map( A1 => n60930, A2 => n62021, B1 => n2768, B2 => 
                           n15100, ZN => n14217);
   U5186 : OAI22_X1 port map( A1 => n60931, A2 => n62035, B1 => n2767, B2 => 
                           n15100, ZN => n14218);
   U5187 : OAI22_X1 port map( A1 => n60931, A2 => n62049, B1 => n2766, B2 => 
                           n15100, ZN => n14219);
   U5188 : OAI22_X1 port map( A1 => n60931, A2 => n62063, B1 => n2765, B2 => 
                           n15100, ZN => n14220);
   U5189 : OAI22_X1 port map( A1 => n60931, A2 => n62077, B1 => n2764, B2 => 
                           n15100, ZN => n14221);
   U5190 : OAI22_X1 port map( A1 => n60931, A2 => n62091, B1 => n2763, B2 => 
                           n15100, ZN => n14222);
   U5191 : OAI22_X1 port map( A1 => n60932, A2 => n62105, B1 => n2762, B2 => 
                           n60929, ZN => n14223);
   U5192 : OAI22_X1 port map( A1 => n60932, A2 => n60958, B1 => n2761, B2 => 
                           n60929, ZN => n14224);
   U5193 : OAI22_X1 port map( A1 => n60932, A2 => n60972, B1 => n2760, B2 => 
                           n60929, ZN => n14225);
   U5194 : OAI22_X1 port map( A1 => n60932, A2 => n60986, B1 => n2759, B2 => 
                           n60929, ZN => n14226);
   U5195 : OAI22_X1 port map( A1 => n60932, A2 => n61000, B1 => n2758, B2 => 
                           n60929, ZN => n14227);
   U5196 : OAI22_X1 port map( A1 => n60933, A2 => n61014, B1 => n2757, B2 => 
                           n60929, ZN => n14228);
   U5197 : OAI22_X1 port map( A1 => n60933, A2 => n61028, B1 => n2756, B2 => 
                           n60929, ZN => n14229);
   U5198 : OAI22_X1 port map( A1 => n60933, A2 => n61042, B1 => n2755, B2 => 
                           n60929, ZN => n14230);
   U5199 : OAI22_X1 port map( A1 => n60933, A2 => n61056, B1 => n2754, B2 => 
                           n60929, ZN => n14231);
   U5200 : OAI22_X1 port map( A1 => n60933, A2 => n61070, B1 => n2753, B2 => 
                           n60929, ZN => n14232);
   U5201 : OAI22_X1 port map( A1 => n60934, A2 => n61084, B1 => n2752, B2 => 
                           n60929, ZN => n14233);
   U5202 : OAI22_X1 port map( A1 => n60934, A2 => n61098, B1 => n2751, B2 => 
                           n60929, ZN => n14234);
   U5203 : OAI22_X1 port map( A1 => n60934, A2 => n61112, B1 => n2750, B2 => 
                           n60929, ZN => n14235);
   U5204 : OAI22_X1 port map( A1 => n60934, A2 => n61126, B1 => n2749, B2 => 
                           n60929, ZN => n14236);
   U5205 : OAI22_X1 port map( A1 => n60372, A2 => n61970, B1 => n2724, B2 => 
                           n60371, ZN => n12229);
   U5206 : OAI22_X1 port map( A1 => n60372, A2 => n61984, B1 => n2723, B2 => 
                           n60371, ZN => n12230);
   U5207 : OAI22_X1 port map( A1 => n60372, A2 => n61998, B1 => n2722, B2 => 
                           n60371, ZN => n12231);
   U5208 : OAI22_X1 port map( A1 => n60372, A2 => n62012, B1 => n2721, B2 => 
                           n60371, ZN => n12232);
   U5209 : OAI22_X1 port map( A1 => n60372, A2 => n62026, B1 => n2720, B2 => 
                           n60371, ZN => n12233);
   U5210 : OAI22_X1 port map( A1 => n60373, A2 => n62040, B1 => n2719, B2 => 
                           n60371, ZN => n12234);
   U5211 : OAI22_X1 port map( A1 => n60373, A2 => n62054, B1 => n2718, B2 => 
                           n60371, ZN => n12235);
   U5212 : OAI22_X1 port map( A1 => n60373, A2 => n62068, B1 => n2717, B2 => 
                           n60371, ZN => n12236);
   U5213 : OAI22_X1 port map( A1 => n60373, A2 => n62082, B1 => n2716, B2 => 
                           n60371, ZN => n12237);
   U5214 : OAI22_X1 port map( A1 => n60373, A2 => n62096, B1 => n2715, B2 => 
                           n60371, ZN => n12238);
   U5215 : OAI22_X1 port map( A1 => n60374, A2 => n62110, B1 => n2714, B2 => 
                           n60371, ZN => n12239);
   U5216 : OAI22_X1 port map( A1 => n60374, A2 => n60963, B1 => n2713, B2 => 
                           n60371, ZN => n12240);
   U5217 : OAI22_X1 port map( A1 => n60374, A2 => n60977, B1 => n2712, B2 => 
                           n15189, ZN => n12241);
   U5218 : OAI22_X1 port map( A1 => n60374, A2 => n60991, B1 => n2711, B2 => 
                           n15189, ZN => n12242);
   U5219 : OAI22_X1 port map( A1 => n60374, A2 => n61005, B1 => n2710, B2 => 
                           n15189, ZN => n12243);
   U5220 : OAI22_X1 port map( A1 => n60375, A2 => n61019, B1 => n2709, B2 => 
                           n15189, ZN => n12244);
   U5221 : OAI22_X1 port map( A1 => n60375, A2 => n61033, B1 => n2708, B2 => 
                           n15189, ZN => n12245);
   U5222 : OAI22_X1 port map( A1 => n60375, A2 => n61047, B1 => n2707, B2 => 
                           n15189, ZN => n12246);
   U5223 : OAI22_X1 port map( A1 => n60375, A2 => n61061, B1 => n2706, B2 => 
                           n15189, ZN => n12247);
   U5224 : OAI22_X1 port map( A1 => n60375, A2 => n61075, B1 => n2705, B2 => 
                           n60371, ZN => n12248);
   U5225 : OAI22_X1 port map( A1 => n60376, A2 => n61089, B1 => n2704, B2 => 
                           n60371, ZN => n12249);
   U5226 : OAI22_X1 port map( A1 => n60376, A2 => n61103, B1 => n2703, B2 => 
                           n60371, ZN => n12250);
   U5227 : OAI22_X1 port map( A1 => n60376, A2 => n61117, B1 => n2702, B2 => 
                           n60371, ZN => n12251);
   U5228 : OAI22_X1 port map( A1 => n60376, A2 => n61131, B1 => n2701, B2 => 
                           n60371, ZN => n12252);
   U5229 : OAI22_X1 port map( A1 => n60365, A2 => n60977, B1 => n2688, B2 => 
                           n60362, ZN => n12209);
   U5230 : OAI22_X1 port map( A1 => n60365, A2 => n60991, B1 => n2687, B2 => 
                           n60362, ZN => n12210);
   U5231 : OAI22_X1 port map( A1 => n60365, A2 => n61005, B1 => n2686, B2 => 
                           n60362, ZN => n12211);
   U5232 : OAI22_X1 port map( A1 => n60366, A2 => n61019, B1 => n2685, B2 => 
                           n60362, ZN => n12212);
   U5233 : OAI22_X1 port map( A1 => n60366, A2 => n61033, B1 => n2684, B2 => 
                           n60362, ZN => n12213);
   U5234 : OAI22_X1 port map( A1 => n60366, A2 => n61047, B1 => n2683, B2 => 
                           n60362, ZN => n12214);
   U5235 : OAI22_X1 port map( A1 => n60366, A2 => n61061, B1 => n2682, B2 => 
                           n60362, ZN => n12215);
   U5236 : OAI22_X1 port map( A1 => n60366, A2 => n61075, B1 => n2681, B2 => 
                           n60362, ZN => n12216);
   U5237 : OAI22_X1 port map( A1 => n60367, A2 => n61089, B1 => n2680, B2 => 
                           n60362, ZN => n12217);
   U5238 : OAI22_X1 port map( A1 => n60367, A2 => n61103, B1 => n2679, B2 => 
                           n60362, ZN => n12218);
   U5239 : OAI22_X1 port map( A1 => n60367, A2 => n61117, B1 => n2678, B2 => 
                           n60362, ZN => n12219);
   U5240 : OAI22_X1 port map( A1 => n60367, A2 => n61131, B1 => n2677, B2 => 
                           n60362, ZN => n12220);
   U5241 : OAI22_X1 port map( A1 => n60345, A2 => n61970, B1 => n2652, B2 => 
                           n60344, ZN => n12133);
   U5242 : OAI22_X1 port map( A1 => n60345, A2 => n61984, B1 => n2644, B2 => 
                           n60344, ZN => n12134);
   U5243 : OAI22_X1 port map( A1 => n60345, A2 => n61998, B1 => n2643, B2 => 
                           n60344, ZN => n12135);
   U5244 : OAI22_X1 port map( A1 => n60345, A2 => n62012, B1 => n2642, B2 => 
                           n60344, ZN => n12136);
   U5245 : OAI22_X1 port map( A1 => n60345, A2 => n62026, B1 => n2641, B2 => 
                           n60344, ZN => n12137);
   U5246 : OAI22_X1 port map( A1 => n60346, A2 => n62040, B1 => n2640, B2 => 
                           n60344, ZN => n12138);
   U5247 : OAI22_X1 port map( A1 => n60346, A2 => n62054, B1 => n2639, B2 => 
                           n60344, ZN => n12139);
   U5248 : OAI22_X1 port map( A1 => n60346, A2 => n62068, B1 => n2638, B2 => 
                           n60344, ZN => n12140);
   U5249 : OAI22_X1 port map( A1 => n60346, A2 => n62082, B1 => n2637, B2 => 
                           n60344, ZN => n12141);
   U5250 : OAI22_X1 port map( A1 => n60346, A2 => n62096, B1 => n2636, B2 => 
                           n60344, ZN => n12142);
   U5251 : OAI22_X1 port map( A1 => n60347, A2 => n62110, B1 => n2635, B2 => 
                           n60344, ZN => n12143);
   U5252 : OAI22_X1 port map( A1 => n60347, A2 => n60963, B1 => n2634, B2 => 
                           n60344, ZN => n12144);
   U5253 : OAI22_X1 port map( A1 => n60347, A2 => n60977, B1 => n2633, B2 => 
                           n15192, ZN => n12145);
   U5254 : OAI22_X1 port map( A1 => n60347, A2 => n60991, B1 => n2632, B2 => 
                           n15192, ZN => n12146);
   U5255 : OAI22_X1 port map( A1 => n60347, A2 => n61005, B1 => n2631, B2 => 
                           n15192, ZN => n12147);
   U5256 : OAI22_X1 port map( A1 => n60348, A2 => n61019, B1 => n2630, B2 => 
                           n15192, ZN => n12148);
   U5257 : OAI22_X1 port map( A1 => n60348, A2 => n61033, B1 => n2629, B2 => 
                           n15192, ZN => n12149);
   U5258 : OAI22_X1 port map( A1 => n60348, A2 => n61047, B1 => n2628, B2 => 
                           n15192, ZN => n12150);
   U5259 : OAI22_X1 port map( A1 => n60348, A2 => n61061, B1 => n2627, B2 => 
                           n15192, ZN => n12151);
   U5260 : OAI22_X1 port map( A1 => n60348, A2 => n61075, B1 => n2626, B2 => 
                           n60344, ZN => n12152);
   U5261 : OAI22_X1 port map( A1 => n60349, A2 => n61089, B1 => n2625, B2 => 
                           n60344, ZN => n12153);
   U5262 : OAI22_X1 port map( A1 => n60349, A2 => n61103, B1 => n2624, B2 => 
                           n60344, ZN => n12154);
   U5263 : OAI22_X1 port map( A1 => n60349, A2 => n61117, B1 => n2623, B2 => 
                           n60344, ZN => n12155);
   U5264 : OAI22_X1 port map( A1 => n60349, A2 => n61131, B1 => n2622, B2 => 
                           n60344, ZN => n12156);
   U5265 : OAI22_X1 port map( A1 => n60336, A2 => n61970, B1 => n2621, B2 => 
                           n60335, ZN => n12101);
   U5266 : OAI22_X1 port map( A1 => n60336, A2 => n61984, B1 => n2620, B2 => 
                           n60335, ZN => n12102);
   U5267 : OAI22_X1 port map( A1 => n60336, A2 => n61998, B1 => n2619, B2 => 
                           n60335, ZN => n12103);
   U5268 : OAI22_X1 port map( A1 => n60336, A2 => n62012, B1 => n2618, B2 => 
                           n60335, ZN => n12104);
   U5269 : OAI22_X1 port map( A1 => n60336, A2 => n62026, B1 => n2617, B2 => 
                           n60335, ZN => n12105);
   U5270 : OAI22_X1 port map( A1 => n60337, A2 => n62040, B1 => n2616, B2 => 
                           n60335, ZN => n12106);
   U5271 : OAI22_X1 port map( A1 => n60337, A2 => n62054, B1 => n2615, B2 => 
                           n60335, ZN => n12107);
   U5272 : OAI22_X1 port map( A1 => n60337, A2 => n62068, B1 => n2614, B2 => 
                           n60335, ZN => n12108);
   U5273 : OAI22_X1 port map( A1 => n60337, A2 => n62082, B1 => n2613, B2 => 
                           n60335, ZN => n12109);
   U5274 : OAI22_X1 port map( A1 => n60337, A2 => n62096, B1 => n2612, B2 => 
                           n60335, ZN => n12110);
   U5275 : OAI22_X1 port map( A1 => n60338, A2 => n62110, B1 => n2611, B2 => 
                           n60335, ZN => n12111);
   U5276 : OAI22_X1 port map( A1 => n60338, A2 => n60963, B1 => n2610, B2 => 
                           n60335, ZN => n12112);
   U5277 : OAI22_X1 port map( A1 => n60338, A2 => n60977, B1 => n2609, B2 => 
                           n15193, ZN => n12113);
   U5278 : OAI22_X1 port map( A1 => n60338, A2 => n60991, B1 => n2608, B2 => 
                           n15193, ZN => n12114);
   U5279 : OAI22_X1 port map( A1 => n60338, A2 => n61005, B1 => n2607, B2 => 
                           n15193, ZN => n12115);
   U5280 : OAI22_X1 port map( A1 => n60339, A2 => n61019, B1 => n2606, B2 => 
                           n15193, ZN => n12116);
   U5281 : OAI22_X1 port map( A1 => n60339, A2 => n61033, B1 => n2605, B2 => 
                           n15193, ZN => n12117);
   U5282 : OAI22_X1 port map( A1 => n60339, A2 => n61047, B1 => n2604, B2 => 
                           n15193, ZN => n12118);
   U5283 : OAI22_X1 port map( A1 => n60339, A2 => n61061, B1 => n2603, B2 => 
                           n15193, ZN => n12119);
   U5284 : OAI22_X1 port map( A1 => n60339, A2 => n61075, B1 => n2602, B2 => 
                           n60335, ZN => n12120);
   U5285 : OAI22_X1 port map( A1 => n60340, A2 => n61089, B1 => n2601, B2 => 
                           n60335, ZN => n12121);
   U5286 : OAI22_X1 port map( A1 => n60340, A2 => n61103, B1 => n2600, B2 => 
                           n60335, ZN => n12122);
   U5287 : OAI22_X1 port map( A1 => n60340, A2 => n61117, B1 => n2599, B2 => 
                           n60335, ZN => n12123);
   U5288 : OAI22_X1 port map( A1 => n60340, A2 => n61131, B1 => n2598, B2 => 
                           n60335, ZN => n12124);
   U5289 : OAI22_X1 port map( A1 => n60309, A2 => n61971, B1 => n2549, B2 => 
                           n60308, ZN => n12005);
   U5290 : OAI22_X1 port map( A1 => n60309, A2 => n61985, B1 => n2548, B2 => 
                           n60308, ZN => n12006);
   U5291 : OAI22_X1 port map( A1 => n60309, A2 => n61999, B1 => n2547, B2 => 
                           n60308, ZN => n12007);
   U5292 : OAI22_X1 port map( A1 => n60309, A2 => n62013, B1 => n2546, B2 => 
                           n60308, ZN => n12008);
   U5293 : OAI22_X1 port map( A1 => n60309, A2 => n62027, B1 => n2545, B2 => 
                           n60308, ZN => n12009);
   U5294 : OAI22_X1 port map( A1 => n60310, A2 => n62041, B1 => n2544, B2 => 
                           n60308, ZN => n12010);
   U5295 : OAI22_X1 port map( A1 => n60310, A2 => n62055, B1 => n2543, B2 => 
                           n60308, ZN => n12011);
   U5296 : OAI22_X1 port map( A1 => n60310, A2 => n62069, B1 => n2542, B2 => 
                           n60308, ZN => n12012);
   U5297 : OAI22_X1 port map( A1 => n60310, A2 => n62083, B1 => n2541, B2 => 
                           n60308, ZN => n12013);
   U5298 : OAI22_X1 port map( A1 => n60310, A2 => n62097, B1 => n2540, B2 => 
                           n60308, ZN => n12014);
   U5299 : OAI22_X1 port map( A1 => n60311, A2 => n62111, B1 => n2539, B2 => 
                           n60308, ZN => n12015);
   U5300 : OAI22_X1 port map( A1 => n60311, A2 => n60964, B1 => n2538, B2 => 
                           n60308, ZN => n12016);
   U5301 : OAI22_X1 port map( A1 => n60311, A2 => n60978, B1 => n2537, B2 => 
                           n15196, ZN => n12017);
   U5302 : OAI22_X1 port map( A1 => n60311, A2 => n60992, B1 => n2536, B2 => 
                           n15196, ZN => n12018);
   U5303 : OAI22_X1 port map( A1 => n60311, A2 => n61006, B1 => n2535, B2 => 
                           n15196, ZN => n12019);
   U5304 : OAI22_X1 port map( A1 => n60312, A2 => n61020, B1 => n2534, B2 => 
                           n15196, ZN => n12020);
   U5305 : OAI22_X1 port map( A1 => n60312, A2 => n61034, B1 => n2533, B2 => 
                           n15196, ZN => n12021);
   U5306 : OAI22_X1 port map( A1 => n60312, A2 => n61048, B1 => n2532, B2 => 
                           n15196, ZN => n12022);
   U5307 : OAI22_X1 port map( A1 => n60312, A2 => n61062, B1 => n2531, B2 => 
                           n15196, ZN => n12023);
   U5308 : OAI22_X1 port map( A1 => n60312, A2 => n61076, B1 => n2530, B2 => 
                           n60308, ZN => n12024);
   U5309 : OAI22_X1 port map( A1 => n60313, A2 => n61090, B1 => n2529, B2 => 
                           n60308, ZN => n12025);
   U5310 : OAI22_X1 port map( A1 => n60313, A2 => n61104, B1 => n2528, B2 => 
                           n60308, ZN => n12026);
   U5311 : OAI22_X1 port map( A1 => n60313, A2 => n61118, B1 => n2527, B2 => 
                           n60308, ZN => n12027);
   U5312 : OAI22_X1 port map( A1 => n60313, A2 => n61132, B1 => n2526, B2 => 
                           n60308, ZN => n12028);
   U5313 : OAI22_X1 port map( A1 => n60300, A2 => n61971, B1 => n2525, B2 => 
                           n60299, ZN => n11973);
   U5314 : OAI22_X1 port map( A1 => n60300, A2 => n61985, B1 => n2524, B2 => 
                           n60299, ZN => n11974);
   U5315 : OAI22_X1 port map( A1 => n60300, A2 => n61999, B1 => n2523, B2 => 
                           n60299, ZN => n11975);
   U5316 : OAI22_X1 port map( A1 => n60300, A2 => n62013, B1 => n2522, B2 => 
                           n60299, ZN => n11976);
   U5317 : OAI22_X1 port map( A1 => n60300, A2 => n62027, B1 => n2521, B2 => 
                           n60299, ZN => n11977);
   U5318 : OAI22_X1 port map( A1 => n60301, A2 => n62041, B1 => n2520, B2 => 
                           n60299, ZN => n11978);
   U5319 : OAI22_X1 port map( A1 => n60301, A2 => n62055, B1 => n2519, B2 => 
                           n60299, ZN => n11979);
   U5320 : OAI22_X1 port map( A1 => n60301, A2 => n62069, B1 => n2518, B2 => 
                           n60299, ZN => n11980);
   U5321 : OAI22_X1 port map( A1 => n60301, A2 => n62083, B1 => n2517, B2 => 
                           n60299, ZN => n11981);
   U5322 : OAI22_X1 port map( A1 => n60301, A2 => n62097, B1 => n2516, B2 => 
                           n60299, ZN => n11982);
   U5323 : OAI22_X1 port map( A1 => n60302, A2 => n62111, B1 => n2515, B2 => 
                           n60299, ZN => n11983);
   U5324 : OAI22_X1 port map( A1 => n60302, A2 => n60964, B1 => n2514, B2 => 
                           n60299, ZN => n11984);
   U5325 : OAI22_X1 port map( A1 => n60302, A2 => n60978, B1 => n2513, B2 => 
                           n15197, ZN => n11985);
   U5326 : OAI22_X1 port map( A1 => n60302, A2 => n60992, B1 => n2512, B2 => 
                           n15197, ZN => n11986);
   U5327 : OAI22_X1 port map( A1 => n60302, A2 => n61006, B1 => n2511, B2 => 
                           n15197, ZN => n11987);
   U5328 : OAI22_X1 port map( A1 => n60303, A2 => n61020, B1 => n2482, B2 => 
                           n15197, ZN => n11988);
   U5329 : OAI22_X1 port map( A1 => n60303, A2 => n61034, B1 => n2481, B2 => 
                           n15197, ZN => n11989);
   U5330 : OAI22_X1 port map( A1 => n60303, A2 => n61048, B1 => n2480, B2 => 
                           n15197, ZN => n11990);
   U5331 : OAI22_X1 port map( A1 => n60303, A2 => n61062, B1 => n2479, B2 => 
                           n15197, ZN => n11991);
   U5332 : OAI22_X1 port map( A1 => n60303, A2 => n61076, B1 => n2478, B2 => 
                           n60299, ZN => n11992);
   U5333 : OAI22_X1 port map( A1 => n60304, A2 => n61090, B1 => n2477, B2 => 
                           n60299, ZN => n11993);
   U5334 : OAI22_X1 port map( A1 => n60304, A2 => n61104, B1 => n2476, B2 => 
                           n60299, ZN => n11994);
   U5335 : OAI22_X1 port map( A1 => n60304, A2 => n61118, B1 => n2475, B2 => 
                           n60299, ZN => n11995);
   U5336 : OAI22_X1 port map( A1 => n60304, A2 => n61132, B1 => n2474, B2 => 
                           n60299, ZN => n11996);
   U5337 : OAI22_X1 port map( A1 => n60273, A2 => n61971, B1 => n2401, B2 => 
                           n60272, ZN => n11877);
   U5338 : OAI22_X1 port map( A1 => n60273, A2 => n61985, B1 => n2400, B2 => 
                           n60272, ZN => n11878);
   U5339 : OAI22_X1 port map( A1 => n60273, A2 => n61999, B1 => n2399, B2 => 
                           n60272, ZN => n11879);
   U5340 : OAI22_X1 port map( A1 => n60273, A2 => n62013, B1 => n2398, B2 => 
                           n60272, ZN => n11880);
   U5341 : OAI22_X1 port map( A1 => n60273, A2 => n62027, B1 => n2397, B2 => 
                           n60272, ZN => n11881);
   U5342 : OAI22_X1 port map( A1 => n60274, A2 => n62041, B1 => n2396, B2 => 
                           n60272, ZN => n11882);
   U5343 : OAI22_X1 port map( A1 => n60274, A2 => n62055, B1 => n2395, B2 => 
                           n60272, ZN => n11883);
   U5344 : OAI22_X1 port map( A1 => n60274, A2 => n62069, B1 => n2394, B2 => 
                           n60272, ZN => n11884);
   U5345 : OAI22_X1 port map( A1 => n60274, A2 => n62083, B1 => n2393, B2 => 
                           n60272, ZN => n11885);
   U5346 : OAI22_X1 port map( A1 => n60274, A2 => n62097, B1 => n2392, B2 => 
                           n60272, ZN => n11886);
   U5347 : OAI22_X1 port map( A1 => n60275, A2 => n62111, B1 => n2391, B2 => 
                           n60272, ZN => n11887);
   U5348 : OAI22_X1 port map( A1 => n60275, A2 => n60964, B1 => n2298, B2 => 
                           n60272, ZN => n11888);
   U5349 : OAI22_X1 port map( A1 => n60275, A2 => n60978, B1 => n2297, B2 => 
                           n15200, ZN => n11889);
   U5350 : OAI22_X1 port map( A1 => n60275, A2 => n60992, B1 => n2296, B2 => 
                           n15200, ZN => n11890);
   U5351 : OAI22_X1 port map( A1 => n60275, A2 => n61006, B1 => n2295, B2 => 
                           n15200, ZN => n11891);
   U5352 : OAI22_X1 port map( A1 => n60276, A2 => n61020, B1 => n2294, B2 => 
                           n15200, ZN => n11892);
   U5353 : OAI22_X1 port map( A1 => n60276, A2 => n61034, B1 => n2293, B2 => 
                           n15200, ZN => n11893);
   U5354 : OAI22_X1 port map( A1 => n60276, A2 => n61048, B1 => n2292, B2 => 
                           n15200, ZN => n11894);
   U5355 : OAI22_X1 port map( A1 => n60276, A2 => n61062, B1 => n2291, B2 => 
                           n15200, ZN => n11895);
   U5356 : OAI22_X1 port map( A1 => n60276, A2 => n61076, B1 => n2290, B2 => 
                           n60272, ZN => n11896);
   U5357 : OAI22_X1 port map( A1 => n60277, A2 => n61090, B1 => n2289, B2 => 
                           n60272, ZN => n11897);
   U5358 : OAI22_X1 port map( A1 => n60277, A2 => n61104, B1 => n2288, B2 => 
                           n60272, ZN => n11898);
   U5359 : OAI22_X1 port map( A1 => n60277, A2 => n61118, B1 => n2287, B2 => 
                           n60272, ZN => n11899);
   U5360 : OAI22_X1 port map( A1 => n60277, A2 => n61132, B1 => n2286, B2 => 
                           n60272, ZN => n11900);
   U5361 : OAI22_X1 port map( A1 => n60264, A2 => n61971, B1 => n2285, B2 => 
                           n60263, ZN => n11845);
   U5362 : OAI22_X1 port map( A1 => n60264, A2 => n61985, B1 => n2284, B2 => 
                           n60263, ZN => n11846);
   U5363 : OAI22_X1 port map( A1 => n60264, A2 => n61999, B1 => n2283, B2 => 
                           n60263, ZN => n11847);
   U5364 : OAI22_X1 port map( A1 => n60264, A2 => n62013, B1 => n2282, B2 => 
                           n60263, ZN => n11848);
   U5365 : OAI22_X1 port map( A1 => n60264, A2 => n62027, B1 => n2281, B2 => 
                           n60263, ZN => n11849);
   U5366 : OAI22_X1 port map( A1 => n60265, A2 => n62041, B1 => n2280, B2 => 
                           n60263, ZN => n11850);
   U5367 : OAI22_X1 port map( A1 => n60265, A2 => n62055, B1 => n2279, B2 => 
                           n60263, ZN => n11851);
   U5368 : OAI22_X1 port map( A1 => n60265, A2 => n62069, B1 => n2278, B2 => 
                           n60263, ZN => n11852);
   U5369 : OAI22_X1 port map( A1 => n60265, A2 => n62083, B1 => n2277, B2 => 
                           n60263, ZN => n11853);
   U5370 : OAI22_X1 port map( A1 => n60265, A2 => n62097, B1 => n2276, B2 => 
                           n60263, ZN => n11854);
   U5371 : OAI22_X1 port map( A1 => n60266, A2 => n62111, B1 => n2275, B2 => 
                           n60263, ZN => n11855);
   U5372 : OAI22_X1 port map( A1 => n60266, A2 => n60964, B1 => n2274, B2 => 
                           n60263, ZN => n11856);
   U5373 : OAI22_X1 port map( A1 => n60266, A2 => n60978, B1 => n2273, B2 => 
                           n15201, ZN => n11857);
   U5374 : OAI22_X1 port map( A1 => n60266, A2 => n60992, B1 => n2272, B2 => 
                           n15201, ZN => n11858);
   U5375 : OAI22_X1 port map( A1 => n60266, A2 => n61006, B1 => n2271, B2 => 
                           n15201, ZN => n11859);
   U5376 : OAI22_X1 port map( A1 => n60267, A2 => n61020, B1 => n2234, B2 => 
                           n15201, ZN => n11860);
   U5377 : OAI22_X1 port map( A1 => n60267, A2 => n61034, B1 => n2233, B2 => 
                           n15201, ZN => n11861);
   U5378 : OAI22_X1 port map( A1 => n60267, A2 => n61048, B1 => n2232, B2 => 
                           n15201, ZN => n11862);
   U5379 : OAI22_X1 port map( A1 => n60267, A2 => n61062, B1 => n2231, B2 => 
                           n15201, ZN => n11863);
   U5380 : OAI22_X1 port map( A1 => n60267, A2 => n61076, B1 => n2230, B2 => 
                           n60263, ZN => n11864);
   U5381 : OAI22_X1 port map( A1 => n60268, A2 => n61090, B1 => n2229, B2 => 
                           n60263, ZN => n11865);
   U5382 : OAI22_X1 port map( A1 => n60268, A2 => n61104, B1 => n2228, B2 => 
                           n60263, ZN => n11866);
   U5383 : OAI22_X1 port map( A1 => n60268, A2 => n61118, B1 => n2227, B2 => 
                           n60263, ZN => n11867);
   U5384 : OAI22_X1 port map( A1 => n60268, A2 => n61132, B1 => n2226, B2 => 
                           n60263, ZN => n11868);
   U5385 : OAI22_X1 port map( A1 => n60237, A2 => n61971, B1 => n2169, B2 => 
                           n60236, ZN => n11749);
   U5386 : OAI22_X1 port map( A1 => n60237, A2 => n61985, B1 => n2168, B2 => 
                           n60236, ZN => n11750);
   U5387 : OAI22_X1 port map( A1 => n60237, A2 => n61999, B1 => n2167, B2 => 
                           n60236, ZN => n11751);
   U5388 : OAI22_X1 port map( A1 => n60237, A2 => n62013, B1 => n2166, B2 => 
                           n60236, ZN => n11752);
   U5389 : OAI22_X1 port map( A1 => n60237, A2 => n62027, B1 => n2165, B2 => 
                           n60236, ZN => n11753);
   U5390 : OAI22_X1 port map( A1 => n60238, A2 => n62041, B1 => n2164, B2 => 
                           n60236, ZN => n11754);
   U5391 : OAI22_X1 port map( A1 => n60238, A2 => n62055, B1 => n2163, B2 => 
                           n60236, ZN => n11755);
   U5392 : OAI22_X1 port map( A1 => n60238, A2 => n62069, B1 => n2162, B2 => 
                           n60236, ZN => n11756);
   U5393 : OAI22_X1 port map( A1 => n60238, A2 => n62083, B1 => n2161, B2 => 
                           n60236, ZN => n11757);
   U5394 : OAI22_X1 port map( A1 => n60238, A2 => n62097, B1 => n2160, B2 => 
                           n60236, ZN => n11758);
   U5395 : OAI22_X1 port map( A1 => n60239, A2 => n62111, B1 => n2159, B2 => 
                           n60236, ZN => n11759);
   U5396 : OAI22_X1 port map( A1 => n60239, A2 => n60964, B1 => n2158, B2 => 
                           n60236, ZN => n11760);
   U5397 : OAI22_X1 port map( A1 => n60239, A2 => n60978, B1 => n2157, B2 => 
                           n15212, ZN => n11761);
   U5398 : OAI22_X1 port map( A1 => n60239, A2 => n60992, B1 => n2156, B2 => 
                           n15212, ZN => n11762);
   U5399 : OAI22_X1 port map( A1 => n60239, A2 => n61006, B1 => n2155, B2 => 
                           n15212, ZN => n11763);
   U5400 : OAI22_X1 port map( A1 => n60240, A2 => n61020, B1 => n2154, B2 => 
                           n15212, ZN => n11764);
   U5401 : OAI22_X1 port map( A1 => n60240, A2 => n61034, B1 => n2153, B2 => 
                           n15212, ZN => n11765);
   U5402 : OAI22_X1 port map( A1 => n60240, A2 => n61048, B1 => n2152, B2 => 
                           n15212, ZN => n11766);
   U5403 : OAI22_X1 port map( A1 => n60240, A2 => n61062, B1 => n2151, B2 => 
                           n15212, ZN => n11767);
   U5404 : OAI22_X1 port map( A1 => n60240, A2 => n61076, B1 => n2150, B2 => 
                           n60236, ZN => n11768);
   U5405 : OAI22_X1 port map( A1 => n60241, A2 => n61090, B1 => n2149, B2 => 
                           n60236, ZN => n11769);
   U5406 : OAI22_X1 port map( A1 => n60241, A2 => n61104, B1 => n2148, B2 => 
                           n60236, ZN => n11770);
   U5407 : OAI22_X1 port map( A1 => n60241, A2 => n61118, B1 => n2147, B2 => 
                           n60236, ZN => n11771);
   U5408 : OAI22_X1 port map( A1 => n60241, A2 => n61132, B1 => n2146, B2 => 
                           n60236, ZN => n11772);
   U5409 : OAI22_X1 port map( A1 => n60228, A2 => n61971, B1 => n2145, B2 => 
                           n60227, ZN => n11717);
   U5410 : OAI22_X1 port map( A1 => n60228, A2 => n61985, B1 => n2144, B2 => 
                           n60227, ZN => n11718);
   U5411 : OAI22_X1 port map( A1 => n60228, A2 => n61999, B1 => n2143, B2 => 
                           n60227, ZN => n11719);
   U5412 : OAI22_X1 port map( A1 => n60228, A2 => n62013, B1 => n2142, B2 => 
                           n60227, ZN => n11720);
   U5413 : OAI22_X1 port map( A1 => n60228, A2 => n62027, B1 => n2141, B2 => 
                           n60227, ZN => n11721);
   U5414 : OAI22_X1 port map( A1 => n60229, A2 => n62041, B1 => n2140, B2 => 
                           n60227, ZN => n11722);
   U5415 : OAI22_X1 port map( A1 => n60229, A2 => n62055, B1 => n2139, B2 => 
                           n60227, ZN => n11723);
   U5416 : OAI22_X1 port map( A1 => n60229, A2 => n62069, B1 => n2138, B2 => 
                           n60227, ZN => n11724);
   U5417 : OAI22_X1 port map( A1 => n60229, A2 => n62083, B1 => n2137, B2 => 
                           n60227, ZN => n11725);
   U5418 : OAI22_X1 port map( A1 => n60229, A2 => n62097, B1 => n2136, B2 => 
                           n60227, ZN => n11726);
   U5419 : OAI22_X1 port map( A1 => n60230, A2 => n62111, B1 => n2135, B2 => 
                           n60227, ZN => n11727);
   U5420 : OAI22_X1 port map( A1 => n60230, A2 => n60964, B1 => n2134, B2 => 
                           n60227, ZN => n11728);
   U5421 : OAI22_X1 port map( A1 => n60230, A2 => n60978, B1 => n2133, B2 => 
                           n15214, ZN => n11729);
   U5422 : OAI22_X1 port map( A1 => n60230, A2 => n60992, B1 => n2132, B2 => 
                           n15214, ZN => n11730);
   U5423 : OAI22_X1 port map( A1 => n60230, A2 => n61006, B1 => n2131, B2 => 
                           n15214, ZN => n11731);
   U5424 : OAI22_X1 port map( A1 => n60231, A2 => n61020, B1 => n2130, B2 => 
                           n15214, ZN => n11732);
   U5425 : OAI22_X1 port map( A1 => n60231, A2 => n61034, B1 => n2129, B2 => 
                           n15214, ZN => n11733);
   U5426 : OAI22_X1 port map( A1 => n60231, A2 => n61048, B1 => n2128, B2 => 
                           n15214, ZN => n11734);
   U5427 : OAI22_X1 port map( A1 => n60231, A2 => n61062, B1 => n2127, B2 => 
                           n15214, ZN => n11735);
   U5428 : OAI22_X1 port map( A1 => n60231, A2 => n61076, B1 => n2126, B2 => 
                           n60227, ZN => n11736);
   U5429 : OAI22_X1 port map( A1 => n60232, A2 => n61090, B1 => n2125, B2 => 
                           n60227, ZN => n11737);
   U5430 : OAI22_X1 port map( A1 => n60232, A2 => n61104, B1 => n2124, B2 => 
                           n60227, ZN => n11738);
   U5431 : OAI22_X1 port map( A1 => n60232, A2 => n61118, B1 => n2123, B2 => 
                           n60227, ZN => n11739);
   U5432 : OAI22_X1 port map( A1 => n60232, A2 => n61132, B1 => n2122, B2 => 
                           n60227, ZN => n11740);
   U5433 : OAI22_X1 port map( A1 => n60210, A2 => n61971, B1 => n2097, B2 => 
                           n60209, ZN => n11653);
   U5434 : OAI22_X1 port map( A1 => n60210, A2 => n61985, B1 => n2096, B2 => 
                           n60209, ZN => n11654);
   U5435 : OAI22_X1 port map( A1 => n60210, A2 => n61999, B1 => n2095, B2 => 
                           n60209, ZN => n11655);
   U5436 : OAI22_X1 port map( A1 => n60210, A2 => n62013, B1 => n2094, B2 => 
                           n60209, ZN => n11656);
   U5437 : OAI22_X1 port map( A1 => n60210, A2 => n62027, B1 => n2093, B2 => 
                           n60209, ZN => n11657);
   U5438 : OAI22_X1 port map( A1 => n60211, A2 => n62041, B1 => n2092, B2 => 
                           n60209, ZN => n11658);
   U5439 : OAI22_X1 port map( A1 => n60211, A2 => n62055, B1 => n2091, B2 => 
                           n60209, ZN => n11659);
   U5440 : OAI22_X1 port map( A1 => n60211, A2 => n62069, B1 => n2090, B2 => 
                           n60209, ZN => n11660);
   U5441 : OAI22_X1 port map( A1 => n60211, A2 => n62083, B1 => n2089, B2 => 
                           n60209, ZN => n11661);
   U5442 : OAI22_X1 port map( A1 => n60211, A2 => n62097, B1 => n2088, B2 => 
                           n60209, ZN => n11662);
   U5443 : OAI22_X1 port map( A1 => n60212, A2 => n62111, B1 => n2087, B2 => 
                           n60209, ZN => n11663);
   U5444 : OAI22_X1 port map( A1 => n60212, A2 => n60964, B1 => n2086, B2 => 
                           n60209, ZN => n11664);
   U5445 : OAI22_X1 port map( A1 => n60212, A2 => n60978, B1 => n2085, B2 => 
                           n15216, ZN => n11665);
   U5446 : OAI22_X1 port map( A1 => n60212, A2 => n60992, B1 => n2084, B2 => 
                           n15216, ZN => n11666);
   U5447 : OAI22_X1 port map( A1 => n60212, A2 => n61006, B1 => n2083, B2 => 
                           n15216, ZN => n11667);
   U5448 : OAI22_X1 port map( A1 => n60213, A2 => n61020, B1 => n2082, B2 => 
                           n15216, ZN => n11668);
   U5449 : OAI22_X1 port map( A1 => n60213, A2 => n61034, B1 => n2081, B2 => 
                           n15216, ZN => n11669);
   U5450 : OAI22_X1 port map( A1 => n60213, A2 => n61048, B1 => n2080, B2 => 
                           n15216, ZN => n11670);
   U5451 : OAI22_X1 port map( A1 => n60213, A2 => n61062, B1 => n2079, B2 => 
                           n15216, ZN => n11671);
   U5452 : OAI22_X1 port map( A1 => n60213, A2 => n61076, B1 => n2074, B2 => 
                           n60209, ZN => n11672);
   U5453 : OAI22_X1 port map( A1 => n60214, A2 => n61090, B1 => n2073, B2 => 
                           n60209, ZN => n11673);
   U5454 : OAI22_X1 port map( A1 => n60214, A2 => n61104, B1 => n2072, B2 => 
                           n60209, ZN => n11674);
   U5455 : OAI22_X1 port map( A1 => n60214, A2 => n61118, B1 => n2071, B2 => 
                           n60209, ZN => n11675);
   U5456 : OAI22_X1 port map( A1 => n60214, A2 => n61132, B1 => n2070, B2 => 
                           n60209, ZN => n11676);
   U5457 : OAI22_X1 port map( A1 => n60192, A2 => n61972, B1 => n2045, B2 => 
                           n60191, ZN => n11589);
   U5458 : OAI22_X1 port map( A1 => n60192, A2 => n61986, B1 => n2044, B2 => 
                           n60191, ZN => n11590);
   U5459 : OAI22_X1 port map( A1 => n60192, A2 => n62000, B1 => n2043, B2 => 
                           n60191, ZN => n11591);
   U5460 : OAI22_X1 port map( A1 => n60192, A2 => n62014, B1 => n2042, B2 => 
                           n60191, ZN => n11592);
   U5461 : OAI22_X1 port map( A1 => n60192, A2 => n62028, B1 => n2041, B2 => 
                           n60191, ZN => n11593);
   U5462 : OAI22_X1 port map( A1 => n60193, A2 => n62042, B1 => n2040, B2 => 
                           n60191, ZN => n11594);
   U5463 : OAI22_X1 port map( A1 => n60193, A2 => n62056, B1 => n2039, B2 => 
                           n60191, ZN => n11595);
   U5464 : OAI22_X1 port map( A1 => n60193, A2 => n62070, B1 => n2038, B2 => 
                           n60191, ZN => n11596);
   U5465 : OAI22_X1 port map( A1 => n60193, A2 => n62084, B1 => n2037, B2 => 
                           n60191, ZN => n11597);
   U5466 : OAI22_X1 port map( A1 => n60193, A2 => n62098, B1 => n2036, B2 => 
                           n60191, ZN => n11598);
   U5467 : OAI22_X1 port map( A1 => n60194, A2 => n62112, B1 => n2035, B2 => 
                           n60191, ZN => n11599);
   U5468 : OAI22_X1 port map( A1 => n60194, A2 => n60965, B1 => n2034, B2 => 
                           n60191, ZN => n11600);
   U5469 : OAI22_X1 port map( A1 => n60194, A2 => n60979, B1 => n2033, B2 => 
                           n15218, ZN => n11601);
   U5470 : OAI22_X1 port map( A1 => n60194, A2 => n60993, B1 => n2032, B2 => 
                           n15218, ZN => n11602);
   U5471 : OAI22_X1 port map( A1 => n60194, A2 => n61007, B1 => n2031, B2 => 
                           n15218, ZN => n11603);
   U5472 : OAI22_X1 port map( A1 => n60195, A2 => n61021, B1 => n2030, B2 => 
                           n15218, ZN => n11604);
   U5473 : OAI22_X1 port map( A1 => n60195, A2 => n61035, B1 => n2029, B2 => 
                           n15218, ZN => n11605);
   U5474 : OAI22_X1 port map( A1 => n60195, A2 => n61049, B1 => n2028, B2 => 
                           n15218, ZN => n11606);
   U5475 : OAI22_X1 port map( A1 => n60195, A2 => n61063, B1 => n2027, B2 => 
                           n15218, ZN => n11607);
   U5476 : OAI22_X1 port map( A1 => n60195, A2 => n61077, B1 => n2026, B2 => 
                           n60191, ZN => n11608);
   U5477 : OAI22_X1 port map( A1 => n60196, A2 => n61091, B1 => n2025, B2 => 
                           n60191, ZN => n11609);
   U5478 : OAI22_X1 port map( A1 => n60196, A2 => n61105, B1 => n2024, B2 => 
                           n60191, ZN => n11610);
   U5479 : OAI22_X1 port map( A1 => n60196, A2 => n61119, B1 => n2023, B2 => 
                           n60191, ZN => n11611);
   U5480 : OAI22_X1 port map( A1 => n60196, A2 => n61133, B1 => n1998, B2 => 
                           n60191, ZN => n11612);
   U5481 : OAI22_X1 port map( A1 => n60183, A2 => n61972, B1 => n1997, B2 => 
                           n60182, ZN => n11557);
   U5482 : OAI22_X1 port map( A1 => n60183, A2 => n61986, B1 => n1996, B2 => 
                           n60182, ZN => n11558);
   U5483 : OAI22_X1 port map( A1 => n60183, A2 => n62000, B1 => n1995, B2 => 
                           n60182, ZN => n11559);
   U5484 : OAI22_X1 port map( A1 => n60183, A2 => n62014, B1 => n1994, B2 => 
                           n60182, ZN => n11560);
   U5485 : OAI22_X1 port map( A1 => n60183, A2 => n62028, B1 => n1993, B2 => 
                           n60182, ZN => n11561);
   U5486 : OAI22_X1 port map( A1 => n60184, A2 => n62042, B1 => n1992, B2 => 
                           n60182, ZN => n11562);
   U5487 : OAI22_X1 port map( A1 => n60184, A2 => n62056, B1 => n1991, B2 => 
                           n60182, ZN => n11563);
   U5488 : OAI22_X1 port map( A1 => n60184, A2 => n62070, B1 => n1990, B2 => 
                           n60182, ZN => n11564);
   U5489 : OAI22_X1 port map( A1 => n60184, A2 => n62084, B1 => n1989, B2 => 
                           n60182, ZN => n11565);
   U5490 : OAI22_X1 port map( A1 => n60184, A2 => n62098, B1 => n1988, B2 => 
                           n60182, ZN => n11566);
   U5491 : OAI22_X1 port map( A1 => n60185, A2 => n62112, B1 => n1987, B2 => 
                           n60182, ZN => n11567);
   U5492 : OAI22_X1 port map( A1 => n60185, A2 => n60965, B1 => n1986, B2 => 
                           n60182, ZN => n11568);
   U5493 : OAI22_X1 port map( A1 => n60185, A2 => n60979, B1 => n1985, B2 => 
                           n15219, ZN => n11569);
   U5494 : OAI22_X1 port map( A1 => n60185, A2 => n60993, B1 => n1984, B2 => 
                           n15219, ZN => n11570);
   U5495 : OAI22_X1 port map( A1 => n60185, A2 => n61007, B1 => n1983, B2 => 
                           n15219, ZN => n11571);
   U5496 : OAI22_X1 port map( A1 => n60186, A2 => n61021, B1 => n1982, B2 => 
                           n15219, ZN => n11572);
   U5497 : OAI22_X1 port map( A1 => n60186, A2 => n61035, B1 => n1981, B2 => 
                           n15219, ZN => n11573);
   U5498 : OAI22_X1 port map( A1 => n60186, A2 => n61049, B1 => n1980, B2 => 
                           n15219, ZN => n11574);
   U5499 : OAI22_X1 port map( A1 => n60186, A2 => n61063, B1 => n1979, B2 => 
                           n15219, ZN => n11575);
   U5500 : OAI22_X1 port map( A1 => n60186, A2 => n61077, B1 => n1978, B2 => 
                           n60182, ZN => n11576);
   U5501 : OAI22_X1 port map( A1 => n60187, A2 => n61091, B1 => n1977, B2 => 
                           n60182, ZN => n11577);
   U5502 : OAI22_X1 port map( A1 => n60187, A2 => n61105, B1 => n1976, B2 => 
                           n60182, ZN => n11578);
   U5503 : OAI22_X1 port map( A1 => n60187, A2 => n61119, B1 => n1975, B2 => 
                           n60182, ZN => n11579);
   U5504 : OAI22_X1 port map( A1 => n60187, A2 => n61133, B1 => n1974, B2 => 
                           n60182, ZN => n11580);
   U5505 : OAI22_X1 port map( A1 => n60156, A2 => n61972, B1 => n1949, B2 => 
                           n60155, ZN => n11461);
   U5506 : OAI22_X1 port map( A1 => n60156, A2 => n61986, B1 => n1948, B2 => 
                           n60155, ZN => n11462);
   U5507 : OAI22_X1 port map( A1 => n60156, A2 => n62000, B1 => n1947, B2 => 
                           n60155, ZN => n11463);
   U5508 : OAI22_X1 port map( A1 => n60156, A2 => n62014, B1 => n1946, B2 => 
                           n60155, ZN => n11464);
   U5509 : OAI22_X1 port map( A1 => n60156, A2 => n62028, B1 => n1945, B2 => 
                           n60155, ZN => n11465);
   U5510 : OAI22_X1 port map( A1 => n60157, A2 => n62042, B1 => n1944, B2 => 
                           n60155, ZN => n11466);
   U5511 : OAI22_X1 port map( A1 => n60157, A2 => n62056, B1 => n1943, B2 => 
                           n60155, ZN => n11467);
   U5512 : OAI22_X1 port map( A1 => n60157, A2 => n62070, B1 => n1942, B2 => 
                           n60155, ZN => n11468);
   U5513 : OAI22_X1 port map( A1 => n60157, A2 => n62084, B1 => n1941, B2 => 
                           n60155, ZN => n11469);
   U5514 : OAI22_X1 port map( A1 => n60157, A2 => n62098, B1 => n1940, B2 => 
                           n60155, ZN => n11470);
   U5515 : OAI22_X1 port map( A1 => n60158, A2 => n62112, B1 => n1939, B2 => 
                           n60155, ZN => n11471);
   U5516 : OAI22_X1 port map( A1 => n60158, A2 => n60965, B1 => n1938, B2 => 
                           n60155, ZN => n11472);
   U5517 : OAI22_X1 port map( A1 => n60158, A2 => n60979, B1 => n1937, B2 => 
                           n15222, ZN => n11473);
   U5518 : OAI22_X1 port map( A1 => n60158, A2 => n60993, B1 => n1936, B2 => 
                           n15222, ZN => n11474);
   U5519 : OAI22_X1 port map( A1 => n60158, A2 => n61007, B1 => n1935, B2 => 
                           n15222, ZN => n11475);
   U5520 : OAI22_X1 port map( A1 => n60159, A2 => n61021, B1 => n1934, B2 => 
                           n15222, ZN => n11476);
   U5521 : OAI22_X1 port map( A1 => n60159, A2 => n61035, B1 => n1933, B2 => 
                           n15222, ZN => n11477);
   U5522 : OAI22_X1 port map( A1 => n60159, A2 => n61049, B1 => n1932, B2 => 
                           n15222, ZN => n11478);
   U5523 : OAI22_X1 port map( A1 => n60159, A2 => n61063, B1 => n1931, B2 => 
                           n15222, ZN => n11479);
   U5524 : OAI22_X1 port map( A1 => n60159, A2 => n61077, B1 => n1930, B2 => 
                           n60155, ZN => n11480);
   U5525 : OAI22_X1 port map( A1 => n60160, A2 => n61091, B1 => n1929, B2 => 
                           n60155, ZN => n11481);
   U5526 : OAI22_X1 port map( A1 => n60160, A2 => n61105, B1 => n1928, B2 => 
                           n60155, ZN => n11482);
   U5527 : OAI22_X1 port map( A1 => n60160, A2 => n61119, B1 => n1927, B2 => 
                           n60155, ZN => n11483);
   U5528 : OAI22_X1 port map( A1 => n60160, A2 => n61133, B1 => n1926, B2 => 
                           n60155, ZN => n11484);
   U5529 : OAI22_X1 port map( A1 => n60147, A2 => n61972, B1 => n1925, B2 => 
                           n60146, ZN => n11429);
   U5530 : OAI22_X1 port map( A1 => n60147, A2 => n61986, B1 => n1924, B2 => 
                           n60146, ZN => n11430);
   U5531 : OAI22_X1 port map( A1 => n60147, A2 => n62000, B1 => n1923, B2 => 
                           n60146, ZN => n11431);
   U5532 : OAI22_X1 port map( A1 => n60147, A2 => n62014, B1 => n1922, B2 => 
                           n60146, ZN => n11432);
   U5533 : OAI22_X1 port map( A1 => n60147, A2 => n62028, B1 => n1921, B2 => 
                           n60146, ZN => n11433);
   U5534 : OAI22_X1 port map( A1 => n60148, A2 => n62042, B1 => n1920, B2 => 
                           n60146, ZN => n11434);
   U5535 : OAI22_X1 port map( A1 => n60148, A2 => n62056, B1 => n1919, B2 => 
                           n60146, ZN => n11435);
   U5536 : OAI22_X1 port map( A1 => n60148, A2 => n62070, B1 => n1918, B2 => 
                           n60146, ZN => n11436);
   U5537 : OAI22_X1 port map( A1 => n60148, A2 => n62084, B1 => n1917, B2 => 
                           n60146, ZN => n11437);
   U5538 : OAI22_X1 port map( A1 => n60148, A2 => n62098, B1 => n1916, B2 => 
                           n60146, ZN => n11438);
   U5539 : OAI22_X1 port map( A1 => n60149, A2 => n62112, B1 => n1915, B2 => 
                           n60146, ZN => n11439);
   U5540 : OAI22_X1 port map( A1 => n60149, A2 => n60965, B1 => n1914, B2 => 
                           n60146, ZN => n11440);
   U5541 : OAI22_X1 port map( A1 => n60149, A2 => n60979, B1 => n1913, B2 => 
                           n15223, ZN => n11441);
   U5542 : OAI22_X1 port map( A1 => n60149, A2 => n60993, B1 => n1912, B2 => 
                           n15223, ZN => n11442);
   U5543 : OAI22_X1 port map( A1 => n60149, A2 => n61007, B1 => n1911, B2 => 
                           n15223, ZN => n11443);
   U5544 : OAI22_X1 port map( A1 => n60150, A2 => n61021, B1 => n1910, B2 => 
                           n15223, ZN => n11444);
   U5545 : OAI22_X1 port map( A1 => n60150, A2 => n61035, B1 => n1909, B2 => 
                           n15223, ZN => n11445);
   U5546 : OAI22_X1 port map( A1 => n60150, A2 => n61049, B1 => n1908, B2 => 
                           n15223, ZN => n11446);
   U5547 : OAI22_X1 port map( A1 => n60150, A2 => n61063, B1 => n1907, B2 => 
                           n15223, ZN => n11447);
   U5548 : OAI22_X1 port map( A1 => n60150, A2 => n61077, B1 => n1906, B2 => 
                           n60146, ZN => n11448);
   U5549 : OAI22_X1 port map( A1 => n60151, A2 => n61091, B1 => n1905, B2 => 
                           n60146, ZN => n11449);
   U5550 : OAI22_X1 port map( A1 => n60151, A2 => n61105, B1 => n1904, B2 => 
                           n60146, ZN => n11450);
   U5551 : OAI22_X1 port map( A1 => n60151, A2 => n61119, B1 => n1903, B2 => 
                           n60146, ZN => n11451);
   U5552 : OAI22_X1 port map( A1 => n60151, A2 => n61133, B1 => n1902, B2 => 
                           n60146, ZN => n11452);
   U5553 : OAI22_X1 port map( A1 => n60121, A2 => n62042, B1 => n1848, B2 => 
                           n15226, ZN => n11338);
   U5554 : OAI22_X1 port map( A1 => n60121, A2 => n62056, B1 => n1847, B2 => 
                           n15226, ZN => n11339);
   U5555 : OAI22_X1 port map( A1 => n60121, A2 => n62070, B1 => n1846, B2 => 
                           n15226, ZN => n11340);
   U5556 : OAI22_X1 port map( A1 => n60121, A2 => n62084, B1 => n1845, B2 => 
                           n15226, ZN => n11341);
   U5557 : OAI22_X1 port map( A1 => n60121, A2 => n62098, B1 => n1844, B2 => 
                           n15226, ZN => n11342);
   U5558 : OAI22_X1 port map( A1 => n60122, A2 => n62112, B1 => n1843, B2 => 
                           n15226, ZN => n11343);
   U5559 : OAI22_X1 port map( A1 => n60122, A2 => n60965, B1 => n1842, B2 => 
                           n15226, ZN => n11344);
   U5560 : OAI22_X1 port map( A1 => n60122, A2 => n60979, B1 => n1841, B2 => 
                           n60119, ZN => n11345);
   U5561 : OAI22_X1 port map( A1 => n60122, A2 => n60993, B1 => n1840, B2 => 
                           n60119, ZN => n11346);
   U5562 : OAI22_X1 port map( A1 => n60122, A2 => n61007, B1 => n1839, B2 => 
                           n60119, ZN => n11347);
   U5563 : OAI22_X1 port map( A1 => n60123, A2 => n61021, B1 => n1838, B2 => 
                           n60119, ZN => n11348);
   U5564 : OAI22_X1 port map( A1 => n60123, A2 => n61035, B1 => n1837, B2 => 
                           n60119, ZN => n11349);
   U5565 : OAI22_X1 port map( A1 => n60123, A2 => n61049, B1 => n1836, B2 => 
                           n60119, ZN => n11350);
   U5566 : OAI22_X1 port map( A1 => n60123, A2 => n61063, B1 => n1835, B2 => 
                           n60119, ZN => n11351);
   U5567 : OAI22_X1 port map( A1 => n60123, A2 => n61077, B1 => n1834, B2 => 
                           n60119, ZN => n11352);
   U5568 : OAI22_X1 port map( A1 => n60124, A2 => n61091, B1 => n1833, B2 => 
                           n60119, ZN => n11353);
   U5569 : OAI22_X1 port map( A1 => n60124, A2 => n61105, B1 => n1832, B2 => 
                           n60119, ZN => n11354);
   U5570 : OAI22_X1 port map( A1 => n60124, A2 => n61119, B1 => n1831, B2 => 
                           n60119, ZN => n11355);
   U5571 : OAI22_X1 port map( A1 => n60124, A2 => n61133, B1 => n1830, B2 => 
                           n60119, ZN => n11356);
   U5572 : OAI22_X1 port map( A1 => n60111, A2 => n61972, B1 => n1829, B2 => 
                           n60110, ZN => n11301);
   U5573 : OAI22_X1 port map( A1 => n60111, A2 => n61986, B1 => n1828, B2 => 
                           n60110, ZN => n11302);
   U5574 : OAI22_X1 port map( A1 => n60111, A2 => n62000, B1 => n1827, B2 => 
                           n60110, ZN => n11303);
   U5575 : OAI22_X1 port map( A1 => n60111, A2 => n62014, B1 => n1826, B2 => 
                           n60110, ZN => n11304);
   U5576 : OAI22_X1 port map( A1 => n60111, A2 => n62028, B1 => n1825, B2 => 
                           n60110, ZN => n11305);
   U5577 : OAI22_X1 port map( A1 => n60112, A2 => n62042, B1 => n1824, B2 => 
                           n60110, ZN => n11306);
   U5578 : OAI22_X1 port map( A1 => n60112, A2 => n62056, B1 => n1823, B2 => 
                           n60110, ZN => n11307);
   U5579 : OAI22_X1 port map( A1 => n60112, A2 => n62070, B1 => n1822, B2 => 
                           n60110, ZN => n11308);
   U5580 : OAI22_X1 port map( A1 => n60112, A2 => n62084, B1 => n1821, B2 => 
                           n60110, ZN => n11309);
   U5581 : OAI22_X1 port map( A1 => n60112, A2 => n62098, B1 => n1820, B2 => 
                           n60110, ZN => n11310);
   U5582 : OAI22_X1 port map( A1 => n60113, A2 => n62112, B1 => n1819, B2 => 
                           n60110, ZN => n11311);
   U5583 : OAI22_X1 port map( A1 => n60113, A2 => n60965, B1 => n1818, B2 => 
                           n60110, ZN => n11312);
   U5584 : OAI22_X1 port map( A1 => n60113, A2 => n60979, B1 => n1817, B2 => 
                           n15227, ZN => n11313);
   U5585 : OAI22_X1 port map( A1 => n60113, A2 => n60993, B1 => n1816, B2 => 
                           n15227, ZN => n11314);
   U5586 : OAI22_X1 port map( A1 => n60113, A2 => n61007, B1 => n1815, B2 => 
                           n15227, ZN => n11315);
   U5587 : OAI22_X1 port map( A1 => n60114, A2 => n61021, B1 => n1814, B2 => 
                           n15227, ZN => n11316);
   U5588 : OAI22_X1 port map( A1 => n60114, A2 => n61035, B1 => n1813, B2 => 
                           n15227, ZN => n11317);
   U5589 : OAI22_X1 port map( A1 => n60103, A2 => n62042, B1 => n1805, B2 => 
                           n60101, ZN => n11274);
   U5590 : OAI22_X1 port map( A1 => n60103, A2 => n62056, B1 => n1804, B2 => 
                           n60101, ZN => n11275);
   U5591 : OAI22_X1 port map( A1 => n60103, A2 => n62070, B1 => n1803, B2 => 
                           n60101, ZN => n11276);
   U5592 : OAI22_X1 port map( A1 => n60103, A2 => n62084, B1 => n1802, B2 => 
                           n60101, ZN => n11277);
   U5593 : OAI22_X1 port map( A1 => n60103, A2 => n62098, B1 => n1801, B2 => 
                           n60101, ZN => n11278);
   U5594 : OAI22_X1 port map( A1 => n60104, A2 => n62112, B1 => n1800, B2 => 
                           n60101, ZN => n11279);
   U5595 : OAI22_X1 port map( A1 => n60104, A2 => n60965, B1 => n1799, B2 => 
                           n60101, ZN => n11280);
   U5596 : OAI22_X1 port map( A1 => n60104, A2 => n60979, B1 => n1798, B2 => 
                           n15228, ZN => n11281);
   U5597 : OAI22_X1 port map( A1 => n60104, A2 => n60993, B1 => n1797, B2 => 
                           n15228, ZN => n11282);
   U5598 : OAI22_X1 port map( A1 => n60104, A2 => n61007, B1 => n1796, B2 => 
                           n15228, ZN => n11283);
   U5599 : OAI22_X1 port map( A1 => n60105, A2 => n61021, B1 => n1795, B2 => 
                           n15228, ZN => n11284);
   U5600 : OAI22_X1 port map( A1 => n60105, A2 => n61035, B1 => n1794, B2 => 
                           n15228, ZN => n11285);
   U5601 : OAI22_X1 port map( A1 => n60105, A2 => n61049, B1 => n1793, B2 => 
                           n15228, ZN => n11286);
   U5602 : OAI22_X1 port map( A1 => n60105, A2 => n61063, B1 => n1792, B2 => 
                           n15228, ZN => n11287);
   U5603 : OAI22_X1 port map( A1 => n60105, A2 => n61077, B1 => n1791, B2 => 
                           n60101, ZN => n11288);
   U5604 : OAI22_X1 port map( A1 => n60106, A2 => n61091, B1 => n1790, B2 => 
                           n60101, ZN => n11289);
   U5605 : OAI22_X1 port map( A1 => n60106, A2 => n61105, B1 => n1789, B2 => 
                           n60101, ZN => n11290);
   U5606 : OAI22_X1 port map( A1 => n60106, A2 => n61119, B1 => n1788, B2 => 
                           n60101, ZN => n11291);
   U5607 : OAI22_X1 port map( A1 => n60106, A2 => n61133, B1 => n1787, B2 => 
                           n60101, ZN => n11292);
   U5608 : OAI22_X1 port map( A1 => n60770, A2 => n61001, B1 => n1738, B2 => 
                           n15134, ZN => n13651);
   U5609 : OAI22_X1 port map( A1 => n60771, A2 => n61015, B1 => n1737, B2 => 
                           n15134, ZN => n13652);
   U5610 : OAI22_X1 port map( A1 => n60771, A2 => n61029, B1 => n1736, B2 => 
                           n15134, ZN => n13653);
   U5611 : OAI22_X1 port map( A1 => n60771, A2 => n61043, B1 => n1735, B2 => 
                           n15134, ZN => n13654);
   U5612 : OAI22_X1 port map( A1 => n60771, A2 => n61057, B1 => n1734, B2 => 
                           n15134, ZN => n13655);
   U5613 : OAI22_X1 port map( A1 => n60771, A2 => n61071, B1 => n1733, B2 => 
                           n15134, ZN => n13656);
   U5614 : OAI22_X1 port map( A1 => n60772, A2 => n61085, B1 => n1732, B2 => 
                           n15134, ZN => n13657);
   U5615 : OAI22_X1 port map( A1 => n60772, A2 => n61099, B1 => n1731, B2 => 
                           n60767, ZN => n13658);
   U5616 : OAI22_X1 port map( A1 => n60772, A2 => n61113, B1 => n1730, B2 => 
                           n60767, ZN => n13659);
   U5617 : OAI22_X1 port map( A1 => n60772, A2 => n61127, B1 => n1729, B2 => 
                           n60767, ZN => n13660);
   U5618 : OAI22_X1 port map( A1 => n60759, A2 => n61966, B1 => n1728, B2 => 
                           n60758, ZN => n13605);
   U5619 : OAI22_X1 port map( A1 => n60759, A2 => n61980, B1 => n1727, B2 => 
                           n60758, ZN => n13606);
   U5620 : OAI22_X1 port map( A1 => n60759, A2 => n61994, B1 => n1726, B2 => 
                           n60758, ZN => n13607);
   U5621 : OAI22_X1 port map( A1 => n60759, A2 => n62008, B1 => n1725, B2 => 
                           n60758, ZN => n13608);
   U5622 : OAI22_X1 port map( A1 => n60759, A2 => n62022, B1 => n1724, B2 => 
                           n60758, ZN => n13609);
   U5623 : OAI22_X1 port map( A1 => n60760, A2 => n62036, B1 => n1723, B2 => 
                           n60758, ZN => n13610);
   U5624 : OAI22_X1 port map( A1 => n60760, A2 => n62050, B1 => n1722, B2 => 
                           n60758, ZN => n13611);
   U5625 : OAI22_X1 port map( A1 => n60760, A2 => n62064, B1 => n1721, B2 => 
                           n60758, ZN => n13612);
   U5626 : OAI22_X1 port map( A1 => n60760, A2 => n62078, B1 => n1720, B2 => 
                           n60758, ZN => n13613);
   U5627 : OAI22_X1 port map( A1 => n60760, A2 => n62092, B1 => n1719, B2 => 
                           n60758, ZN => n13614);
   U5628 : OAI22_X1 port map( A1 => n60761, A2 => n62106, B1 => n1718, B2 => 
                           n60758, ZN => n13615);
   U5629 : OAI22_X1 port map( A1 => n60761, A2 => n60959, B1 => n1717, B2 => 
                           n60758, ZN => n13616);
   U5630 : OAI22_X1 port map( A1 => n60761, A2 => n60973, B1 => n1716, B2 => 
                           n15135, ZN => n13617);
   U5631 : OAI22_X1 port map( A1 => n60761, A2 => n60987, B1 => n1715, B2 => 
                           n15135, ZN => n13618);
   U5632 : OAI22_X1 port map( A1 => n60761, A2 => n61001, B1 => n1714, B2 => 
                           n15135, ZN => n13619);
   U5633 : OAI22_X1 port map( A1 => n60762, A2 => n61015, B1 => n1713, B2 => 
                           n15135, ZN => n13620);
   U5634 : OAI22_X1 port map( A1 => n60762, A2 => n61029, B1 => n1712, B2 => 
                           n15135, ZN => n13621);
   U5635 : OAI22_X1 port map( A1 => n60762, A2 => n61043, B1 => n1711, B2 => 
                           n15135, ZN => n13622);
   U5636 : OAI22_X1 port map( A1 => n60762, A2 => n61057, B1 => n1710, B2 => 
                           n15135, ZN => n13623);
   U5637 : OAI22_X1 port map( A1 => n60762, A2 => n61071, B1 => n1709, B2 => 
                           n60758, ZN => n13624);
   U5638 : OAI22_X1 port map( A1 => n60763, A2 => n61085, B1 => n1708, B2 => 
                           n60758, ZN => n13625);
   U5639 : OAI22_X1 port map( A1 => n60763, A2 => n61099, B1 => n1707, B2 => 
                           n60758, ZN => n13626);
   U5640 : OAI22_X1 port map( A1 => n60763, A2 => n61113, B1 => n1706, B2 => 
                           n60758, ZN => n13627);
   U5641 : OAI22_X1 port map( A1 => n60763, A2 => n61127, B1 => n1705, B2 => 
                           n60758, ZN => n13628);
   U5642 : OAI22_X1 port map( A1 => n60732, A2 => n61967, B1 => n1616, B2 => 
                           n60731, ZN => n13509);
   U5643 : OAI22_X1 port map( A1 => n60732, A2 => n61981, B1 => n1615, B2 => 
                           n60731, ZN => n13510);
   U5644 : OAI22_X1 port map( A1 => n60732, A2 => n61995, B1 => n1614, B2 => 
                           n60731, ZN => n13511);
   U5645 : OAI22_X1 port map( A1 => n60732, A2 => n62009, B1 => n1613, B2 => 
                           n60731, ZN => n13512);
   U5646 : OAI22_X1 port map( A1 => n60732, A2 => n62023, B1 => n1612, B2 => 
                           n60731, ZN => n13513);
   U5647 : OAI22_X1 port map( A1 => n60733, A2 => n62037, B1 => n1611, B2 => 
                           n60731, ZN => n13514);
   U5648 : OAI22_X1 port map( A1 => n60733, A2 => n62051, B1 => n1610, B2 => 
                           n60731, ZN => n13515);
   U5649 : OAI22_X1 port map( A1 => n60733, A2 => n62065, B1 => n1609, B2 => 
                           n60731, ZN => n13516);
   U5650 : OAI22_X1 port map( A1 => n60733, A2 => n62079, B1 => n1608, B2 => 
                           n60731, ZN => n13517);
   U5651 : OAI22_X1 port map( A1 => n60733, A2 => n62093, B1 => n1607, B2 => 
                           n60731, ZN => n13518);
   U5652 : OAI22_X1 port map( A1 => n60734, A2 => n62107, B1 => n1590, B2 => 
                           n60731, ZN => n13519);
   U5653 : OAI22_X1 port map( A1 => n60734, A2 => n60960, B1 => n1589, B2 => 
                           n60731, ZN => n13520);
   U5654 : OAI22_X1 port map( A1 => n60734, A2 => n60974, B1 => n1558, B2 => 
                           n15138, ZN => n13521);
   U5655 : OAI22_X1 port map( A1 => n60734, A2 => n60988, B1 => n1557, B2 => 
                           n15138, ZN => n13522);
   U5656 : OAI22_X1 port map( A1 => n60734, A2 => n61002, B1 => n1556, B2 => 
                           n15138, ZN => n13523);
   U5657 : OAI22_X1 port map( A1 => n60735, A2 => n61016, B1 => n1555, B2 => 
                           n15138, ZN => n13524);
   U5658 : OAI22_X1 port map( A1 => n60735, A2 => n61030, B1 => n1554, B2 => 
                           n15138, ZN => n13525);
   U5659 : OAI22_X1 port map( A1 => n60735, A2 => n61044, B1 => n1553, B2 => 
                           n15138, ZN => n13526);
   U5660 : OAI22_X1 port map( A1 => n60735, A2 => n61058, B1 => n1552, B2 => 
                           n15138, ZN => n13527);
   U5661 : OAI22_X1 port map( A1 => n60735, A2 => n61072, B1 => n1551, B2 => 
                           n60731, ZN => n13528);
   U5662 : OAI22_X1 port map( A1 => n60736, A2 => n61086, B1 => n1550, B2 => 
                           n60731, ZN => n13529);
   U5663 : OAI22_X1 port map( A1 => n60736, A2 => n61100, B1 => n1549, B2 => 
                           n60731, ZN => n13530);
   U5664 : OAI22_X1 port map( A1 => n60736, A2 => n61114, B1 => n1548, B2 => 
                           n60731, ZN => n13531);
   U5665 : OAI22_X1 port map( A1 => n60736, A2 => n61128, B1 => n1547, B2 => 
                           n60731, ZN => n13532);
   U5666 : OAI22_X1 port map( A1 => n60723, A2 => n61967, B1 => n1546, B2 => 
                           n60722, ZN => n13477);
   U5667 : OAI22_X1 port map( A1 => n60723, A2 => n61981, B1 => n1544, B2 => 
                           n60722, ZN => n13478);
   U5668 : OAI22_X1 port map( A1 => n60723, A2 => n61995, B1 => n1542, B2 => 
                           n60722, ZN => n13479);
   U5669 : OAI22_X1 port map( A1 => n60723, A2 => n62009, B1 => n1540, B2 => 
                           n60722, ZN => n13480);
   U5670 : OAI22_X1 port map( A1 => n60723, A2 => n62023, B1 => n1538, B2 => 
                           n60722, ZN => n13481);
   U5671 : OAI22_X1 port map( A1 => n60724, A2 => n62037, B1 => n1536, B2 => 
                           n60722, ZN => n13482);
   U5672 : OAI22_X1 port map( A1 => n60724, A2 => n62051, B1 => n1534, B2 => 
                           n60722, ZN => n13483);
   U5673 : OAI22_X1 port map( A1 => n60724, A2 => n62065, B1 => n1532, B2 => 
                           n60722, ZN => n13484);
   U5674 : OAI22_X1 port map( A1 => n60724, A2 => n62079, B1 => n1530, B2 => 
                           n60722, ZN => n13485);
   U5675 : OAI22_X1 port map( A1 => n60724, A2 => n62093, B1 => n1528, B2 => 
                           n60722, ZN => n13486);
   U5676 : OAI22_X1 port map( A1 => n60725, A2 => n62107, B1 => n1526, B2 => 
                           n60722, ZN => n13487);
   U5677 : OAI22_X1 port map( A1 => n60725, A2 => n60960, B1 => n1524, B2 => 
                           n60722, ZN => n13488);
   U5678 : OAI22_X1 port map( A1 => n60725, A2 => n60974, B1 => n1522, B2 => 
                           n15139, ZN => n13489);
   U5679 : OAI22_X1 port map( A1 => n60725, A2 => n60988, B1 => n1520, B2 => 
                           n15139, ZN => n13490);
   U5680 : OAI22_X1 port map( A1 => n60725, A2 => n61002, B1 => n1517, B2 => 
                           n15139, ZN => n13491);
   U5681 : OAI22_X1 port map( A1 => n60726, A2 => n61016, B1 => n1516, B2 => 
                           n15139, ZN => n13492);
   U5682 : OAI22_X1 port map( A1 => n60726, A2 => n61030, B1 => n1515, B2 => 
                           n15139, ZN => n13493);
   U5683 : OAI22_X1 port map( A1 => n60726, A2 => n61044, B1 => n1514, B2 => 
                           n15139, ZN => n13494);
   U5684 : OAI22_X1 port map( A1 => n60726, A2 => n61058, B1 => n1513, B2 => 
                           n15139, ZN => n13495);
   U5685 : OAI22_X1 port map( A1 => n60726, A2 => n61072, B1 => n1512, B2 => 
                           n60722, ZN => n13496);
   U5686 : OAI22_X1 port map( A1 => n60727, A2 => n61086, B1 => n1511, B2 => 
                           n60722, ZN => n13497);
   U5687 : OAI22_X1 port map( A1 => n60727, A2 => n61100, B1 => n1510, B2 => 
                           n60722, ZN => n13498);
   U5688 : OAI22_X1 port map( A1 => n60727, A2 => n61114, B1 => n1509, B2 => 
                           n60722, ZN => n13499);
   U5689 : OAI22_X1 port map( A1 => n60727, A2 => n61128, B1 => n1508, B2 => 
                           n60722, ZN => n13500);
   U5690 : OAI22_X1 port map( A1 => n60696, A2 => n61967, B1 => n1506, B2 => 
                           n60695, ZN => n13381);
   U5691 : OAI22_X1 port map( A1 => n60696, A2 => n61981, B1 => n1505, B2 => 
                           n60695, ZN => n13382);
   U5692 : OAI22_X1 port map( A1 => n60696, A2 => n61995, B1 => n1504, B2 => 
                           n60695, ZN => n13383);
   U5693 : OAI22_X1 port map( A1 => n60696, A2 => n62009, B1 => n1503, B2 => 
                           n60695, ZN => n13384);
   U5694 : OAI22_X1 port map( A1 => n60696, A2 => n62023, B1 => n1502, B2 => 
                           n60695, ZN => n13385);
   U5695 : OAI22_X1 port map( A1 => n60697, A2 => n62037, B1 => n1501, B2 => 
                           n60695, ZN => n13386);
   U5696 : OAI22_X1 port map( A1 => n60697, A2 => n62051, B1 => n1500, B2 => 
                           n60695, ZN => n13387);
   U5697 : OAI22_X1 port map( A1 => n60697, A2 => n62065, B1 => n1499, B2 => 
                           n60695, ZN => n13388);
   U5698 : OAI22_X1 port map( A1 => n60697, A2 => n62079, B1 => n1498, B2 => 
                           n60695, ZN => n13389);
   U5699 : OAI22_X1 port map( A1 => n60697, A2 => n62093, B1 => n1497, B2 => 
                           n60695, ZN => n13390);
   U5700 : OAI22_X1 port map( A1 => n60698, A2 => n62107, B1 => n1496, B2 => 
                           n60695, ZN => n13391);
   U5701 : OAI22_X1 port map( A1 => n60698, A2 => n60960, B1 => n1495, B2 => 
                           n60695, ZN => n13392);
   U5702 : OAI22_X1 port map( A1 => n60698, A2 => n60974, B1 => n1494, B2 => 
                           n15142, ZN => n13393);
   U5703 : OAI22_X1 port map( A1 => n60698, A2 => n60988, B1 => n1493, B2 => 
                           n15142, ZN => n13394);
   U5704 : OAI22_X1 port map( A1 => n60698, A2 => n61002, B1 => n1492, B2 => 
                           n15142, ZN => n13395);
   U5705 : OAI22_X1 port map( A1 => n60699, A2 => n61016, B1 => n1491, B2 => 
                           n15142, ZN => n13396);
   U5706 : OAI22_X1 port map( A1 => n60699, A2 => n61030, B1 => n1490, B2 => 
                           n15142, ZN => n13397);
   U5707 : OAI22_X1 port map( A1 => n60699, A2 => n61044, B1 => n1489, B2 => 
                           n15142, ZN => n13398);
   U5708 : OAI22_X1 port map( A1 => n60699, A2 => n61058, B1 => n1488, B2 => 
                           n15142, ZN => n13399);
   U5709 : OAI22_X1 port map( A1 => n60699, A2 => n61072, B1 => n1487, B2 => 
                           n60695, ZN => n13400);
   U5710 : OAI22_X1 port map( A1 => n60700, A2 => n61086, B1 => n1486, B2 => 
                           n60695, ZN => n13401);
   U5711 : OAI22_X1 port map( A1 => n60700, A2 => n61100, B1 => n1485, B2 => 
                           n60695, ZN => n13402);
   U5712 : OAI22_X1 port map( A1 => n60700, A2 => n61114, B1 => n1484, B2 => 
                           n60695, ZN => n13403);
   U5713 : OAI22_X1 port map( A1 => n60700, A2 => n61128, B1 => n1483, B2 => 
                           n60695, ZN => n13404);
   U5714 : OAI22_X1 port map( A1 => n60687, A2 => n61967, B1 => n1482, B2 => 
                           n60686, ZN => n13349);
   U5715 : OAI22_X1 port map( A1 => n60687, A2 => n61981, B1 => n1481, B2 => 
                           n60686, ZN => n13350);
   U5716 : OAI22_X1 port map( A1 => n60687, A2 => n61995, B1 => n1480, B2 => 
                           n60686, ZN => n13351);
   U5717 : OAI22_X1 port map( A1 => n60687, A2 => n62009, B1 => n1479, B2 => 
                           n60686, ZN => n13352);
   U5718 : OAI22_X1 port map( A1 => n60687, A2 => n62023, B1 => n1478, B2 => 
                           n60686, ZN => n13353);
   U5719 : OAI22_X1 port map( A1 => n60688, A2 => n62037, B1 => n1477, B2 => 
                           n60686, ZN => n13354);
   U5720 : OAI22_X1 port map( A1 => n60688, A2 => n62051, B1 => n1476, B2 => 
                           n60686, ZN => n13355);
   U5721 : OAI22_X1 port map( A1 => n60688, A2 => n62065, B1 => n1475, B2 => 
                           n60686, ZN => n13356);
   U5722 : OAI22_X1 port map( A1 => n60688, A2 => n62079, B1 => n1474, B2 => 
                           n60686, ZN => n13357);
   U5723 : OAI22_X1 port map( A1 => n60688, A2 => n62093, B1 => n1473, B2 => 
                           n60686, ZN => n13358);
   U5724 : OAI22_X1 port map( A1 => n60689, A2 => n62107, B1 => n1472, B2 => 
                           n60686, ZN => n13359);
   U5725 : OAI22_X1 port map( A1 => n60689, A2 => n60960, B1 => n1471, B2 => 
                           n60686, ZN => n13360);
   U5726 : OAI22_X1 port map( A1 => n60689, A2 => n60974, B1 => n1470, B2 => 
                           n15143, ZN => n13361);
   U5727 : OAI22_X1 port map( A1 => n60689, A2 => n60988, B1 => n1469, B2 => 
                           n15143, ZN => n13362);
   U5728 : OAI22_X1 port map( A1 => n60689, A2 => n61002, B1 => n1468, B2 => 
                           n15143, ZN => n13363);
   U5729 : OAI22_X1 port map( A1 => n60690, A2 => n61016, B1 => n1467, B2 => 
                           n15143, ZN => n13364);
   U5730 : OAI22_X1 port map( A1 => n60690, A2 => n61030, B1 => n1466, B2 => 
                           n15143, ZN => n13365);
   U5731 : OAI22_X1 port map( A1 => n60690, A2 => n61044, B1 => n1465, B2 => 
                           n15143, ZN => n13366);
   U5732 : OAI22_X1 port map( A1 => n60690, A2 => n61058, B1 => n1464, B2 => 
                           n15143, ZN => n13367);
   U5733 : OAI22_X1 port map( A1 => n60690, A2 => n61072, B1 => n1463, B2 => 
                           n60686, ZN => n13368);
   U5734 : OAI22_X1 port map( A1 => n60691, A2 => n61086, B1 => n1462, B2 => 
                           n60686, ZN => n13369);
   U5735 : OAI22_X1 port map( A1 => n60691, A2 => n61100, B1 => n1461, B2 => 
                           n60686, ZN => n13370);
   U5736 : OAI22_X1 port map( A1 => n60691, A2 => n61114, B1 => n1460, B2 => 
                           n60686, ZN => n13371);
   U5737 : OAI22_X1 port map( A1 => n60691, A2 => n61128, B1 => n1459, B2 => 
                           n60686, ZN => n13372);
   U5738 : OAI22_X1 port map( A1 => n59796, A2 => n61975, B1 => n1410, B2 => 
                           n59795, ZN => n10181);
   U5739 : OAI22_X1 port map( A1 => n59796, A2 => n61989, B1 => n1409, B2 => 
                           n59795, ZN => n10182);
   U5740 : OAI22_X1 port map( A1 => n59796, A2 => n62003, B1 => n1408, B2 => 
                           n59795, ZN => n10183);
   U5741 : OAI22_X1 port map( A1 => n59796, A2 => n62017, B1 => n1407, B2 => 
                           n59795, ZN => n10184);
   U5742 : OAI22_X1 port map( A1 => n59796, A2 => n62031, B1 => n1406, B2 => 
                           n59795, ZN => n10185);
   U5743 : OAI22_X1 port map( A1 => n59797, A2 => n62045, B1 => n1405, B2 => 
                           n59795, ZN => n10186);
   U5744 : OAI22_X1 port map( A1 => n59797, A2 => n62059, B1 => n1404, B2 => 
                           n59795, ZN => n10187);
   U5745 : OAI22_X1 port map( A1 => n59797, A2 => n62073, B1 => n1403, B2 => 
                           n59795, ZN => n10188);
   U5746 : OAI22_X1 port map( A1 => n59797, A2 => n62087, B1 => n1402, B2 => 
                           n59795, ZN => n10189);
   U5747 : OAI22_X1 port map( A1 => n59797, A2 => n62101, B1 => n1401, B2 => 
                           n59795, ZN => n10190);
   U5748 : OAI22_X1 port map( A1 => n59798, A2 => n62115, B1 => n1400, B2 => 
                           n59795, ZN => n10191);
   U5749 : OAI22_X1 port map( A1 => n59798, A2 => n60968, B1 => n1399, B2 => 
                           n59795, ZN => n10192);
   U5750 : OAI22_X1 port map( A1 => n59798, A2 => n60982, B1 => n1398, B2 => 
                           n15280, ZN => n10193);
   U5751 : OAI22_X1 port map( A1 => n59798, A2 => n60996, B1 => n1397, B2 => 
                           n15280, ZN => n10194);
   U5752 : OAI22_X1 port map( A1 => n59798, A2 => n61010, B1 => n1396, B2 => 
                           n15280, ZN => n10195);
   U5753 : OAI22_X1 port map( A1 => n59799, A2 => n61024, B1 => n1395, B2 => 
                           n15280, ZN => n10196);
   U5754 : OAI22_X1 port map( A1 => n59799, A2 => n61038, B1 => n1394, B2 => 
                           n15280, ZN => n10197);
   U5755 : OAI22_X1 port map( A1 => n59799, A2 => n61052, B1 => n1393, B2 => 
                           n15280, ZN => n10198);
   U5756 : OAI22_X1 port map( A1 => n59799, A2 => n61066, B1 => n1392, B2 => 
                           n15280, ZN => n10199);
   U5757 : OAI22_X1 port map( A1 => n59799, A2 => n61080, B1 => n1391, B2 => 
                           n59795, ZN => n10200);
   U5758 : OAI22_X1 port map( A1 => n59800, A2 => n61094, B1 => n1390, B2 => 
                           n59795, ZN => n10201);
   U5759 : OAI22_X1 port map( A1 => n59800, A2 => n61108, B1 => n1389, B2 => 
                           n59795, ZN => n10202);
   U5760 : OAI22_X1 port map( A1 => n59800, A2 => n61122, B1 => n1388, B2 => 
                           n59795, ZN => n10203);
   U5761 : OAI22_X1 port map( A1 => n59800, A2 => n61136, B1 => n1387, B2 => 
                           n59795, ZN => n10204);
   U5762 : OAI22_X1 port map( A1 => n59787, A2 => n61975, B1 => n1386, B2 => 
                           n59786, ZN => n10149);
   U5763 : OAI22_X1 port map( A1 => n59787, A2 => n61989, B1 => n1385, B2 => 
                           n59786, ZN => n10150);
   U5764 : OAI22_X1 port map( A1 => n59787, A2 => n62003, B1 => n1384, B2 => 
                           n59786, ZN => n10151);
   U5765 : OAI22_X1 port map( A1 => n59787, A2 => n62017, B1 => n1383, B2 => 
                           n59786, ZN => n10152);
   U5766 : OAI22_X1 port map( A1 => n59787, A2 => n62031, B1 => n1382, B2 => 
                           n59786, ZN => n10153);
   U5767 : OAI22_X1 port map( A1 => n59788, A2 => n62045, B1 => n1381, B2 => 
                           n59786, ZN => n10154);
   U5768 : OAI22_X1 port map( A1 => n59788, A2 => n62059, B1 => n1380, B2 => 
                           n59786, ZN => n10155);
   U5769 : OAI22_X1 port map( A1 => n59788, A2 => n62073, B1 => n1379, B2 => 
                           n59786, ZN => n10156);
   U5770 : OAI22_X1 port map( A1 => n59788, A2 => n62087, B1 => n1378, B2 => 
                           n59786, ZN => n10157);
   U5771 : OAI22_X1 port map( A1 => n59788, A2 => n62101, B1 => n1377, B2 => 
                           n59786, ZN => n10158);
   U5772 : OAI22_X1 port map( A1 => n59789, A2 => n62115, B1 => n1376, B2 => 
                           n59786, ZN => n10159);
   U5773 : OAI22_X1 port map( A1 => n59789, A2 => n60968, B1 => n1375, B2 => 
                           n59786, ZN => n10160);
   U5774 : OAI22_X1 port map( A1 => n59789, A2 => n60982, B1 => n1374, B2 => 
                           n15281, ZN => n10161);
   U5775 : OAI22_X1 port map( A1 => n59789, A2 => n60996, B1 => n1373, B2 => 
                           n15281, ZN => n10162);
   U5776 : OAI22_X1 port map( A1 => n59789, A2 => n61010, B1 => n1372, B2 => 
                           n15281, ZN => n10163);
   U5777 : OAI22_X1 port map( A1 => n59790, A2 => n61024, B1 => n1371, B2 => 
                           n15281, ZN => n10164);
   U5778 : OAI22_X1 port map( A1 => n59790, A2 => n61038, B1 => n1370, B2 => 
                           n15281, ZN => n10165);
   U5779 : OAI22_X1 port map( A1 => n59790, A2 => n61052, B1 => n1369, B2 => 
                           n15281, ZN => n10166);
   U5780 : OAI22_X1 port map( A1 => n59790, A2 => n61066, B1 => n1368, B2 => 
                           n15281, ZN => n10167);
   U5781 : OAI22_X1 port map( A1 => n59790, A2 => n61080, B1 => n1367, B2 => 
                           n59786, ZN => n10168);
   U5782 : OAI22_X1 port map( A1 => n59791, A2 => n61094, B1 => n1366, B2 => 
                           n59786, ZN => n10169);
   U5783 : OAI22_X1 port map( A1 => n59791, A2 => n61108, B1 => n1365, B2 => 
                           n59786, ZN => n10170);
   U5784 : OAI22_X1 port map( A1 => n59791, A2 => n61122, B1 => n1364, B2 => 
                           n59786, ZN => n10171);
   U5785 : OAI22_X1 port map( A1 => n59791, A2 => n61136, B1 => n1363, B2 => 
                           n59786, ZN => n10172);
   U5786 : OAI22_X1 port map( A1 => n59780, A2 => n60968, B1 => n1362, B2 => 
                           n15282, ZN => n10128);
   U5787 : OAI22_X1 port map( A1 => n59780, A2 => n60982, B1 => n1361, B2 => 
                           n59777, ZN => n10129);
   U5788 : OAI22_X1 port map( A1 => n59780, A2 => n60996, B1 => n1360, B2 => 
                           n59777, ZN => n10130);
   U5789 : OAI22_X1 port map( A1 => n59780, A2 => n61010, B1 => n1359, B2 => 
                           n59777, ZN => n10131);
   U5790 : OAI22_X1 port map( A1 => n59781, A2 => n61024, B1 => n1358, B2 => 
                           n59777, ZN => n10132);
   U5791 : OAI22_X1 port map( A1 => n59781, A2 => n61038, B1 => n1357, B2 => 
                           n59777, ZN => n10133);
   U5792 : OAI22_X1 port map( A1 => n59781, A2 => n61052, B1 => n1356, B2 => 
                           n59777, ZN => n10134);
   U5793 : OAI22_X1 port map( A1 => n59781, A2 => n61066, B1 => n1355, B2 => 
                           n59777, ZN => n10135);
   U5794 : OAI22_X1 port map( A1 => n59781, A2 => n61080, B1 => n1354, B2 => 
                           n59777, ZN => n10136);
   U5795 : OAI22_X1 port map( A1 => n59782, A2 => n61094, B1 => n1353, B2 => 
                           n59777, ZN => n10137);
   U5796 : OAI22_X1 port map( A1 => n59782, A2 => n61108, B1 => n1352, B2 => 
                           n59777, ZN => n10138);
   U5797 : OAI22_X1 port map( A1 => n59782, A2 => n61122, B1 => n1351, B2 => 
                           n59777, ZN => n10139);
   U5798 : OAI22_X1 port map( A1 => n59782, A2 => n61136, B1 => n1350, B2 => 
                           n59777, ZN => n10140);
   U5799 : OAI22_X1 port map( A1 => n59769, A2 => n61975, B1 => n1349, B2 => 
                           n59768, ZN => n10085);
   U5800 : OAI22_X1 port map( A1 => n59769, A2 => n61989, B1 => n1348, B2 => 
                           n59768, ZN => n10086);
   U5801 : OAI22_X1 port map( A1 => n59769, A2 => n62003, B1 => n1347, B2 => 
                           n59768, ZN => n10087);
   U5802 : OAI22_X1 port map( A1 => n59769, A2 => n62017, B1 => n1346, B2 => 
                           n59768, ZN => n10088);
   U5803 : OAI22_X1 port map( A1 => n59769, A2 => n62031, B1 => n1345, B2 => 
                           n59768, ZN => n10089);
   U5804 : OAI22_X1 port map( A1 => n59770, A2 => n62045, B1 => n1344, B2 => 
                           n59768, ZN => n10090);
   U5805 : OAI22_X1 port map( A1 => n59770, A2 => n62059, B1 => n1343, B2 => 
                           n59768, ZN => n10091);
   U5806 : OAI22_X1 port map( A1 => n59770, A2 => n62073, B1 => n1342, B2 => 
                           n59768, ZN => n10092);
   U5807 : OAI22_X1 port map( A1 => n59770, A2 => n62087, B1 => n1341, B2 => 
                           n59768, ZN => n10093);
   U5808 : OAI22_X1 port map( A1 => n59770, A2 => n62101, B1 => n1340, B2 => 
                           n59768, ZN => n10094);
   U5809 : OAI22_X1 port map( A1 => n59771, A2 => n62115, B1 => n1339, B2 => 
                           n59768, ZN => n10095);
   U5810 : OAI22_X1 port map( A1 => n59778, A2 => n61976, B1 => n1338, B2 => 
                           n15282, ZN => n10117);
   U5811 : OAI22_X1 port map( A1 => n59778, A2 => n61990, B1 => n1337, B2 => 
                           n15282, ZN => n10118);
   U5812 : OAI22_X1 port map( A1 => n59778, A2 => n62004, B1 => n1336, B2 => 
                           n15282, ZN => n10119);
   U5813 : OAI22_X1 port map( A1 => n59778, A2 => n62018, B1 => n1335, B2 => 
                           n15282, ZN => n10120);
   U5814 : OAI22_X1 port map( A1 => n59778, A2 => n62032, B1 => n1334, B2 => 
                           n15282, ZN => n10121);
   U5815 : OAI22_X1 port map( A1 => n59779, A2 => n62046, B1 => n1333, B2 => 
                           n15282, ZN => n10122);
   U5816 : OAI22_X1 port map( A1 => n59779, A2 => n62060, B1 => n1332, B2 => 
                           n59777, ZN => n10123);
   U5817 : OAI22_X1 port map( A1 => n59779, A2 => n62074, B1 => n1331, B2 => 
                           n59777, ZN => n10124);
   U5818 : OAI22_X1 port map( A1 => n59779, A2 => n62088, B1 => n1330, B2 => 
                           n59777, ZN => n10125);
   U5819 : OAI22_X1 port map( A1 => n59779, A2 => n62102, B1 => n1329, B2 => 
                           n59777, ZN => n10126);
   U5820 : OAI22_X1 port map( A1 => n59780, A2 => n62116, B1 => n1328, B2 => 
                           n59777, ZN => n10127);
   U5821 : OAI22_X1 port map( A1 => n59771, A2 => n60969, B1 => n1327, B2 => 
                           n59768, ZN => n10096);
   U5822 : OAI22_X1 port map( A1 => n59771, A2 => n60983, B1 => n1326, B2 => 
                           n15283, ZN => n10097);
   U5823 : OAI22_X1 port map( A1 => n59771, A2 => n60997, B1 => n1325, B2 => 
                           n15283, ZN => n10098);
   U5824 : OAI22_X1 port map( A1 => n59771, A2 => n61011, B1 => n1324, B2 => 
                           n15283, ZN => n10099);
   U5825 : OAI22_X1 port map( A1 => n59772, A2 => n61025, B1 => n1323, B2 => 
                           n15283, ZN => n10100);
   U5826 : OAI22_X1 port map( A1 => n59772, A2 => n61039, B1 => n1322, B2 => 
                           n15283, ZN => n10101);
   U5827 : OAI22_X1 port map( A1 => n59772, A2 => n61053, B1 => n1321, B2 => 
                           n15283, ZN => n10102);
   U5828 : OAI22_X1 port map( A1 => n59772, A2 => n61067, B1 => n1320, B2 => 
                           n15283, ZN => n10103);
   U5829 : OAI22_X1 port map( A1 => n59772, A2 => n61081, B1 => n1319, B2 => 
                           n59768, ZN => n10104);
   U5830 : OAI22_X1 port map( A1 => n59773, A2 => n61095, B1 => n1318, B2 => 
                           n59768, ZN => n10105);
   U5831 : OAI22_X1 port map( A1 => n59773, A2 => n61109, B1 => n1317, B2 => 
                           n59768, ZN => n10106);
   U5832 : OAI22_X1 port map( A1 => n59773, A2 => n61123, B1 => n1316, B2 => 
                           n59768, ZN => n10107);
   U5833 : OAI22_X1 port map( A1 => n59773, A2 => n61137, B1 => n1315, B2 => 
                           n59768, ZN => n10108);
   U5834 : AND2_X1 port map( A1 => ADDR_WR(3), A2 => ADDR_WR(2), ZN => n15265);
   U5835 : OAI21_X1 port map( B1 => n15270, B2 => n15107, A => n62197, ZN => 
                           n15286);
   U5836 : INV_X1 port map( A => ADDR_WR(0), ZN => n5283);
   U5837 : INV_X1 port map( A => ADDR_WR(1), ZN => n5282);
   U5838 : INV_X1 port map( A => n15269, ZN => n59812);
   U5839 : OAI21_X1 port map( B1 => n15270, B2 => n15095, A => n62197, ZN => 
                           n15269);
   U5840 : INV_X1 port map( A => n15280, ZN => n59803);
   U5841 : OAI21_X1 port map( B1 => n15270, B2 => n15097, A => n62197, ZN => 
                           n15280);
   U5842 : INV_X1 port map( A => n15281, ZN => n59794);
   U5843 : OAI21_X1 port map( B1 => n15270, B2 => n15099, A => n62197, ZN => 
                           n15281);
   U5844 : INV_X1 port map( A => n15282, ZN => n59785);
   U5845 : OAI21_X1 port map( B1 => n15270, B2 => n15101, A => n62197, ZN => 
                           n15282);
   U5846 : INV_X1 port map( A => n15283, ZN => n59776);
   U5847 : OAI21_X1 port map( B1 => n15270, B2 => n15103, A => n62198, ZN => 
                           n15283);
   U5848 : INV_X1 port map( A => n15285, ZN => n59767);
   U5849 : OAI21_X1 port map( B1 => n15270, B2 => n15105, A => n62198, ZN => 
                           n15285);
   U5850 : INV_X1 port map( A => ADDR_WR(2), ZN => n5281);
   U5851 : BUF_X1 port map( A => n5374, Z => n61959);
   U5852 : BUF_X1 port map( A => n5374, Z => n61961);
   U5853 : BUF_X1 port map( A => n5374, Z => n61960);
   U5854 : BUF_X1 port map( A => n5374, Z => n61957);
   U5855 : BUF_X1 port map( A => n5374, Z => n61958);
   U5856 : BUF_X1 port map( A => n5373, Z => n61963);
   U5857 : BUF_X1 port map( A => n5372, Z => n61977);
   U5858 : BUF_X1 port map( A => n5371, Z => n61991);
   U5859 : BUF_X1 port map( A => n5370, Z => n62005);
   U5860 : BUF_X1 port map( A => n5369, Z => n62019);
   U5861 : BUF_X1 port map( A => n5368, Z => n62033);
   U5862 : BUF_X1 port map( A => n5367, Z => n62047);
   U5863 : BUF_X1 port map( A => n5366, Z => n62061);
   U5864 : BUF_X1 port map( A => n5365, Z => n62075);
   U5865 : BUF_X1 port map( A => n5364, Z => n62089);
   U5866 : BUF_X1 port map( A => n5363, Z => n62103);
   U5867 : BUF_X1 port map( A => n15093, Z => n60956);
   U5868 : BUF_X1 port map( A => n15092, Z => n60970);
   U5869 : BUF_X1 port map( A => n15091, Z => n60984);
   U5870 : BUF_X1 port map( A => n15090, Z => n60998);
   U5871 : BUF_X1 port map( A => n15089, Z => n61012);
   U5872 : BUF_X1 port map( A => n15088, Z => n61026);
   U5873 : BUF_X1 port map( A => n15087, Z => n61040);
   U5874 : BUF_X1 port map( A => n15086, Z => n61054);
   U5875 : BUF_X1 port map( A => n15085, Z => n61068);
   U5876 : BUF_X1 port map( A => n15084, Z => n61082);
   U5877 : BUF_X1 port map( A => n15083, Z => n61096);
   U5878 : BUF_X1 port map( A => n15082, Z => n61110);
   U5879 : BUF_X1 port map( A => n15081, Z => n61124);
   U5880 : BUF_X1 port map( A => n15080, Z => n61138);
   U5881 : BUF_X1 port map( A => n15079, Z => n61152);
   U5882 : BUF_X1 port map( A => n15078, Z => n61166);
   U5883 : BUF_X1 port map( A => n15077, Z => n61180);
   U5884 : BUF_X1 port map( A => n15076, Z => n61194);
   U5885 : BUF_X1 port map( A => n15075, Z => n61208);
   U5886 : BUF_X1 port map( A => n15074, Z => n61222);
   U5887 : BUF_X1 port map( A => n15072, Z => n61245);
   U5888 : BUF_X1 port map( A => n5373, Z => n61964);
   U5889 : BUF_X1 port map( A => n5372, Z => n61978);
   U5890 : BUF_X1 port map( A => n5371, Z => n61992);
   U5891 : BUF_X1 port map( A => n5370, Z => n62006);
   U5892 : BUF_X1 port map( A => n5369, Z => n62020);
   U5893 : BUF_X1 port map( A => n5368, Z => n62034);
   U5894 : BUF_X1 port map( A => n5367, Z => n62048);
   U5895 : BUF_X1 port map( A => n5366, Z => n62062);
   U5896 : BUF_X1 port map( A => n5365, Z => n62076);
   U5897 : BUF_X1 port map( A => n5364, Z => n62090);
   U5898 : BUF_X1 port map( A => n5363, Z => n62104);
   U5899 : BUF_X1 port map( A => n15085, Z => n61069);
   U5900 : BUF_X1 port map( A => n15084, Z => n61083);
   U5901 : BUF_X1 port map( A => n15083, Z => n61097);
   U5902 : BUF_X1 port map( A => n15082, Z => n61111);
   U5903 : BUF_X1 port map( A => n15081, Z => n61125);
   U5904 : BUF_X1 port map( A => n15093, Z => n60957);
   U5905 : BUF_X1 port map( A => n15092, Z => n60971);
   U5906 : BUF_X1 port map( A => n15091, Z => n60985);
   U5907 : BUF_X1 port map( A => n15090, Z => n60999);
   U5908 : BUF_X1 port map( A => n15089, Z => n61013);
   U5909 : BUF_X1 port map( A => n15088, Z => n61027);
   U5910 : BUF_X1 port map( A => n15087, Z => n61041);
   U5911 : BUF_X1 port map( A => n15086, Z => n61055);
   U5912 : BUF_X1 port map( A => n15080, Z => n61139);
   U5913 : BUF_X1 port map( A => n15079, Z => n61153);
   U5914 : BUF_X1 port map( A => n15078, Z => n61167);
   U5915 : BUF_X1 port map( A => n15077, Z => n61181);
   U5916 : BUF_X1 port map( A => n15076, Z => n61195);
   U5917 : BUF_X1 port map( A => n15075, Z => n61209);
   U5918 : BUF_X1 port map( A => n15074, Z => n61223);
   U5919 : BUF_X1 port map( A => n15072, Z => n61246);
   U5920 : BUF_X1 port map( A => n7943, Z => n61669);
   U5921 : BUF_X1 port map( A => n7943, Z => n61671);
   U5922 : BUF_X1 port map( A => n7943, Z => n61670);
   U5923 : BUF_X1 port map( A => n7943, Z => n61667);
   U5924 : BUF_X1 port map( A => n7943, Z => n61668);
   U5925 : BUF_X1 port map( A => n5276, Z => n62183);
   U5926 : BUF_X1 port map( A => n5276, Z => n62182);
   U5927 : BUF_X1 port map( A => n5276, Z => n62184);
   U5928 : NAND4_X1 port map( A1 => n15127, A2 => n5280, A3 => ADDR_WR(7), A4 
                           => n15287, ZN => n15270);
   U5929 : AND2_X1 port map( A1 => EN, A2 => WR, ZN => n15287);
   U5930 : AOI222_X1 port map( A1 => n16232, A2 => n5288, B1 => n15602, B2 => 
                           n5293, C1 => n16231, C2 => n5289, ZN => n6733);
   U5931 : AOI222_X1 port map( A1 => n16238, A2 => n5288, B1 => n15603, B2 => 
                           n5293, C1 => n16237, C2 => n5289, ZN => n6658);
   U5932 : AOI222_X1 port map( A1 => n16244, A2 => n5288, B1 => n15604, B2 => 
                           n5293, C1 => n16243, C2 => n5289, ZN => n6583);
   U5933 : AOI222_X1 port map( A1 => n16250, A2 => n5288, B1 => n15605, B2 => 
                           n5293, C1 => n16249, C2 => n5289, ZN => n6508);
   U5934 : AOI222_X1 port map( A1 => n16256, A2 => n5288, B1 => n15606, B2 => 
                           n5293, C1 => n16255, C2 => n5289, ZN => n6433);
   U5935 : AOI222_X1 port map( A1 => n16190, A2 => n5288, B1 => n15607, B2 => 
                           n5293, C1 => n16189, C2 => n5289, ZN => n6358);
   U5936 : AOI222_X1 port map( A1 => n16196, A2 => n5288, B1 => n15608, B2 => 
                           n5293, C1 => n16195, C2 => n5289, ZN => n6283);
   U5937 : AOI222_X1 port map( A1 => n16202, A2 => n5288, B1 => n15609, B2 => 
                           n5293, C1 => n16201, C2 => n5289, ZN => n6208);
   U5938 : AOI222_X1 port map( A1 => n16208, A2 => n5288, B1 => n15610, B2 => 
                           n5293, C1 => n16207, C2 => n5289, ZN => n6133);
   U5939 : AOI222_X1 port map( A1 => n16280, A2 => n5288, B1 => n15601, B2 => 
                           n5293, C1 => n16279, C2 => n5289, ZN => n6808);
   U5940 : AOI222_X1 port map( A1 => n54260, A2 => n62128, B1 => n54236, B2 => 
                           n61835, C1 => n54513, C2 => n62130, ZN => n6761);
   U5941 : AOI222_X1 port map( A1 => n54259, A2 => n62128, B1 => n54235, B2 => 
                           n61835, C1 => n54514, C2 => n62130, ZN => n6686);
   U5942 : AOI222_X1 port map( A1 => n54258, A2 => n62128, B1 => n54234, B2 => 
                           n61835, C1 => n54515, C2 => n62130, ZN => n6611);
   U5943 : AOI222_X1 port map( A1 => n54257, A2 => n62128, B1 => n54233, B2 => 
                           n61835, C1 => n54516, C2 => n62130, ZN => n6536);
   U5944 : AOI222_X1 port map( A1 => n54256, A2 => n62128, B1 => n54232, B2 => 
                           n61835, C1 => n54517, C2 => n62130, ZN => n6461);
   U5945 : AOI222_X1 port map( A1 => n54255, A2 => n62128, B1 => n54231, B2 => 
                           n61835, C1 => n54518, C2 => n62130, ZN => n6386);
   U5946 : AOI222_X1 port map( A1 => n54254, A2 => n62128, B1 => n54230, B2 => 
                           n61835, C1 => n54519, C2 => n62130, ZN => n6311);
   U5947 : AOI222_X1 port map( A1 => n54253, A2 => n62128, B1 => n54229, B2 => 
                           n61835, C1 => n54520, C2 => n62130, ZN => n6236);
   U5948 : AOI222_X1 port map( A1 => n54252, A2 => n62128, B1 => n54228, B2 => 
                           n61835, C1 => n54521, C2 => n62130, ZN => n6161);
   U5949 : AOI222_X1 port map( A1 => n54265, A2 => n62129, B1 => n54241, B2 => 
                           n61834, C1 => n54524, C2 => n62131, ZN => n7136);
   U5950 : AOI222_X1 port map( A1 => n54264, A2 => n62129, B1 => n54240, B2 => 
                           n61834, C1 => n54525, C2 => n62131, ZN => n7061);
   U5951 : AOI222_X1 port map( A1 => n54262, A2 => n62128, B1 => n54238, B2 => 
                           n61835, C1 => n54511, C2 => n62130, ZN => n6911);
   U5952 : AOI222_X1 port map( A1 => n54261, A2 => n62128, B1 => n54237, B2 => 
                           n61835, C1 => n54512, C2 => n62130, ZN => n6836);
   U5953 : AOI222_X1 port map( A1 => n54267, A2 => n62129, B1 => n54243, B2 => 
                           n61834, C1 => n54508, C2 => n62131, ZN => n7286);
   U5954 : AOI222_X1 port map( A1 => n54275, A2 => n62129, B1 => n54251, B2 => 
                           n61834, C1 => n54527, C2 => n62131, ZN => n7913);
   U5955 : AOI222_X1 port map( A1 => n54274, A2 => n62129, B1 => n54250, B2 => 
                           n61834, C1 => n54504, C2 => n62131, ZN => n7811);
   U5956 : AOI222_X1 port map( A1 => n54273, A2 => n62129, B1 => n54249, B2 => 
                           n61834, C1 => n54505, C2 => n62131, ZN => n7736);
   U5957 : AOI222_X1 port map( A1 => n54272, A2 => n62129, B1 => n54248, B2 => 
                           n61834, C1 => n54506, C2 => n62131, ZN => n7661);
   U5958 : AOI222_X1 port map( A1 => n54271, A2 => n62129, B1 => n54247, B2 => 
                           n61834, C1 => n54507, C2 => n62131, ZN => n7586);
   U5959 : AOI222_X1 port map( A1 => n54270, A2 => n62129, B1 => n54246, B2 => 
                           n61834, C1 => n54509, C2 => n62131, ZN => n7511);
   U5960 : AOI222_X1 port map( A1 => n54269, A2 => n62129, B1 => n54245, B2 => 
                           n61834, C1 => n54510, C2 => n62131, ZN => n7436);
   U5961 : AOI222_X1 port map( A1 => n54268, A2 => n62129, B1 => n54244, B2 => 
                           n61834, C1 => n54522, C2 => n62131, ZN => n7361);
   U5962 : AOI222_X1 port map( A1 => n54266, A2 => n62129, B1 => n54242, B2 => 
                           n61834, C1 => n54523, C2 => n62131, ZN => n7211);
   U5963 : AOI222_X1 port map( A1 => n54263, A2 => n62128, B1 => n54239, B2 => 
                           n61835, C1 => n54526, C2 => n62130, ZN => n6986);
   U5964 : AOI222_X1 port map( A1 => n2799, A2 => n61781, B1 => n2823, B2 => 
                           n61778, C1 => n53712, C2 => n61775, ZN => n6777);
   U5965 : AOI222_X1 port map( A1 => n2798, A2 => n61781, B1 => n2822, B2 => 
                           n61778, C1 => n53711, C2 => n61775, ZN => n6702);
   U5966 : AOI222_X1 port map( A1 => n2797, A2 => n61781, B1 => n2821, B2 => 
                           n61778, C1 => n53710, C2 => n61775, ZN => n6627);
   U5967 : AOI222_X1 port map( A1 => n2796, A2 => n61781, B1 => n2820, B2 => 
                           n61778, C1 => n53709, C2 => n61775, ZN => n6552);
   U5968 : AOI222_X1 port map( A1 => n52772, A2 => n61742, B1 => n54570, B2 => 
                           n61739, C1 => n52788, C2 => n61735, ZN => n6485);
   U5969 : AOI222_X1 port map( A1 => n2795, A2 => n61781, B1 => n2819, B2 => 
                           n61778, C1 => n53708, C2 => n61775, ZN => n6477);
   U5970 : AOI222_X1 port map( A1 => n52771, A2 => n61741, B1 => n54571, B2 => 
                           n61739, C1 => n52787, C2 => n61735, ZN => n6410);
   U5971 : AOI222_X1 port map( A1 => n2794, A2 => n61781, B1 => n2818, B2 => 
                           n61778, C1 => n53707, C2 => n61775, ZN => n6402);
   U5972 : AOI222_X1 port map( A1 => n52770, A2 => n61741, B1 => n54572, B2 => 
                           n61739, C1 => n52786, C2 => n61735, ZN => n6335);
   U5973 : AOI222_X1 port map( A1 => n2793, A2 => n61781, B1 => n2817, B2 => 
                           n61778, C1 => n53706, C2 => n61775, ZN => n6327);
   U5974 : AOI222_X1 port map( A1 => n52769, A2 => n61741, B1 => n54573, B2 => 
                           n61739, C1 => n52785, C2 => n61735, ZN => n6260);
   U5975 : AOI222_X1 port map( A1 => n2792, A2 => n61781, B1 => n2816, B2 => 
                           n61778, C1 => n53705, C2 => n61775, ZN => n6252);
   U5976 : AOI222_X1 port map( A1 => n52768, A2 => n61741, B1 => n54574, B2 => 
                           n61738, C1 => n52784, C2 => n61735, ZN => n6185);
   U5977 : AOI222_X1 port map( A1 => n2791, A2 => n61781, B1 => n2815, B2 => 
                           n61778, C1 => n53704, C2 => n61775, ZN => n6177);
   U5978 : AOI222_X1 port map( A1 => n2804, A2 => n61780, B1 => n2828, B2 => 
                           n61777, C1 => n53717, C2 => n61774, ZN => n7152);
   U5979 : AOI222_X1 port map( A1 => n2803, A2 => n61780, B1 => n2827, B2 => 
                           n61777, C1 => n53716, C2 => n61774, ZN => n7077);
   U5980 : AOI222_X1 port map( A1 => n2801, A2 => n61781, B1 => n2825, B2 => 
                           n61778, C1 => n53714, C2 => n61775, ZN => n6927);
   U5981 : AOI222_X1 port map( A1 => n2800, A2 => n61781, B1 => n2824, B2 => 
                           n61778, C1 => n53713, C2 => n61775, ZN => n6852);
   U5982 : AOI222_X1 port map( A1 => n52767, A2 => n61741, B1 => n51783, B2 => 
                           n61738, C1 => n61737, C2 => n3939, ZN => n6110);
   U5983 : AOI222_X1 port map( A1 => n52766, A2 => n61741, B1 => n51782, B2 => 
                           n61738, C1 => n61737, C2 => n3938, ZN => n6004);
   U5984 : AOI222_X1 port map( A1 => n52765, A2 => n61741, B1 => n51781, B2 => 
                           n61738, C1 => n61737, C2 => n3937, ZN => n5929);
   U5985 : AOI222_X1 port map( A1 => n52764, A2 => n61741, B1 => n51780, B2 => 
                           n61738, C1 => n61737, C2 => n3936, ZN => n5854);
   U5986 : AOI222_X1 port map( A1 => n52763, A2 => n61741, B1 => n51779, B2 => 
                           n61738, C1 => n61737, C2 => n3935, ZN => n5779);
   U5987 : AOI222_X1 port map( A1 => n52762, A2 => n61741, B1 => n51778, B2 => 
                           n61738, C1 => n52238, C2 => n61735, ZN => n5704);
   U5988 : AOI222_X1 port map( A1 => n52761, A2 => n61741, B1 => n51777, B2 => 
                           n61738, C1 => n52237, C2 => n61735, ZN => n5629);
   U5989 : AOI222_X1 port map( A1 => n52760, A2 => n61741, B1 => n51776, B2 => 
                           n61738, C1 => n52236, C2 => n61736, ZN => n5551);
   U5990 : AOI222_X1 port map( A1 => n2806, A2 => n61780, B1 => n2830, B2 => 
                           n61777, C1 => n53719, C2 => n61774, ZN => n7302);
   U5991 : AOI222_X1 port map( A1 => n61743, A2 => n52783, B1 => n54575, B2 => 
                           n61738, C1 => n52807, C2 => n61735, ZN => n7942);
   U5992 : AOI222_X1 port map( A1 => n2814, A2 => n61780, B1 => n2838, B2 => 
                           n61777, C1 => n53727, C2 => n61774, ZN => n7933);
   U5993 : AOI222_X1 port map( A1 => n61743, A2 => n52782, B1 => n54563, B2 => 
                           n61738, C1 => n52806, C2 => n61737, ZN => n7835);
   U5994 : AOI222_X1 port map( A1 => n2813, A2 => n61780, B1 => n2837, B2 => 
                           n61777, C1 => n53726, C2 => n61774, ZN => n7827);
   U5995 : AOI222_X1 port map( A1 => n61743, A2 => n52781, B1 => n54564, B2 => 
                           n61738, C1 => n52805, C2 => n61737, ZN => n7760);
   U5996 : AOI222_X1 port map( A1 => n2812, A2 => n61780, B1 => n2836, B2 => 
                           n61777, C1 => n53725, C2 => n61774, ZN => n7752);
   U5997 : AOI222_X1 port map( A1 => n61743, A2 => n52780, B1 => n61739, B2 => 
                           n59676, C1 => n52804, C2 => n61737, ZN => n7685);
   U5998 : AOI222_X1 port map( A1 => n2811, A2 => n61780, B1 => n2835, B2 => 
                           n61777, C1 => n53724, C2 => n61774, ZN => n7677);
   U5999 : AOI222_X1 port map( A1 => n2810, A2 => n61780, B1 => n2834, B2 => 
                           n61777, C1 => n53723, C2 => n61774, ZN => n7602);
   U6000 : AOI222_X1 port map( A1 => n2809, A2 => n61780, B1 => n2833, B2 => 
                           n61777, C1 => n53722, C2 => n61774, ZN => n7527);
   U6001 : AOI222_X1 port map( A1 => n2808, A2 => n61780, B1 => n2832, B2 => 
                           n61777, C1 => n53721, C2 => n61774, ZN => n7452);
   U6002 : AOI222_X1 port map( A1 => n2807, A2 => n61780, B1 => n2831, B2 => 
                           n61777, C1 => n53720, C2 => n61774, ZN => n7377);
   U6003 : AOI222_X1 port map( A1 => n2805, A2 => n61780, B1 => n2829, B2 => 
                           n61777, C1 => n53718, C2 => n61774, ZN => n7227);
   U6004 : AOI222_X1 port map( A1 => n61266, A2 => n52772, B1 => n61263, B2 => 
                           n54570, C1 => n61260, C2 => n52788, ZN => n9054);
   U6005 : AOI222_X1 port map( A1 => n61266, A2 => n52771, B1 => n61262, B2 => 
                           n54571, C1 => n61259, C2 => n52787, ZN => n8979);
   U6006 : AOI222_X1 port map( A1 => n61266, A2 => n52770, B1 => n61262, B2 => 
                           n54572, C1 => n61259, C2 => n52786, ZN => n8904);
   U6007 : AOI222_X1 port map( A1 => n61266, A2 => n52769, B1 => n61262, B2 => 
                           n54573, C1 => n61259, C2 => n52785, ZN => n8829);
   U6008 : AOI222_X1 port map( A1 => n61266, A2 => n52768, B1 => n61262, B2 => 
                           n54574, C1 => n61259, C2 => n52784, ZN => n8754);
   U6009 : AOI222_X1 port map( A1 => n61267, A2 => n52767, B1 => n61262, B2 => 
                           n51783, C1 => n61259, C2 => n3939, ZN => n8679);
   U6010 : AOI222_X1 port map( A1 => n61267, A2 => n52766, B1 => n61262, B2 => 
                           n51782, C1 => n61259, C2 => n3938, ZN => n8604);
   U6011 : AOI222_X1 port map( A1 => n61267, A2 => n52765, B1 => n61262, B2 => 
                           n51781, C1 => n61259, C2 => n3937, ZN => n8529);
   U6012 : AOI222_X1 port map( A1 => n61267, A2 => n52764, B1 => n61262, B2 => 
                           n51780, C1 => n61259, C2 => n3936, ZN => n8454);
   U6013 : AOI222_X1 port map( A1 => n61267, A2 => n52763, B1 => n61262, B2 => 
                           n51779, C1 => n61259, C2 => n3935, ZN => n8379);
   U6014 : AOI222_X1 port map( A1 => n61267, A2 => n52762, B1 => n61262, B2 => 
                           n51778, C1 => n61259, C2 => n52238, ZN => n8304);
   U6015 : AOI222_X1 port map( A1 => n61267, A2 => n52761, B1 => n61262, B2 => 
                           n51777, C1 => n61259, C2 => n52237, ZN => n8229);
   U6016 : AOI222_X1 port map( A1 => n61267, A2 => n52760, B1 => n61262, B2 => 
                           n51776, C1 => n61259, C2 => n52236, ZN => n8151);
   U6017 : AOI222_X1 port map( A1 => n61265, A2 => n52783, B1 => n61264, B2 => 
                           n54575, C1 => n61261, C2 => n52807, ZN => n15071);
   U6018 : AOI222_X1 port map( A1 => n61265, A2 => n52782, B1 => n61264, B2 => 
                           n54563, C1 => n61261, C2 => n52806, ZN => n14964);
   U6019 : AOI222_X1 port map( A1 => n61265, A2 => n52781, B1 => n61264, B2 => 
                           n54564, C1 => n61261, C2 => n52805, ZN => n14889);
   U6020 : AOI222_X1 port map( A1 => n2802, A2 => n61781, B1 => n2826, B2 => 
                           n61778, C1 => n53715, C2 => n61775, ZN => n7002);
   U6021 : AOI222_X1 port map( A1 => n61470, A2 => n54383, B1 => n61467, B2 => 
                           n54558, C1 => n61464, C2 => n54407, ZN => n9623);
   U6022 : AOI222_X1 port map( A1 => n61470, A2 => n54382, B1 => n61467, B2 => 
                           n54543, C1 => n61464, C2 => n54406, ZN => n9532);
   U6023 : AOI222_X1 port map( A1 => n61470, A2 => n54381, B1 => n61467, B2 => 
                           n54544, C1 => n61464, C2 => n54405, ZN => n9457);
   U6024 : AOI222_X1 port map( A1 => n61470, A2 => n54380, B1 => n61467, B2 => 
                           n54545, C1 => n61464, C2 => n54404, ZN => n9382);
   U6025 : AOI222_X1 port map( A1 => n61470, A2 => n54379, B1 => n61467, B2 => 
                           n54546, C1 => n61464, C2 => n54403, ZN => n9243);
   U6026 : AOI222_X1 port map( A1 => n61470, A2 => n54378, B1 => n61467, B2 => 
                           n54547, C1 => n61464, C2 => n54402, ZN => n9168);
   U6027 : AOI222_X1 port map( A1 => n61470, A2 => n54377, B1 => n61467, B2 => 
                           n54548, C1 => n61464, C2 => n54401, ZN => n9093);
   U6028 : AOI222_X1 port map( A1 => n61470, A2 => n54376, B1 => n61467, B2 => 
                           n54549, C1 => n61464, C2 => n54400, ZN => n9018);
   U6029 : AOI222_X1 port map( A1 => n61470, A2 => n54375, B1 => n61466, B2 => 
                           n54550, C1 => n61463, C2 => n54399, ZN => n8943);
   U6030 : AOI222_X1 port map( A1 => n61470, A2 => n54374, B1 => n61466, B2 => 
                           n54551, C1 => n61463, C2 => n54398, ZN => n8868);
   U6031 : AOI222_X1 port map( A1 => n61470, A2 => n54373, B1 => n61466, B2 => 
                           n54552, C1 => n61463, C2 => n54397, ZN => n8793);
   U6032 : AOI222_X1 port map( A1 => n61470, A2 => n54372, B1 => n61466, B2 => 
                           n54553, C1 => n61463, C2 => n54396, ZN => n8718);
   U6033 : AOI222_X1 port map( A1 => n54531, A2 => n61742, B1 => n61739, B2 => 
                           n59684, C1 => n52792, C2 => n61735, ZN => n6785);
   U6034 : AOI222_X1 port map( A1 => n54532, A2 => n61742, B1 => n61739, B2 => 
                           n59685, C1 => n52791, C2 => n61735, ZN => n6710);
   U6035 : AOI222_X1 port map( A1 => n54533, A2 => n61742, B1 => n61739, B2 => 
                           n59686, C1 => n52790, C2 => n61735, ZN => n6635);
   U6036 : AOI222_X1 port map( A1 => n54534, A2 => n61742, B1 => n61739, B2 => 
                           n59687, C1 => n52789, C2 => n61735, ZN => n6560);
   U6037 : AOI222_X1 port map( A1 => n61742, A2 => n52773, B1 => n61740, B2 => 
                           n59675, C1 => n52797, C2 => n61736, ZN => n7160);
   U6038 : AOI222_X1 port map( A1 => n54535, A2 => n61742, B1 => n61740, B2 => 
                           n59681, C1 => n52796, C2 => n61736, ZN => n7085);
   U6039 : AOI222_X1 port map( A1 => n54529, A2 => n61742, B1 => n61739, B2 => 
                           n59682, C1 => n52794, C2 => n61736, ZN => n6935);
   U6040 : AOI222_X1 port map( A1 => n54530, A2 => n61742, B1 => n61739, B2 => 
                           n59683, C1 => n52793, C2 => n61736, ZN => n6860);
   U6041 : AOI222_X1 port map( A1 => n530, A2 => n61869, B1 => n538, B2 => 
                           n61698, C1 => n52275, C2 => n59645, ZN => n6060);
   U6042 : AOI222_X1 port map( A1 => n61876, A2 => n4264, B1 => n52358, B2 => 
                           n61710, C1 => n52315, C2 => n61712, ZN => n6046);
   U6043 : AOI222_X1 port map( A1 => n51735, A2 => n61836, B1 => n1646, B2 => 
                           n61690, C1 => n59648, C2 => n4035, ZN => n6076);
   U6044 : AOI222_X1 port map( A1 => n529, A2 => n61869, B1 => n537, B2 => 
                           n61698, C1 => n52274, C2 => n59645, ZN => n5968);
   U6045 : AOI222_X1 port map( A1 => n61876, A2 => n4263, B1 => n52357, B2 => 
                           n61710, C1 => n52314, C2 => n61712, ZN => n5960);
   U6046 : AOI222_X1 port map( A1 => n51734, A2 => n61836, B1 => n1645, B2 => 
                           n61690, C1 => n59648, C2 => n4034, ZN => n5980);
   U6047 : AOI222_X1 port map( A1 => n528, A2 => n61869, B1 => n536, B2 => 
                           n61698, C1 => n52273, C2 => n59645, ZN => n5893);
   U6048 : AOI222_X1 port map( A1 => n61876, A2 => n4262, B1 => n52356, B2 => 
                           n61710, C1 => n52313, C2 => n61712, ZN => n5885);
   U6049 : AOI222_X1 port map( A1 => n51733, A2 => n61836, B1 => n1644, B2 => 
                           n61690, C1 => n59648, C2 => n4033, ZN => n5905);
   U6050 : AOI222_X1 port map( A1 => n527, A2 => n61869, B1 => n535, B2 => 
                           n61698, C1 => n52272, C2 => n59645, ZN => n5818);
   U6051 : AOI222_X1 port map( A1 => n61876, A2 => n4261, B1 => n52355, B2 => 
                           n61710, C1 => n52312, C2 => n61712, ZN => n5810);
   U6052 : AOI222_X1 port map( A1 => n51732, A2 => n61836, B1 => n1643, B2 => 
                           n61690, C1 => n59648, C2 => n4032, ZN => n5830);
   U6053 : AOI222_X1 port map( A1 => n526, A2 => n61869, B1 => n534, B2 => 
                           n61698, C1 => n52271, C2 => n59645, ZN => n5743);
   U6054 : AOI222_X1 port map( A1 => n61876, A2 => n4260, B1 => n52354, B2 => 
                           n61710, C1 => n52311, C2 => n61712, ZN => n5735);
   U6055 : AOI222_X1 port map( A1 => n51731, A2 => n61836, B1 => n1642, B2 => 
                           n61690, C1 => n59648, C2 => n4031, ZN => n5755);
   U6056 : AOI222_X1 port map( A1 => n525, A2 => n61869, B1 => n533, B2 => 
                           n61698, C1 => n52270, C2 => n59645, ZN => n5668);
   U6057 : AOI222_X1 port map( A1 => n61876, A2 => n4259, B1 => n52353, B2 => 
                           n61710, C1 => n52310, C2 => n61712, ZN => n5660);
   U6058 : AOI222_X1 port map( A1 => n51730, A2 => n61836, B1 => n1641, B2 => 
                           n61690, C1 => n59648, C2 => n4030, ZN => n5680);
   U6059 : AOI222_X1 port map( A1 => n524, A2 => n61869, B1 => n532, B2 => 
                           n61698, C1 => n52269, C2 => n59645, ZN => n5593);
   U6060 : AOI222_X1 port map( A1 => n61876, A2 => n4258, B1 => n52352, B2 => 
                           n61710, C1 => n52309, C2 => n61712, ZN => n5585);
   U6061 : AOI222_X1 port map( A1 => n51729, A2 => n61836, B1 => n1640, B2 => 
                           n61690, C1 => n59648, C2 => n4029, ZN => n5605);
   U6062 : AOI222_X1 port map( A1 => n523, A2 => n61869, B1 => n531, B2 => 
                           n61698, C1 => n52268, C2 => n59645, ZN => n5461);
   U6063 : AOI222_X1 port map( A1 => n61876, A2 => n4257, B1 => n52351, B2 => 
                           n61710, C1 => n52308, C2 => n61712, ZN => n5442);
   U6064 : AOI222_X1 port map( A1 => n51728, A2 => n61836, B1 => n1639, B2 => 
                           n61690, C1 => n59648, C2 => n4028, ZN => n5486);
   U6065 : AOI222_X1 port map( A1 => n61742, A2 => n52775, B1 => n61739, B2 => 
                           n59673, C1 => n52799, C2 => n61736, ZN => n7310);
   U6066 : AOI222_X1 port map( A1 => n61743, A2 => n52779, B1 => n61740, B2 => 
                           n59677, C1 => n52803, C2 => n61736, ZN => n7610);
   U6067 : AOI222_X1 port map( A1 => n61743, A2 => n52778, B1 => n61740, B2 => 
                           n59678, C1 => n52802, C2 => n61736, ZN => n7535);
   U6068 : AOI222_X1 port map( A1 => n61743, A2 => n52777, B1 => n61740, B2 => 
                           n59679, C1 => n52801, C2 => n61736, ZN => n7460);
   U6069 : AOI222_X1 port map( A1 => n61743, A2 => n52776, B1 => n61740, B2 => 
                           n59680, C1 => n52800, C2 => n61736, ZN => n7385);
   U6070 : AOI222_X1 port map( A1 => n61742, A2 => n52774, B1 => n61740, B2 => 
                           n59674, C1 => n52798, C2 => n61736, ZN => n7235);
   U6071 : AOI222_X1 port map( A1 => n61469, A2 => n54387, B1 => n61467, B2 => 
                           n59718, C1 => n61464, C2 => n54411, ZN => n14403);
   U6072 : AOI222_X1 port map( A1 => n61265, A2 => n52775, B1 => n61263, B2 => 
                           n59673, C1 => n61260, C2 => n52799, ZN => n14439);
   U6073 : AOI222_X1 port map( A1 => n61469, A2 => n54386, B1 => n61467, B2 => 
                           n59719, C1 => n61464, C2 => n54410, ZN => n9912);
   U6074 : AOI222_X1 port map( A1 => n61265, A2 => n52774, B1 => n61263, B2 => 
                           n59674, C1 => n61260, C2 => n52798, ZN => n14364);
   U6075 : AOI222_X1 port map( A1 => n61469, A2 => n54385, B1 => n61467, B2 => 
                           n59720, C1 => n61464, C2 => n54409, ZN => n9837);
   U6076 : AOI222_X1 port map( A1 => n61265, A2 => n52773, B1 => n61263, B2 => 
                           n59675, C1 => n61260, C2 => n52797, ZN => n9873);
   U6077 : AOI222_X1 port map( A1 => n61469, A2 => n54384, B1 => n61467, B2 => 
                           n59721, C1 => n61464, C2 => n54408, ZN => n9698);
   U6078 : AOI222_X1 port map( A1 => n61265, A2 => n54535, B1 => n61263, B2 => 
                           n59681, C1 => n61260, C2 => n52796, ZN => n9734);
   U6079 : AOI222_X1 port map( A1 => n61266, A2 => n54528, B1 => n61263, B2 => 
                           n59688, C1 => n61260, C2 => n52795, ZN => n9659);
   U6080 : AOI222_X1 port map( A1 => n61266, A2 => n54529, B1 => n61263, B2 => 
                           n59682, C1 => n61260, C2 => n52794, ZN => n9568);
   U6081 : AOI222_X1 port map( A1 => n61266, A2 => n54530, B1 => n61263, B2 => 
                           n59683, C1 => n61260, C2 => n52793, ZN => n9493);
   U6082 : AOI222_X1 port map( A1 => n61266, A2 => n54531, B1 => n61263, B2 => 
                           n59684, C1 => n61260, C2 => n52792, ZN => n9418);
   U6083 : AOI222_X1 port map( A1 => n61266, A2 => n54532, B1 => n61263, B2 => 
                           n59685, C1 => n61260, C2 => n52791, ZN => n9279);
   U6084 : AOI222_X1 port map( A1 => n61266, A2 => n54533, B1 => n61263, B2 => 
                           n59686, C1 => n61260, C2 => n52790, ZN => n9204);
   U6085 : AOI222_X1 port map( A1 => n61266, A2 => n54534, B1 => n61263, B2 => 
                           n59687, C1 => n61260, C2 => n52789, ZN => n9129);
   U6086 : AOI222_X1 port map( A1 => n61471, A2 => n4083, B1 => n61466, B2 => 
                           n4091, C1 => n61463, C2 => n4099, ZN => n8643);
   U6087 : AOI222_X1 port map( A1 => n61471, A2 => n4082, B1 => n61466, B2 => 
                           n4090, C1 => n61463, C2 => n4098, ZN => n8568);
   U6088 : AOI222_X1 port map( A1 => n61471, A2 => n4081, B1 => n61466, B2 => 
                           n4089, C1 => n61463, C2 => n4097, ZN => n8493);
   U6089 : AOI222_X1 port map( A1 => n61471, A2 => n4080, B1 => n61466, B2 => 
                           n4088, C1 => n61463, C2 => n4096, ZN => n8418);
   U6090 : AOI222_X1 port map( A1 => n61471, A2 => n4079, B1 => n61466, B2 => 
                           n4087, C1 => n61463, C2 => n4095, ZN => n8343);
   U6091 : AOI222_X1 port map( A1 => n61471, A2 => n4078, B1 => n61466, B2 => 
                           n4086, C1 => n61463, C2 => n4094, ZN => n8268);
   U6092 : AOI222_X1 port map( A1 => n61471, A2 => n4077, B1 => n61466, B2 => 
                           n4085, C1 => n61463, C2 => n4093, ZN => n8193);
   U6093 : AOI222_X1 port map( A1 => n61471, A2 => n4076, B1 => n61466, B2 => 
                           n4084, C1 => n61463, C2 => n4092, ZN => n8047);
   U6094 : AOI222_X1 port map( A1 => n61469, A2 => n54395, B1 => n61468, B2 => 
                           n59722, C1 => n61465, C2 => n54419, ZN => n15025);
   U6095 : AOI222_X1 port map( A1 => n61469, A2 => n54394, B1 => n61468, B2 => 
                           n59723, C1 => n61465, C2 => n54418, ZN => n14928);
   U6096 : AOI222_X1 port map( A1 => n61469, A2 => n54393, B1 => n61468, B2 => 
                           n59724, C1 => n61465, C2 => n54417, ZN => n14853);
   U6097 : AOI222_X1 port map( A1 => n61469, A2 => n54392, B1 => n61468, B2 => 
                           n59725, C1 => n61465, C2 => n54416, ZN => n14778);
   U6098 : AOI222_X1 port map( A1 => n61265, A2 => n52780, B1 => n61264, B2 => 
                           n59676, C1 => n61261, C2 => n52804, ZN => n14814);
   U6099 : AOI222_X1 port map( A1 => n61469, A2 => n54391, B1 => n61468, B2 => 
                           n59726, C1 => n61465, C2 => n54415, ZN => n14703);
   U6100 : AOI222_X1 port map( A1 => n61265, A2 => n52779, B1 => n61264, B2 => 
                           n59677, C1 => n61261, C2 => n52803, ZN => n14739);
   U6101 : AOI222_X1 port map( A1 => n61469, A2 => n54390, B1 => n61468, B2 => 
                           n59727, C1 => n61465, C2 => n54414, ZN => n14628);
   U6102 : AOI222_X1 port map( A1 => n61265, A2 => n52778, B1 => n61264, B2 => 
                           n59678, C1 => n61261, C2 => n52802, ZN => n14664);
   U6103 : AOI222_X1 port map( A1 => n61469, A2 => n54389, B1 => n61468, B2 => 
                           n59728, C1 => n61465, C2 => n54413, ZN => n14553);
   U6104 : AOI222_X1 port map( A1 => n61265, A2 => n52777, B1 => n61264, B2 => 
                           n59679, C1 => n61261, C2 => n52801, ZN => n14589);
   U6105 : AOI222_X1 port map( A1 => n61469, A2 => n54388, B1 => n61468, B2 => 
                           n59729, C1 => n61465, C2 => n54412, ZN => n14478);
   U6106 : AOI222_X1 port map( A1 => n61265, A2 => n52776, B1 => n61264, B2 => 
                           n59680, C1 => n61261, C2 => n52800, ZN => n14514);
   U6107 : AOI222_X1 port map( A1 => n54528, A2 => n61742, B1 => n61739, B2 => 
                           n59688, C1 => n52795, C2 => n61736, ZN => n7010);
   U6108 : NOR4_X1 port map( A1 => n6718, A2 => n6719, A3 => n6720, A4 => n6721
                           , ZN => n6717);
   U6109 : OAI221_X1 port map( B1 => n2235, B2 => n6021, C1 => n2257, C2 => 
                           n61730, A => n6724, ZN => n6719);
   U6110 : OAI221_X1 port map( B1 => n61718, B2 => n1713, C1 => n52936, C2 => 
                           n61910, A => n6722, ZN => n6721);
   U6111 : OAI221_X1 port map( B1 => n896, B2 => n6018, C1 => n872, C2 => 
                           n61734, A => n6723, ZN => n6720);
   U6112 : NOR4_X1 port map( A1 => n6643, A2 => n6644, A3 => n6645, A4 => n6646
                           , ZN => n6642);
   U6113 : OAI221_X1 port map( B1 => n2220, B2 => n6021, C1 => n2256, C2 => 
                           n61730, A => n6649, ZN => n6644);
   U6114 : OAI221_X1 port map( B1 => n61718, B2 => n1712, C1 => n52935, C2 => 
                           n61910, A => n6647, ZN => n6646);
   U6115 : OAI221_X1 port map( B1 => n895, B2 => n6018, C1 => n871, C2 => 
                           n61734, A => n6648, ZN => n6645);
   U6116 : NOR4_X1 port map( A1 => n6568, A2 => n6569, A3 => n6570, A4 => n6571
                           , ZN => n6567);
   U6117 : OAI221_X1 port map( B1 => n2219, B2 => n6021, C1 => n2255, C2 => 
                           n61730, A => n6574, ZN => n6569);
   U6118 : OAI221_X1 port map( B1 => n61718, B2 => n1711, C1 => n52934, C2 => 
                           n61910, A => n6572, ZN => n6571);
   U6119 : OAI221_X1 port map( B1 => n894, B2 => n6018, C1 => n870, C2 => 
                           n61734, A => n6573, ZN => n6570);
   U6120 : NOR4_X1 port map( A1 => n6493, A2 => n6494, A3 => n6495, A4 => n6496
                           , ZN => n6492);
   U6121 : OAI221_X1 port map( B1 => n2218, B2 => n6021, C1 => n2254, C2 => 
                           n61730, A => n6499, ZN => n6494);
   U6122 : OAI221_X1 port map( B1 => n61718, B2 => n1710, C1 => n52933, C2 => 
                           n61910, A => n6497, ZN => n6496);
   U6123 : OAI221_X1 port map( B1 => n893, B2 => n6018, C1 => n869, C2 => 
                           n61734, A => n6498, ZN => n6495);
   U6124 : NOR4_X1 port map( A1 => n6418, A2 => n6419, A3 => n6420, A4 => n6421
                           , ZN => n6417);
   U6125 : OAI221_X1 port map( B1 => n2217, B2 => n6021, C1 => n2253, C2 => 
                           n61730, A => n6424, ZN => n6419);
   U6126 : OAI221_X1 port map( B1 => n61718, B2 => n1709, C1 => n52932, C2 => 
                           n61910, A => n6422, ZN => n6421);
   U6127 : OAI221_X1 port map( B1 => n892, B2 => n6018, C1 => n868, C2 => 
                           n61734, A => n6423, ZN => n6420);
   U6128 : NOR4_X1 port map( A1 => n6343, A2 => n6344, A3 => n6345, A4 => n6346
                           , ZN => n6342);
   U6129 : OAI221_X1 port map( B1 => n2216, B2 => n6021, C1 => n2252, C2 => 
                           n61730, A => n6349, ZN => n6344);
   U6130 : OAI221_X1 port map( B1 => n61718, B2 => n1708, C1 => n52931, C2 => 
                           n61910, A => n6347, ZN => n6346);
   U6131 : OAI221_X1 port map( B1 => n891, B2 => n6018, C1 => n867, C2 => 
                           n61734, A => n6348, ZN => n6345);
   U6132 : NOR4_X1 port map( A1 => n6268, A2 => n6269, A3 => n6270, A4 => n6271
                           , ZN => n6267);
   U6133 : OAI221_X1 port map( B1 => n2215, B2 => n6021, C1 => n2251, C2 => 
                           n61730, A => n6274, ZN => n6269);
   U6134 : OAI221_X1 port map( B1 => n61718, B2 => n1707, C1 => n52930, C2 => 
                           n61910, A => n6272, ZN => n6271);
   U6135 : OAI221_X1 port map( B1 => n890, B2 => n6018, C1 => n866, C2 => 
                           n61734, A => n6273, ZN => n6270);
   U6136 : NOR4_X1 port map( A1 => n6193, A2 => n6194, A3 => n6195, A4 => n6196
                           , ZN => n6192);
   U6137 : OAI221_X1 port map( B1 => n2214, B2 => n6021, C1 => n2250, C2 => 
                           n61730, A => n6199, ZN => n6194);
   U6138 : OAI221_X1 port map( B1 => n61718, B2 => n1706, C1 => n52929, C2 => 
                           n61910, A => n6197, ZN => n6196);
   U6139 : OAI221_X1 port map( B1 => n889, B2 => n6018, C1 => n865, C2 => 
                           n61734, A => n6198, ZN => n6195);
   U6140 : NOR4_X1 port map( A1 => n6118, A2 => n6119, A3 => n6120, A4 => n6121
                           , ZN => n6117);
   U6141 : OAI221_X1 port map( B1 => n2213, B2 => n6021, C1 => n2249, C2 => 
                           n61730, A => n6124, ZN => n6119);
   U6142 : OAI221_X1 port map( B1 => n61718, B2 => n1705, C1 => n52928, C2 => 
                           n61910, A => n6122, ZN => n6121);
   U6143 : OAI221_X1 port map( B1 => n888, B2 => n6018, C1 => n864, C2 => 
                           n61734, A => n6123, ZN => n6120);
   U6144 : NOR4_X1 port map( A1 => n7093, A2 => n7094, A3 => n7095, A4 => n7096
                           , ZN => n7092);
   U6145 : OAI221_X1 port map( B1 => n2239, B2 => n61727, C1 => n2261, C2 => 
                           n61729, A => n7099, ZN => n7094);
   U6146 : OAI221_X1 port map( B1 => n61717, B2 => n1718, C1 => n52941, C2 => 
                           n61909, A => n7097, ZN => n7096);
   U6147 : OAI221_X1 port map( B1 => n901, B2 => n61731, C1 => n877, C2 => 
                           n61733, A => n7098, ZN => n7095);
   U6148 : NOR4_X1 port map( A1 => n7018, A2 => n7019, A3 => n7020, A4 => n7021
                           , ZN => n7017);
   U6149 : OAI221_X1 port map( B1 => n2075, B2 => n61727, C1 => n2077, C2 => 
                           n61729, A => n7024, ZN => n7019);
   U6150 : OAI221_X1 port map( B1 => n61717, B2 => n1717, C1 => n52940, C2 => 
                           n61909, A => n7022, ZN => n7021);
   U6151 : OAI221_X1 port map( B1 => n900, B2 => n61731, C1 => n876, C2 => 
                           n61733, A => n7023, ZN => n7020);
   U6152 : NOR4_X1 port map( A1 => n6868, A2 => n6869, A3 => n6870, A4 => n6871
                           , ZN => n6867);
   U6153 : OAI221_X1 port map( B1 => n2237, B2 => n6021, C1 => n2259, C2 => 
                           n61730, A => n6874, ZN => n6869);
   U6154 : OAI221_X1 port map( B1 => n61718, B2 => n1715, C1 => n52938, C2 => 
                           n61910, A => n6872, ZN => n6871);
   U6155 : OAI221_X1 port map( B1 => n898, B2 => n6018, C1 => n874, C2 => 
                           n61734, A => n6873, ZN => n6870);
   U6156 : NOR4_X1 port map( A1 => n6793, A2 => n6794, A3 => n6795, A4 => n6796
                           , ZN => n6792);
   U6157 : OAI221_X1 port map( B1 => n2236, B2 => n6021, C1 => n2258, C2 => 
                           n61730, A => n6799, ZN => n6794);
   U6158 : OAI221_X1 port map( B1 => n61718, B2 => n1714, C1 => n52937, C2 => 
                           n61910, A => n6797, ZN => n6796);
   U6159 : OAI221_X1 port map( B1 => n897, B2 => n6018, C1 => n873, C2 => 
                           n61734, A => n6798, ZN => n6795);
   U6160 : NOR4_X1 port map( A1 => n7243, A2 => n7244, A3 => n7245, A4 => n7246
                           , ZN => n7242);
   U6161 : OAI221_X1 port map( B1 => n2241, B2 => n61727, C1 => n2263, C2 => 
                           n61729, A => n7249, ZN => n7244);
   U6162 : OAI221_X1 port map( B1 => n61717, B2 => n1720, C1 => n52943, C2 => 
                           n61909, A => n7247, ZN => n7246);
   U6163 : OAI221_X1 port map( B1 => n903, B2 => n61731, C1 => n879, C2 => 
                           n61733, A => n7248, ZN => n7245);
   U6164 : NOR4_X1 port map( A1 => n7843, A2 => n7844, A3 => n7845, A4 => n7846
                           , ZN => n7842);
   U6165 : OAI221_X1 port map( B1 => n2076, B2 => n61727, C1 => n2078, C2 => 
                           n61729, A => n7858, ZN => n7844);
   U6166 : OAI221_X1 port map( B1 => n61717, B2 => n1728, C1 => n52951, C2 => 
                           n61909, A => n7847, ZN => n7846);
   U6167 : OAI221_X1 port map( B1 => n911, B2 => n61731, C1 => n887, C2 => 
                           n61733, A => n7854, ZN => n7845);
   U6168 : NOR4_X1 port map( A1 => n7768, A2 => n7769, A3 => n7770, A4 => n7771
                           , ZN => n7767);
   U6169 : OAI221_X1 port map( B1 => n2248, B2 => n61727, C1 => n2270, C2 => 
                           n61729, A => n7774, ZN => n7769);
   U6170 : OAI221_X1 port map( B1 => n61717, B2 => n1727, C1 => n52950, C2 => 
                           n61909, A => n7772, ZN => n7771);
   U6171 : OAI221_X1 port map( B1 => n910, B2 => n61731, C1 => n886, C2 => 
                           n61733, A => n7773, ZN => n7770);
   U6172 : NOR4_X1 port map( A1 => n7693, A2 => n7694, A3 => n7695, A4 => n7696
                           , ZN => n7692);
   U6173 : OAI221_X1 port map( B1 => n2247, B2 => n61727, C1 => n2269, C2 => 
                           n61729, A => n7699, ZN => n7694);
   U6174 : OAI221_X1 port map( B1 => n61717, B2 => n1726, C1 => n52949, C2 => 
                           n61909, A => n7697, ZN => n7696);
   U6175 : OAI221_X1 port map( B1 => n909, B2 => n61731, C1 => n885, C2 => 
                           n61733, A => n7698, ZN => n7695);
   U6176 : NOR4_X1 port map( A1 => n7618, A2 => n7619, A3 => n7620, A4 => n7621
                           , ZN => n7617);
   U6177 : OAI221_X1 port map( B1 => n2246, B2 => n61727, C1 => n2268, C2 => 
                           n61729, A => n7624, ZN => n7619);
   U6178 : OAI221_X1 port map( B1 => n61717, B2 => n1725, C1 => n52948, C2 => 
                           n61909, A => n7622, ZN => n7621);
   U6179 : OAI221_X1 port map( B1 => n908, B2 => n61731, C1 => n884, C2 => 
                           n61733, A => n7623, ZN => n7620);
   U6180 : NOR4_X1 port map( A1 => n7543, A2 => n7544, A3 => n7545, A4 => n7546
                           , ZN => n7542);
   U6181 : OAI221_X1 port map( B1 => n2245, B2 => n61727, C1 => n2267, C2 => 
                           n61729, A => n7549, ZN => n7544);
   U6182 : OAI221_X1 port map( B1 => n61717, B2 => n1724, C1 => n52947, C2 => 
                           n61909, A => n7547, ZN => n7546);
   U6183 : OAI221_X1 port map( B1 => n907, B2 => n61731, C1 => n883, C2 => 
                           n61733, A => n7548, ZN => n7545);
   U6184 : NOR4_X1 port map( A1 => n7468, A2 => n7469, A3 => n7470, A4 => n7471
                           , ZN => n7467);
   U6185 : OAI221_X1 port map( B1 => n2244, B2 => n61727, C1 => n2266, C2 => 
                           n61729, A => n7474, ZN => n7469);
   U6186 : OAI221_X1 port map( B1 => n61717, B2 => n1723, C1 => n52946, C2 => 
                           n61909, A => n7472, ZN => n7471);
   U6187 : OAI221_X1 port map( B1 => n906, B2 => n61731, C1 => n882, C2 => 
                           n61733, A => n7473, ZN => n7470);
   U6188 : NOR4_X1 port map( A1 => n7393, A2 => n7394, A3 => n7395, A4 => n7396
                           , ZN => n7392);
   U6189 : OAI221_X1 port map( B1 => n2243, B2 => n61727, C1 => n2265, C2 => 
                           n61729, A => n7399, ZN => n7394);
   U6190 : OAI221_X1 port map( B1 => n61717, B2 => n1722, C1 => n52945, C2 => 
                           n61909, A => n7397, ZN => n7396);
   U6191 : OAI221_X1 port map( B1 => n905, B2 => n61731, C1 => n881, C2 => 
                           n61733, A => n7398, ZN => n7395);
   U6192 : NOR4_X1 port map( A1 => n7318, A2 => n7319, A3 => n7320, A4 => n7321
                           , ZN => n7317);
   U6193 : OAI221_X1 port map( B1 => n2242, B2 => n61727, C1 => n2264, C2 => 
                           n61729, A => n7324, ZN => n7319);
   U6194 : OAI221_X1 port map( B1 => n61717, B2 => n1721, C1 => n52944, C2 => 
                           n61909, A => n7322, ZN => n7321);
   U6195 : OAI221_X1 port map( B1 => n904, B2 => n61731, C1 => n880, C2 => 
                           n61733, A => n7323, ZN => n7320);
   U6196 : NOR4_X1 port map( A1 => n7168, A2 => n7169, A3 => n7170, A4 => n7171
                           , ZN => n7167);
   U6197 : OAI221_X1 port map( B1 => n2240, B2 => n61727, C1 => n2262, C2 => 
                           n61729, A => n7174, ZN => n7169);
   U6198 : OAI221_X1 port map( B1 => n61717, B2 => n1719, C1 => n52942, C2 => 
                           n61909, A => n7172, ZN => n7171);
   U6199 : OAI221_X1 port map( B1 => n902, B2 => n61731, C1 => n878, C2 => 
                           n61733, A => n7173, ZN => n7170);
   U6200 : NOR4_X1 port map( A1 => n6943, A2 => n6944, A3 => n6945, A4 => n6946
                           , ZN => n6942);
   U6201 : OAI221_X1 port map( B1 => n2238, B2 => n6021, C1 => n2260, C2 => 
                           n61730, A => n6949, ZN => n6944);
   U6202 : OAI221_X1 port map( B1 => n61718, B2 => n1716, C1 => n52939, C2 => 
                           n61910, A => n6947, ZN => n6946);
   U6203 : OAI221_X1 port map( B1 => n899, B2 => n6018, C1 => n875, C2 => 
                           n61734, A => n6948, ZN => n6945);
   U6204 : NOR4_X1 port map( A1 => n6012, A2 => n6013, A3 => n6014, A4 => n6015
                           , ZN => n6011);
   U6205 : OAI221_X1 port map( B1 => n5386, B2 => n1045, C1 => n5387, C2 => 
                           n3955, A => n6016, ZN => n6015);
   U6206 : OAI221_X1 port map( B1 => n61956, B2 => n4155, C1 => n61953, C2 => 
                           n4163, A => n6019, ZN => n6014);
   U6207 : OAI221_X1 port map( B1 => n51647, B2 => n61949, C1 => n51639, C2 => 
                           n61946, A => n6022, ZN => n6013);
   U6208 : NOR4_X1 port map( A1 => n5937, A2 => n5938, A3 => n5939, A4 => n5940
                           , ZN => n5936);
   U6209 : OAI221_X1 port map( B1 => n5386, B2 => n1044, C1 => n5387, C2 => 
                           n3954, A => n5941, ZN => n5940);
   U6210 : OAI221_X1 port map( B1 => n61956, B2 => n4154, C1 => n61953, C2 => 
                           n4162, A => n5942, ZN => n5939);
   U6211 : OAI221_X1 port map( B1 => n51646, B2 => n61950, C1 => n51638, C2 => 
                           n61946, A => n5943, ZN => n5938);
   U6212 : NOR4_X1 port map( A1 => n5787, A2 => n5788, A3 => n5789, A4 => n5790
                           , ZN => n5786);
   U6213 : OAI221_X1 port map( B1 => n5386, B2 => n1042, C1 => n5387, C2 => 
                           n3952, A => n5791, ZN => n5790);
   U6214 : OAI221_X1 port map( B1 => n61956, B2 => n4152, C1 => n61953, C2 => 
                           n4160, A => n5792, ZN => n5789);
   U6215 : OAI221_X1 port map( B1 => n51644, B2 => n61950, C1 => n51636, C2 => 
                           n61946, A => n5793, ZN => n5788);
   U6216 : NOR4_X1 port map( A1 => n5562, A2 => n5563, A3 => n5564, A4 => n5565
                           , ZN => n5561);
   U6217 : OAI221_X1 port map( B1 => n5386, B2 => n1039, C1 => n5387, C2 => 
                           n3949, A => n5566, ZN => n5565);
   U6218 : OAI221_X1 port map( B1 => n61956, B2 => n4149, C1 => n61953, C2 => 
                           n4157, A => n5567, ZN => n5564);
   U6219 : OAI221_X1 port map( B1 => n51641, B2 => n61950, C1 => n51633, C2 => 
                           n61946, A => n5568, ZN => n5563);
   U6220 : NOR4_X1 port map( A1 => n5382, A2 => n5383, A3 => n5384, A4 => n5385
                           , ZN => n5381);
   U6221 : OAI221_X1 port map( B1 => n5386, B2 => n1038, C1 => n5387, C2 => 
                           n3948, A => n5388, ZN => n5385);
   U6222 : OAI221_X1 port map( B1 => n61956, B2 => n4148, C1 => n61953, C2 => 
                           n4156, A => n5391, ZN => n5384);
   U6223 : OAI221_X1 port map( B1 => n51640, B2 => n61949, C1 => n51632, C2 => 
                           n61946, A => n5394, ZN => n5383);
   U6224 : NOR4_X1 port map( A1 => n14372, A2 => n14373, A3 => n14374, A4 => 
                           n14375, ZN => n14371);
   U6225 : OAI221_X1 port map( B1 => n4591, B2 => n61640, C1 => n4615, C2 => 
                           n61637, A => n14378, ZN => n14373);
   U6226 : OAI221_X1 port map( B1 => n4663, B2 => n61652, C1 => n4687, C2 => 
                           n61649, A => n14377, ZN => n14374);
   U6227 : OAI221_X1 port map( B1 => n2241, B2 => n61664, C1 => n2263, C2 => 
                           n61661, A => n14376, ZN => n14375);
   U6228 : NOR4_X1 port map( A1 => n9881, A2 => n9882, A3 => n9883, A4 => n9884
                           , ZN => n9880);
   U6229 : OAI221_X1 port map( B1 => n4590, B2 => n61640, C1 => n4614, C2 => 
                           n61637, A => n9887, ZN => n9882);
   U6230 : OAI221_X1 port map( B1 => n4662, B2 => n61652, C1 => n4686, C2 => 
                           n61649, A => n9886, ZN => n9883);
   U6231 : OAI221_X1 port map( B1 => n2240, B2 => n61664, C1 => n2262, C2 => 
                           n61661, A => n9885, ZN => n9884);
   U6232 : NOR4_X1 port map( A1 => n9742, A2 => n9743, A3 => n9744, A4 => n9745
                           , ZN => n9741);
   U6233 : OAI221_X1 port map( B1 => n4589, B2 => n61640, C1 => n4613, C2 => 
                           n61637, A => n9812, ZN => n9743);
   U6234 : OAI221_X1 port map( B1 => n4661, B2 => n61652, C1 => n4685, C2 => 
                           n61649, A => n9811, ZN => n9744);
   U6235 : OAI221_X1 port map( B1 => n2239, B2 => n61664, C1 => n2261, C2 => 
                           n61661, A => n9746, ZN => n9745);
   U6236 : NOR4_X1 port map( A1 => n9667, A2 => n9668, A3 => n9669, A4 => n9670
                           , ZN => n9666);
   U6237 : OAI221_X1 port map( B1 => n4588, B2 => n61640, C1 => n4612, C2 => 
                           n61637, A => n9673, ZN => n9668);
   U6238 : OAI221_X1 port map( B1 => n4660, B2 => n61652, C1 => n4684, C2 => 
                           n61649, A => n9672, ZN => n9669);
   U6239 : OAI221_X1 port map( B1 => n2075, B2 => n61664, C1 => n2077, C2 => 
                           n61661, A => n9671, ZN => n9670);
   U6240 : NOR4_X1 port map( A1 => n9576, A2 => n9577, A3 => n9578, A4 => n9579
                           , ZN => n9575);
   U6241 : OAI221_X1 port map( B1 => n4587, B2 => n61641, C1 => n4611, C2 => 
                           n61638, A => n9582, ZN => n9577);
   U6242 : OAI221_X1 port map( B1 => n4659, B2 => n61653, C1 => n4683, C2 => 
                           n61650, A => n9581, ZN => n9578);
   U6243 : OAI221_X1 port map( B1 => n2238, B2 => n61665, C1 => n2260, C2 => 
                           n61662, A => n9580, ZN => n9579);
   U6244 : NOR4_X1 port map( A1 => n9501, A2 => n9502, A3 => n9503, A4 => n9504
                           , ZN => n9500);
   U6245 : OAI221_X1 port map( B1 => n4586, B2 => n61641, C1 => n4610, C2 => 
                           n61638, A => n9507, ZN => n9502);
   U6246 : OAI221_X1 port map( B1 => n4658, B2 => n61653, C1 => n4682, C2 => 
                           n61650, A => n9506, ZN => n9503);
   U6247 : OAI221_X1 port map( B1 => n2237, B2 => n61665, C1 => n2259, C2 => 
                           n61662, A => n9505, ZN => n9504);
   U6248 : NOR4_X1 port map( A1 => n9426, A2 => n9427, A3 => n9428, A4 => n9429
                           , ZN => n9425);
   U6249 : OAI221_X1 port map( B1 => n4585, B2 => n61641, C1 => n4609, C2 => 
                           n61638, A => n9432, ZN => n9427);
   U6250 : OAI221_X1 port map( B1 => n4657, B2 => n61653, C1 => n4681, C2 => 
                           n61650, A => n9431, ZN => n9428);
   U6251 : OAI221_X1 port map( B1 => n2236, B2 => n61665, C1 => n2258, C2 => 
                           n61662, A => n9430, ZN => n9429);
   U6252 : NOR4_X1 port map( A1 => n9351, A2 => n9352, A3 => n9353, A4 => n9354
                           , ZN => n9350);
   U6253 : OAI221_X1 port map( B1 => n4584, B2 => n61641, C1 => n4608, C2 => 
                           n61638, A => n9357, ZN => n9352);
   U6254 : OAI221_X1 port map( B1 => n4656, B2 => n61653, C1 => n4680, C2 => 
                           n61650, A => n9356, ZN => n9353);
   U6255 : OAI221_X1 port map( B1 => n2235, B2 => n61665, C1 => n2257, C2 => 
                           n61662, A => n9355, ZN => n9354);
   U6256 : NOR4_X1 port map( A1 => n9212, A2 => n9213, A3 => n9214, A4 => n9215
                           , ZN => n9211);
   U6257 : OAI221_X1 port map( B1 => n4583, B2 => n61641, C1 => n4607, C2 => 
                           n61638, A => n9218, ZN => n9213);
   U6258 : OAI221_X1 port map( B1 => n4655, B2 => n61653, C1 => n4679, C2 => 
                           n61650, A => n9217, ZN => n9214);
   U6259 : OAI221_X1 port map( B1 => n2220, B2 => n61665, C1 => n2256, C2 => 
                           n61662, A => n9216, ZN => n9215);
   U6260 : NOR4_X1 port map( A1 => n9137, A2 => n9138, A3 => n9139, A4 => n9140
                           , ZN => n9136);
   U6261 : OAI221_X1 port map( B1 => n4582, B2 => n61641, C1 => n4606, C2 => 
                           n61638, A => n9143, ZN => n9138);
   U6262 : OAI221_X1 port map( B1 => n4654, B2 => n61653, C1 => n4678, C2 => 
                           n61650, A => n9142, ZN => n9139);
   U6263 : OAI221_X1 port map( B1 => n2219, B2 => n61665, C1 => n2255, C2 => 
                           n61662, A => n9141, ZN => n9140);
   U6264 : NOR4_X1 port map( A1 => n9062, A2 => n9063, A3 => n9064, A4 => n9065
                           , ZN => n9061);
   U6265 : OAI221_X1 port map( B1 => n4581, B2 => n61641, C1 => n4605, C2 => 
                           n61638, A => n9068, ZN => n9063);
   U6266 : OAI221_X1 port map( B1 => n4653, B2 => n61653, C1 => n4677, C2 => 
                           n61650, A => n9067, ZN => n9064);
   U6267 : OAI221_X1 port map( B1 => n2218, B2 => n61665, C1 => n2254, C2 => 
                           n61662, A => n9066, ZN => n9065);
   U6268 : NOR4_X1 port map( A1 => n8987, A2 => n8988, A3 => n8989, A4 => n8990
                           , ZN => n8986);
   U6269 : OAI221_X1 port map( B1 => n4580, B2 => n61641, C1 => n4604, C2 => 
                           n61638, A => n8993, ZN => n8988);
   U6270 : OAI221_X1 port map( B1 => n4652, B2 => n61653, C1 => n4676, C2 => 
                           n61650, A => n8992, ZN => n8989);
   U6271 : OAI221_X1 port map( B1 => n2217, B2 => n61665, C1 => n2253, C2 => 
                           n61662, A => n8991, ZN => n8990);
   U6272 : NOR4_X1 port map( A1 => n8912, A2 => n8913, A3 => n8914, A4 => n8915
                           , ZN => n8911);
   U6273 : OAI221_X1 port map( B1 => n4579, B2 => n61641, C1 => n4603, C2 => 
                           n61638, A => n8918, ZN => n8913);
   U6274 : OAI221_X1 port map( B1 => n4651, B2 => n61653, C1 => n4675, C2 => 
                           n61650, A => n8917, ZN => n8914);
   U6275 : OAI221_X1 port map( B1 => n2216, B2 => n61665, C1 => n2252, C2 => 
                           n61662, A => n8916, ZN => n8915);
   U6276 : NOR4_X1 port map( A1 => n8837, A2 => n8838, A3 => n8839, A4 => n8840
                           , ZN => n8836);
   U6277 : OAI221_X1 port map( B1 => n4578, B2 => n61641, C1 => n4602, C2 => 
                           n61638, A => n8843, ZN => n8838);
   U6278 : OAI221_X1 port map( B1 => n4650, B2 => n61653, C1 => n4674, C2 => 
                           n61650, A => n8842, ZN => n8839);
   U6279 : OAI221_X1 port map( B1 => n2215, B2 => n61665, C1 => n2251, C2 => 
                           n61662, A => n8841, ZN => n8840);
   U6280 : NOR4_X1 port map( A1 => n8762, A2 => n8763, A3 => n8764, A4 => n8765
                           , ZN => n8761);
   U6281 : OAI221_X1 port map( B1 => n4577, B2 => n61641, C1 => n4601, C2 => 
                           n61638, A => n8768, ZN => n8763);
   U6282 : OAI221_X1 port map( B1 => n4649, B2 => n61653, C1 => n4673, C2 => 
                           n61650, A => n8767, ZN => n8764);
   U6283 : OAI221_X1 port map( B1 => n2214, B2 => n61665, C1 => n2250, C2 => 
                           n61662, A => n8766, ZN => n8765);
   U6284 : NOR4_X1 port map( A1 => n8687, A2 => n8688, A3 => n8689, A4 => n8690
                           , ZN => n8686);
   U6285 : OAI221_X1 port map( B1 => n4576, B2 => n61641, C1 => n4600, C2 => 
                           n61638, A => n8693, ZN => n8688);
   U6286 : OAI221_X1 port map( B1 => n4648, B2 => n61653, C1 => n4672, C2 => 
                           n61650, A => n8692, ZN => n8689);
   U6287 : OAI221_X1 port map( B1 => n2213, B2 => n61665, C1 => n2249, C2 => 
                           n61662, A => n8691, ZN => n8690);
   U6288 : NOR4_X1 port map( A1 => n14972, A2 => n14973, A3 => n14974, A4 => 
                           n14975, ZN => n14971);
   U6289 : OAI221_X1 port map( B1 => n4599, B2 => n61640, C1 => n4623, C2 => 
                           n61637, A => n14989, ZN => n14973);
   U6290 : OAI221_X1 port map( B1 => n4671, B2 => n61652, C1 => n4695, C2 => 
                           n61649, A => n14982, ZN => n14974);
   U6291 : OAI221_X1 port map( B1 => n2076, B2 => n61664, C1 => n2078, C2 => 
                           n61661, A => n14976, ZN => n14975);
   U6292 : NOR4_X1 port map( A1 => n14897, A2 => n14898, A3 => n14899, A4 => 
                           n14900, ZN => n14896);
   U6293 : OAI221_X1 port map( B1 => n4598, B2 => n61640, C1 => n4622, C2 => 
                           n61637, A => n14903, ZN => n14898);
   U6294 : OAI221_X1 port map( B1 => n4670, B2 => n61652, C1 => n4694, C2 => 
                           n61649, A => n14902, ZN => n14899);
   U6295 : OAI221_X1 port map( B1 => n2248, B2 => n61664, C1 => n2270, C2 => 
                           n61661, A => n14901, ZN => n14900);
   U6296 : NOR4_X1 port map( A1 => n14822, A2 => n14823, A3 => n14824, A4 => 
                           n14825, ZN => n14821);
   U6297 : OAI221_X1 port map( B1 => n4597, B2 => n61640, C1 => n4621, C2 => 
                           n61637, A => n14828, ZN => n14823);
   U6298 : OAI221_X1 port map( B1 => n4669, B2 => n61652, C1 => n4693, C2 => 
                           n61649, A => n14827, ZN => n14824);
   U6299 : OAI221_X1 port map( B1 => n2247, B2 => n61664, C1 => n2269, C2 => 
                           n61661, A => n14826, ZN => n14825);
   U6300 : NOR4_X1 port map( A1 => n14747, A2 => n14748, A3 => n14749, A4 => 
                           n14750, ZN => n14746);
   U6301 : OAI221_X1 port map( B1 => n4596, B2 => n61640, C1 => n4620, C2 => 
                           n61637, A => n14753, ZN => n14748);
   U6302 : OAI221_X1 port map( B1 => n4668, B2 => n61652, C1 => n4692, C2 => 
                           n61649, A => n14752, ZN => n14749);
   U6303 : OAI221_X1 port map( B1 => n2246, B2 => n61664, C1 => n2268, C2 => 
                           n61661, A => n14751, ZN => n14750);
   U6304 : NOR4_X1 port map( A1 => n14672, A2 => n14673, A3 => n14674, A4 => 
                           n14675, ZN => n14671);
   U6305 : OAI221_X1 port map( B1 => n4595, B2 => n61640, C1 => n4619, C2 => 
                           n61637, A => n14678, ZN => n14673);
   U6306 : OAI221_X1 port map( B1 => n4667, B2 => n61652, C1 => n4691, C2 => 
                           n61649, A => n14677, ZN => n14674);
   U6307 : OAI221_X1 port map( B1 => n2245, B2 => n61664, C1 => n2267, C2 => 
                           n61661, A => n14676, ZN => n14675);
   U6308 : NOR4_X1 port map( A1 => n14597, A2 => n14598, A3 => n14599, A4 => 
                           n14600, ZN => n14596);
   U6309 : OAI221_X1 port map( B1 => n4594, B2 => n61640, C1 => n4618, C2 => 
                           n61637, A => n14603, ZN => n14598);
   U6310 : OAI221_X1 port map( B1 => n4666, B2 => n61652, C1 => n4690, C2 => 
                           n61649, A => n14602, ZN => n14599);
   U6311 : OAI221_X1 port map( B1 => n2244, B2 => n61664, C1 => n2266, C2 => 
                           n61661, A => n14601, ZN => n14600);
   U6312 : NOR4_X1 port map( A1 => n14522, A2 => n14523, A3 => n14524, A4 => 
                           n14525, ZN => n14521);
   U6313 : OAI221_X1 port map( B1 => n4593, B2 => n61640, C1 => n4617, C2 => 
                           n61637, A => n14528, ZN => n14523);
   U6314 : OAI221_X1 port map( B1 => n4665, B2 => n61652, C1 => n4689, C2 => 
                           n61649, A => n14527, ZN => n14524);
   U6315 : OAI221_X1 port map( B1 => n2243, B2 => n61664, C1 => n2265, C2 => 
                           n61661, A => n14526, ZN => n14525);
   U6316 : NOR4_X1 port map( A1 => n14447, A2 => n14448, A3 => n14449, A4 => 
                           n14450, ZN => n14446);
   U6317 : OAI221_X1 port map( B1 => n4592, B2 => n61640, C1 => n4616, C2 => 
                           n61637, A => n14453, ZN => n14448);
   U6318 : OAI221_X1 port map( B1 => n4664, B2 => n61652, C1 => n4688, C2 => 
                           n61649, A => n14452, ZN => n14449);
   U6319 : OAI221_X1 port map( B1 => n2242, B2 => n61664, C1 => n2264, C2 => 
                           n61661, A => n14451, ZN => n14450);
   U6320 : NOR4_X1 port map( A1 => n6067, A2 => n6068, A3 => n6069, A4 => n6070
                           , ZN => n6066);
   U6321 : OAI221_X1 port map( B1 => n61864, B2 => n388, C1 => n505, C2 => 
                           n61863, A => n6071, ZN => n6070);
   U6322 : OAI221_X1 port map( B1 => n61848, B2 => n4051, C1 => n61845, C2 => 
                           n4059, A => n6075, ZN => n6068);
   U6323 : OAI221_X1 port map( B1 => n5484, B2 => n276, C1 => n5485, C2 => n300
                           , A => n6076, ZN => n6067);
   U6324 : NOR4_X1 port map( A1 => n5862, A2 => n5863, A3 => n5864, A4 => n5865
                           , ZN => n5861);
   U6325 : OAI221_X1 port map( B1 => n5386, B2 => n1043, C1 => n5387, C2 => 
                           n3953, A => n5866, ZN => n5865);
   U6326 : OAI221_X1 port map( B1 => n61956, B2 => n4153, C1 => n61953, C2 => 
                           n4161, A => n5867, ZN => n5864);
   U6327 : OAI221_X1 port map( B1 => n51645, B2 => n61950, C1 => n51637, C2 => 
                           n61945, A => n5868, ZN => n5863);
   U6328 : NOR4_X1 port map( A1 => n5823, A2 => n5824, A3 => n5825, A4 => n5826
                           , ZN => n5822);
   U6329 : OAI221_X1 port map( B1 => n61864, B2 => n369, C1 => n502, C2 => 
                           n61863, A => n5827, ZN => n5826);
   U6330 : OAI221_X1 port map( B1 => n61848, B2 => n4048, C1 => n61845, C2 => 
                           n4056, A => n5829, ZN => n5824);
   U6331 : OAI221_X1 port map( B1 => n5484, B2 => n273, C1 => n5485, C2 => n297
                           , A => n5830, ZN => n5823);
   U6332 : NOR4_X1 port map( A1 => n5712, A2 => n5713, A3 => n5714, A4 => n5715
                           , ZN => n5711);
   U6333 : OAI221_X1 port map( B1 => n5386, B2 => n1041, C1 => n5387, C2 => 
                           n3951, A => n5716, ZN => n5715);
   U6334 : OAI221_X1 port map( B1 => n61956, B2 => n4151, C1 => n61953, C2 => 
                           n4159, A => n5717, ZN => n5714);
   U6335 : OAI221_X1 port map( B1 => n51643, B2 => n61950, C1 => n51635, C2 => 
                           n61945, A => n5718, ZN => n5713);
   U6336 : NOR4_X1 port map( A1 => n5637, A2 => n5638, A3 => n5639, A4 => n5640
                           , ZN => n5636);
   U6337 : OAI221_X1 port map( B1 => n5386, B2 => n1040, C1 => n5387, C2 => 
                           n3950, A => n5641, ZN => n5640);
   U6338 : OAI221_X1 port map( B1 => n61956, B2 => n4150, C1 => n61953, C2 => 
                           n4158, A => n5642, ZN => n5639);
   U6339 : OAI221_X1 port map( B1 => n51642, B2 => n61950, C1 => n51634, C2 => 
                           n61946, A => n5643, ZN => n5638);
   U6340 : NOR4_X1 port map( A1 => n5973, A2 => n5974, A3 => n5975, A4 => n5976
                           , ZN => n5972);
   U6341 : OAI221_X1 port map( B1 => n61864, B2 => n371, C1 => n504, C2 => 
                           n61863, A => n5977, ZN => n5976);
   U6342 : OAI221_X1 port map( B1 => n61848, B2 => n4050, C1 => n61845, C2 => 
                           n4058, A => n5979, ZN => n5974);
   U6343 : OAI221_X1 port map( B1 => n5484, B2 => n275, C1 => n5485, C2 => n299
                           , A => n5980, ZN => n5973);
   U6344 : NOR4_X1 port map( A1 => n5898, A2 => n5899, A3 => n5900, A4 => n5901
                           , ZN => n5897);
   U6345 : OAI221_X1 port map( B1 => n61864, B2 => n370, C1 => n503, C2 => 
                           n61863, A => n5902, ZN => n5901);
   U6346 : OAI221_X1 port map( B1 => n61848, B2 => n4049, C1 => n61845, C2 => 
                           n4057, A => n5904, ZN => n5899);
   U6347 : OAI221_X1 port map( B1 => n5484, B2 => n274, C1 => n5485, C2 => n298
                           , A => n5905, ZN => n5898);
   U6348 : NOR4_X1 port map( A1 => n5748, A2 => n5749, A3 => n5750, A4 => n5751
                           , ZN => n5747);
   U6349 : OAI221_X1 port map( B1 => n61864, B2 => n368, C1 => n501, C2 => 
                           n61863, A => n5752, ZN => n5751);
   U6350 : OAI221_X1 port map( B1 => n61848, B2 => n4047, C1 => n61845, C2 => 
                           n4055, A => n5754, ZN => n5749);
   U6351 : OAI221_X1 port map( B1 => n5484, B2 => n272, C1 => n5485, C2 => n296
                           , A => n5755, ZN => n5748);
   U6352 : NOR4_X1 port map( A1 => n5673, A2 => n5674, A3 => n5675, A4 => n5676
                           , ZN => n5672);
   U6353 : OAI221_X1 port map( B1 => n61864, B2 => n367, C1 => n500, C2 => 
                           n61863, A => n5677, ZN => n5676);
   U6354 : OAI221_X1 port map( B1 => n61848, B2 => n4046, C1 => n61845, C2 => 
                           n4054, A => n5679, ZN => n5674);
   U6355 : OAI221_X1 port map( B1 => n5484, B2 => n271, C1 => n5485, C2 => n295
                           , A => n5680, ZN => n5673);
   U6356 : NOR4_X1 port map( A1 => n5598, A2 => n5599, A3 => n5600, A4 => n5601
                           , ZN => n5597);
   U6357 : OAI221_X1 port map( B1 => n61864, B2 => n366, C1 => n475, C2 => 
                           n61863, A => n5602, ZN => n5601);
   U6358 : OAI221_X1 port map( B1 => n61848, B2 => n4045, C1 => n61845, C2 => 
                           n4053, A => n5604, ZN => n5599);
   U6359 : OAI221_X1 port map( B1 => n5484, B2 => n270, C1 => n5485, C2 => n294
                           , A => n5605, ZN => n5598);
   U6360 : NOR4_X1 port map( A1 => n5467, A2 => n5468, A3 => n5469, A4 => n5470
                           , ZN => n5466);
   U6361 : OAI221_X1 port map( B1 => n61864, B2 => n365, C1 => n474, C2 => 
                           n61863, A => n5473, ZN => n5470);
   U6362 : OAI221_X1 port map( B1 => n61848, B2 => n4044, C1 => n61845, C2 => 
                           n4052, A => n5481, ZN => n5468);
   U6363 : OAI221_X1 port map( B1 => n5484, B2 => n269, C1 => n5485, C2 => n293
                           , A => n5486, ZN => n5467);
   U6364 : NOR4_X1 port map( A1 => n6762, A2 => n6763, A3 => n6764, A4 => n6765
                           , ZN => n6752);
   U6365 : OAI221_X1 port map( B1 => n6078, B2 => n2154, C1 => n61692, C2 => 
                           n2082, A => n6766, ZN => n6765);
   U6366 : OAI221_X1 port map( B1 => n61826, B2 => n2030, C1 => n61823, C2 => 
                           n1982, A => n6768, ZN => n6763);
   U6367 : OAI221_X1 port map( B1 => n173, B2 => n6086, C1 => n197, C2 => 
                           n61688, A => n6767, ZN => n6764);
   U6368 : NOR4_X1 port map( A1 => n6687, A2 => n6688, A3 => n6689, A4 => n6690
                           , ZN => n6677);
   U6369 : OAI221_X1 port map( B1 => n6078, B2 => n2153, C1 => n61692, C2 => 
                           n2081, A => n6691, ZN => n6690);
   U6370 : OAI221_X1 port map( B1 => n61826, B2 => n2029, C1 => n61823, C2 => 
                           n1981, A => n6693, ZN => n6688);
   U6371 : OAI221_X1 port map( B1 => n172, B2 => n6086, C1 => n196, C2 => 
                           n61688, A => n6692, ZN => n6689);
   U6372 : NOR4_X1 port map( A1 => n6612, A2 => n6613, A3 => n6614, A4 => n6615
                           , ZN => n6602);
   U6373 : OAI221_X1 port map( B1 => n6078, B2 => n2152, C1 => n61692, C2 => 
                           n2080, A => n6616, ZN => n6615);
   U6374 : OAI221_X1 port map( B1 => n61826, B2 => n2028, C1 => n61823, C2 => 
                           n1980, A => n6618, ZN => n6613);
   U6375 : OAI221_X1 port map( B1 => n171, B2 => n6086, C1 => n195, C2 => 
                           n61688, A => n6617, ZN => n6614);
   U6376 : NOR4_X1 port map( A1 => n6537, A2 => n6538, A3 => n6539, A4 => n6540
                           , ZN => n6527);
   U6377 : OAI221_X1 port map( B1 => n6078, B2 => n2151, C1 => n61692, C2 => 
                           n2079, A => n6541, ZN => n6540);
   U6378 : OAI221_X1 port map( B1 => n61826, B2 => n2027, C1 => n61823, C2 => 
                           n1979, A => n6543, ZN => n6538);
   U6379 : OAI221_X1 port map( B1 => n170, B2 => n6086, C1 => n194, C2 => 
                           n61688, A => n6542, ZN => n6539);
   U6380 : NOR4_X1 port map( A1 => n6462, A2 => n6463, A3 => n6464, A4 => n6465
                           , ZN => n6452);
   U6381 : OAI221_X1 port map( B1 => n6078, B2 => n2150, C1 => n61692, C2 => 
                           n2074, A => n6466, ZN => n6465);
   U6382 : OAI221_X1 port map( B1 => n61826, B2 => n2026, C1 => n61823, C2 => 
                           n1978, A => n6468, ZN => n6463);
   U6383 : OAI221_X1 port map( B1 => n169, B2 => n6086, C1 => n193, C2 => 
                           n61688, A => n6467, ZN => n6464);
   U6384 : NOR4_X1 port map( A1 => n6387, A2 => n6388, A3 => n6389, A4 => n6390
                           , ZN => n6377);
   U6385 : OAI221_X1 port map( B1 => n6078, B2 => n2149, C1 => n61692, C2 => 
                           n2073, A => n6391, ZN => n6390);
   U6386 : OAI221_X1 port map( B1 => n61826, B2 => n2025, C1 => n61823, C2 => 
                           n1977, A => n6393, ZN => n6388);
   U6387 : OAI221_X1 port map( B1 => n168, B2 => n6086, C1 => n192, C2 => 
                           n61688, A => n6392, ZN => n6389);
   U6388 : NOR4_X1 port map( A1 => n6312, A2 => n6313, A3 => n6314, A4 => n6315
                           , ZN => n6302);
   U6389 : OAI221_X1 port map( B1 => n6078, B2 => n2148, C1 => n61692, C2 => 
                           n2072, A => n6316, ZN => n6315);
   U6390 : OAI221_X1 port map( B1 => n61826, B2 => n2024, C1 => n61823, C2 => 
                           n1976, A => n6318, ZN => n6313);
   U6391 : OAI221_X1 port map( B1 => n167, B2 => n6086, C1 => n191, C2 => 
                           n61688, A => n6317, ZN => n6314);
   U6392 : NOR4_X1 port map( A1 => n6237, A2 => n6238, A3 => n6239, A4 => n6240
                           , ZN => n6227);
   U6393 : OAI221_X1 port map( B1 => n6078, B2 => n2147, C1 => n61692, C2 => 
                           n2071, A => n6241, ZN => n6240);
   U6394 : OAI221_X1 port map( B1 => n61826, B2 => n2023, C1 => n61823, C2 => 
                           n1975, A => n6243, ZN => n6238);
   U6395 : OAI221_X1 port map( B1 => n166, B2 => n6086, C1 => n190, C2 => 
                           n61688, A => n6242, ZN => n6239);
   U6396 : NOR4_X1 port map( A1 => n6162, A2 => n6163, A3 => n6164, A4 => n6165
                           , ZN => n6152);
   U6397 : OAI221_X1 port map( B1 => n6078, B2 => n2146, C1 => n61692, C2 => 
                           n2070, A => n6166, ZN => n6165);
   U6398 : OAI221_X1 port map( B1 => n61826, B2 => n1998, C1 => n61823, C2 => 
                           n1974, A => n6168, ZN => n6163);
   U6399 : OAI221_X1 port map( B1 => n165, B2 => n6086, C1 => n189, C2 => 
                           n61688, A => n6167, ZN => n6164);
   U6400 : NOR4_X1 port map( A1 => n7137, A2 => n7138, A3 => n7139, A4 => n7140
                           , ZN => n7127);
   U6401 : OAI221_X1 port map( B1 => n61689, B2 => n2159, C1 => n61691, C2 => 
                           n2087, A => n7141, ZN => n7140);
   U6402 : OAI221_X1 port map( B1 => n61825, B2 => n2035, C1 => n61822, C2 => 
                           n1987, A => n7143, ZN => n7138);
   U6403 : OAI221_X1 port map( B1 => n178, B2 => n61685, C1 => n202, C2 => 
                           n61687, A => n7142, ZN => n7139);
   U6404 : NOR4_X1 port map( A1 => n7062, A2 => n7063, A3 => n7064, A4 => n7065
                           , ZN => n7052);
   U6405 : OAI221_X1 port map( B1 => n61689, B2 => n2158, C1 => n61691, C2 => 
                           n2086, A => n7066, ZN => n7065);
   U6406 : OAI221_X1 port map( B1 => n61825, B2 => n2034, C1 => n61822, C2 => 
                           n1986, A => n7068, ZN => n7063);
   U6407 : OAI221_X1 port map( B1 => n177, B2 => n61685, C1 => n201, C2 => 
                           n61687, A => n7067, ZN => n7064);
   U6408 : NOR4_X1 port map( A1 => n6912, A2 => n6913, A3 => n6914, A4 => n6915
                           , ZN => n6902);
   U6409 : OAI221_X1 port map( B1 => n6078, B2 => n2156, C1 => n61692, C2 => 
                           n2084, A => n6916, ZN => n6915);
   U6410 : OAI221_X1 port map( B1 => n61826, B2 => n2032, C1 => n61823, C2 => 
                           n1984, A => n6918, ZN => n6913);
   U6411 : OAI221_X1 port map( B1 => n175, B2 => n6086, C1 => n199, C2 => 
                           n61688, A => n6917, ZN => n6914);
   U6412 : NOR4_X1 port map( A1 => n6837, A2 => n6838, A3 => n6839, A4 => n6840
                           , ZN => n6827);
   U6413 : OAI221_X1 port map( B1 => n6078, B2 => n2155, C1 => n61692, C2 => 
                           n2083, A => n6841, ZN => n6840);
   U6414 : OAI221_X1 port map( B1 => n61826, B2 => n2031, C1 => n61823, C2 => 
                           n1983, A => n6843, ZN => n6838);
   U6415 : OAI221_X1 port map( B1 => n174, B2 => n6086, C1 => n198, C2 => 
                           n61688, A => n6842, ZN => n6839);
   U6416 : NOR4_X1 port map( A1 => n7287, A2 => n7288, A3 => n7289, A4 => n7290
                           , ZN => n7277);
   U6417 : OAI221_X1 port map( B1 => n61689, B2 => n2161, C1 => n61691, C2 => 
                           n2089, A => n7291, ZN => n7290);
   U6418 : OAI221_X1 port map( B1 => n61825, B2 => n2037, C1 => n61822, C2 => 
                           n1989, A => n7293, ZN => n7288);
   U6419 : OAI221_X1 port map( B1 => n180, B2 => n61685, C1 => n204, C2 => 
                           n61687, A => n7292, ZN => n7289);
   U6420 : NOR4_X1 port map( A1 => n7915, A2 => n7916, A3 => n7917, A4 => n7918
                           , ZN => n7902);
   U6421 : OAI221_X1 port map( B1 => n61689, B2 => n2169, C1 => n61691, C2 => 
                           n2097, A => n7919, ZN => n7918);
   U6422 : OAI221_X1 port map( B1 => n61825, B2 => n2045, C1 => n61822, C2 => 
                           n1997, A => n7922, ZN => n7916);
   U6423 : OAI221_X1 port map( B1 => n188, B2 => n61685, C1 => n212, C2 => 
                           n61687, A => n7921, ZN => n7917);
   U6424 : NOR4_X1 port map( A1 => n7812, A2 => n7813, A3 => n7814, A4 => n7815
                           , ZN => n7802);
   U6425 : OAI221_X1 port map( B1 => n61689, B2 => n2168, C1 => n61691, C2 => 
                           n2096, A => n7816, ZN => n7815);
   U6426 : OAI221_X1 port map( B1 => n61825, B2 => n2044, C1 => n61822, C2 => 
                           n1996, A => n7818, ZN => n7813);
   U6427 : OAI221_X1 port map( B1 => n187, B2 => n61685, C1 => n211, C2 => 
                           n61687, A => n7817, ZN => n7814);
   U6428 : NOR4_X1 port map( A1 => n7737, A2 => n7738, A3 => n7739, A4 => n7740
                           , ZN => n7727);
   U6429 : OAI221_X1 port map( B1 => n61689, B2 => n2167, C1 => n61691, C2 => 
                           n2095, A => n7741, ZN => n7740);
   U6430 : OAI221_X1 port map( B1 => n61825, B2 => n2043, C1 => n61822, C2 => 
                           n1995, A => n7743, ZN => n7738);
   U6431 : OAI221_X1 port map( B1 => n186, B2 => n61685, C1 => n210, C2 => 
                           n61687, A => n7742, ZN => n7739);
   U6432 : NOR4_X1 port map( A1 => n7662, A2 => n7663, A3 => n7664, A4 => n7665
                           , ZN => n7652);
   U6433 : OAI221_X1 port map( B1 => n61689, B2 => n2166, C1 => n61691, C2 => 
                           n2094, A => n7666, ZN => n7665);
   U6434 : OAI221_X1 port map( B1 => n61825, B2 => n2042, C1 => n61822, C2 => 
                           n1994, A => n7668, ZN => n7663);
   U6435 : OAI221_X1 port map( B1 => n185, B2 => n61685, C1 => n209, C2 => 
                           n61687, A => n7667, ZN => n7664);
   U6436 : NOR4_X1 port map( A1 => n7587, A2 => n7588, A3 => n7589, A4 => n7590
                           , ZN => n7577);
   U6437 : OAI221_X1 port map( B1 => n61689, B2 => n2165, C1 => n61691, C2 => 
                           n2093, A => n7591, ZN => n7590);
   U6438 : OAI221_X1 port map( B1 => n61825, B2 => n2041, C1 => n61822, C2 => 
                           n1993, A => n7593, ZN => n7588);
   U6439 : OAI221_X1 port map( B1 => n184, B2 => n61685, C1 => n208, C2 => 
                           n61687, A => n7592, ZN => n7589);
   U6440 : NOR4_X1 port map( A1 => n7512, A2 => n7513, A3 => n7514, A4 => n7515
                           , ZN => n7502);
   U6441 : OAI221_X1 port map( B1 => n61689, B2 => n2164, C1 => n61691, C2 => 
                           n2092, A => n7516, ZN => n7515);
   U6442 : OAI221_X1 port map( B1 => n61825, B2 => n2040, C1 => n61822, C2 => 
                           n1992, A => n7518, ZN => n7513);
   U6443 : OAI221_X1 port map( B1 => n183, B2 => n61685, C1 => n207, C2 => 
                           n61687, A => n7517, ZN => n7514);
   U6444 : NOR4_X1 port map( A1 => n7437, A2 => n7438, A3 => n7439, A4 => n7440
                           , ZN => n7427);
   U6445 : OAI221_X1 port map( B1 => n61689, B2 => n2163, C1 => n61691, C2 => 
                           n2091, A => n7441, ZN => n7440);
   U6446 : OAI221_X1 port map( B1 => n61825, B2 => n2039, C1 => n61822, C2 => 
                           n1991, A => n7443, ZN => n7438);
   U6447 : OAI221_X1 port map( B1 => n182, B2 => n61685, C1 => n206, C2 => 
                           n61687, A => n7442, ZN => n7439);
   U6448 : NOR4_X1 port map( A1 => n7362, A2 => n7363, A3 => n7364, A4 => n7365
                           , ZN => n7352);
   U6449 : OAI221_X1 port map( B1 => n61689, B2 => n2162, C1 => n61691, C2 => 
                           n2090, A => n7366, ZN => n7365);
   U6450 : OAI221_X1 port map( B1 => n61825, B2 => n2038, C1 => n61822, C2 => 
                           n1990, A => n7368, ZN => n7363);
   U6451 : OAI221_X1 port map( B1 => n181, B2 => n61685, C1 => n205, C2 => 
                           n61687, A => n7367, ZN => n7364);
   U6452 : NOR4_X1 port map( A1 => n7212, A2 => n7213, A3 => n7214, A4 => n7215
                           , ZN => n7202);
   U6453 : OAI221_X1 port map( B1 => n61689, B2 => n2160, C1 => n61691, C2 => 
                           n2088, A => n7216, ZN => n7215);
   U6454 : OAI221_X1 port map( B1 => n61825, B2 => n2036, C1 => n61822, C2 => 
                           n1988, A => n7218, ZN => n7213);
   U6455 : OAI221_X1 port map( B1 => n179, B2 => n61685, C1 => n203, C2 => 
                           n61687, A => n7217, ZN => n7214);
   U6456 : NOR4_X1 port map( A1 => n6987, A2 => n6988, A3 => n6989, A4 => n6990
                           , ZN => n6977);
   U6457 : OAI221_X1 port map( B1 => n6078, B2 => n2157, C1 => n61692, C2 => 
                           n2085, A => n6991, ZN => n6990);
   U6458 : OAI221_X1 port map( B1 => n61826, B2 => n2033, C1 => n61823, C2 => 
                           n1985, A => n6993, ZN => n6988);
   U6459 : OAI221_X1 port map( B1 => n176, B2 => n6086, C1 => n200, C2 => 
                           n61688, A => n6992, ZN => n6989);
   U6460 : NOR4_X1 port map( A1 => n6726, A2 => n6727, A3 => n6728, A4 => n6729
                           , ZN => n6716);
   U6461 : OAI221_X1 port map( B1 => n53156, B2 => n61922, C1 => n53180, C2 => 
                           n61918, A => n6732, ZN => n6727);
   U6462 : OAI221_X1 port map( B1 => n3417, B2 => n61934, C1 => n3441, C2 => 
                           n61931, A => n6731, ZN => n6728);
   U6463 : OAI221_X1 port map( B1 => n52964, B2 => n6034, C1 => n52988, C2 => 
                           n6033, A => n6733, ZN => n6726);
   U6464 : NOR4_X1 port map( A1 => n6651, A2 => n6652, A3 => n6653, A4 => n6654
                           , ZN => n6641);
   U6465 : OAI221_X1 port map( B1 => n53155, B2 => n61922, C1 => n53179, C2 => 
                           n61918, A => n6657, ZN => n6652);
   U6466 : OAI221_X1 port map( B1 => n3416, B2 => n61934, C1 => n3440, C2 => 
                           n61931, A => n6656, ZN => n6653);
   U6467 : OAI221_X1 port map( B1 => n52963, B2 => n6034, C1 => n52987, C2 => 
                           n6033, A => n6658, ZN => n6651);
   U6468 : NOR4_X1 port map( A1 => n6576, A2 => n6577, A3 => n6578, A4 => n6579
                           , ZN => n6566);
   U6469 : OAI221_X1 port map( B1 => n53154, B2 => n61922, C1 => n53178, C2 => 
                           n61918, A => n6582, ZN => n6577);
   U6470 : OAI221_X1 port map( B1 => n3415, B2 => n61934, C1 => n3439, C2 => 
                           n61931, A => n6581, ZN => n6578);
   U6471 : OAI221_X1 port map( B1 => n52962, B2 => n6034, C1 => n52986, C2 => 
                           n6033, A => n6583, ZN => n6576);
   U6472 : NOR4_X1 port map( A1 => n6501, A2 => n6502, A3 => n6503, A4 => n6504
                           , ZN => n6491);
   U6473 : OAI221_X1 port map( B1 => n53153, B2 => n61922, C1 => n53177, C2 => 
                           n61918, A => n6507, ZN => n6502);
   U6474 : OAI221_X1 port map( B1 => n3414, B2 => n61934, C1 => n3438, C2 => 
                           n61931, A => n6506, ZN => n6503);
   U6475 : OAI221_X1 port map( B1 => n52961, B2 => n6034, C1 => n52985, C2 => 
                           n6033, A => n6508, ZN => n6501);
   U6476 : NOR4_X1 port map( A1 => n6426, A2 => n6427, A3 => n6428, A4 => n6429
                           , ZN => n6416);
   U6477 : OAI221_X1 port map( B1 => n53152, B2 => n61922, C1 => n53176, C2 => 
                           n61919, A => n6432, ZN => n6427);
   U6478 : OAI221_X1 port map( B1 => n3413, B2 => n61934, C1 => n3437, C2 => 
                           n61931, A => n6431, ZN => n6428);
   U6479 : OAI221_X1 port map( B1 => n52960, B2 => n6034, C1 => n52984, C2 => 
                           n6033, A => n6433, ZN => n6426);
   U6480 : NOR4_X1 port map( A1 => n6351, A2 => n6352, A3 => n6353, A4 => n6354
                           , ZN => n6341);
   U6481 : OAI221_X1 port map( B1 => n53151, B2 => n61921, C1 => n53175, C2 => 
                           n61919, A => n6357, ZN => n6352);
   U6482 : OAI221_X1 port map( B1 => n3412, B2 => n61934, C1 => n3436, C2 => 
                           n61931, A => n6356, ZN => n6353);
   U6483 : OAI221_X1 port map( B1 => n52959, B2 => n6034, C1 => n52983, C2 => 
                           n6033, A => n6358, ZN => n6351);
   U6484 : NOR4_X1 port map( A1 => n6276, A2 => n6277, A3 => n6278, A4 => n6279
                           , ZN => n6266);
   U6485 : OAI221_X1 port map( B1 => n53150, B2 => n61921, C1 => n53174, C2 => 
                           n61918, A => n6282, ZN => n6277);
   U6486 : OAI221_X1 port map( B1 => n3411, B2 => n61934, C1 => n3435, C2 => 
                           n61931, A => n6281, ZN => n6278);
   U6487 : OAI221_X1 port map( B1 => n52958, B2 => n6034, C1 => n52982, C2 => 
                           n6033, A => n6283, ZN => n6276);
   U6488 : NOR4_X1 port map( A1 => n6201, A2 => n6202, A3 => n6203, A4 => n6204
                           , ZN => n6191);
   U6489 : OAI221_X1 port map( B1 => n53149, B2 => n61921, C1 => n53173, C2 => 
                           n61918, A => n6207, ZN => n6202);
   U6490 : OAI221_X1 port map( B1 => n3410, B2 => n61934, C1 => n3434, C2 => 
                           n61931, A => n6206, ZN => n6203);
   U6491 : OAI221_X1 port map( B1 => n52957, B2 => n6034, C1 => n52981, C2 => 
                           n6033, A => n6208, ZN => n6201);
   U6492 : NOR4_X1 port map( A1 => n6126, A2 => n6127, A3 => n6128, A4 => n6129
                           , ZN => n6116);
   U6493 : OAI221_X1 port map( B1 => n53148, B2 => n61921, C1 => n53172, C2 => 
                           n61918, A => n6132, ZN => n6127);
   U6494 : OAI221_X1 port map( B1 => n3409, B2 => n61934, C1 => n3433, C2 => 
                           n61931, A => n6131, ZN => n6128);
   U6495 : OAI221_X1 port map( B1 => n52956, B2 => n6034, C1 => n52980, C2 => 
                           n6033, A => n6133, ZN => n6126);
   U6496 : NOR4_X1 port map( A1 => n7101, A2 => n7102, A3 => n7103, A4 => n7104
                           , ZN => n7091);
   U6497 : OAI221_X1 port map( B1 => n53161, B2 => n61922, C1 => n53185, C2 => 
                           n61918, A => n7107, ZN => n7102);
   U6498 : OAI221_X1 port map( B1 => n3422, B2 => n61933, C1 => n3446, C2 => 
                           n61930, A => n7106, ZN => n7103);
   U6499 : OAI221_X1 port map( B1 => n52969, B2 => n61719, C1 => n52993, C2 => 
                           n61721, A => n1525, ZN => n7101);
   U6500 : NOR4_X1 port map( A1 => n7026, A2 => n7027, A3 => n7028, A4 => n7029
                           , ZN => n7016);
   U6501 : OAI221_X1 port map( B1 => n53160, B2 => n61922, C1 => n53184, C2 => 
                           n61918, A => n7032, ZN => n7027);
   U6502 : OAI221_X1 port map( B1 => n3421, B2 => n61933, C1 => n3445, C2 => 
                           n61930, A => n7031, ZN => n7028);
   U6503 : OAI221_X1 port map( B1 => n52968, B2 => n61719, C1 => n52992, C2 => 
                           n61721, A => n1523, ZN => n7026);
   U6504 : NOR4_X1 port map( A1 => n6876, A2 => n6877, A3 => n6878, A4 => n6879
                           , ZN => n6866);
   U6505 : OAI221_X1 port map( B1 => n53158, B2 => n61922, C1 => n53182, C2 => 
                           n61918, A => n6882, ZN => n6877);
   U6506 : OAI221_X1 port map( B1 => n3419, B2 => n61934, C1 => n3443, C2 => 
                           n61931, A => n6881, ZN => n6878);
   U6507 : OAI221_X1 port map( B1 => n52966, B2 => n6034, C1 => n52990, C2 => 
                           n6033, A => n1519, ZN => n6876);
   U6508 : NOR4_X1 port map( A1 => n6801, A2 => n6802, A3 => n6803, A4 => n6804
                           , ZN => n6791);
   U6509 : OAI221_X1 port map( B1 => n53157, B2 => n61922, C1 => n53181, C2 => 
                           n61918, A => n6807, ZN => n6802);
   U6510 : OAI221_X1 port map( B1 => n3418, B2 => n61934, C1 => n3442, C2 => 
                           n61931, A => n6806, ZN => n6803);
   U6511 : OAI221_X1 port map( B1 => n52965, B2 => n6034, C1 => n52989, C2 => 
                           n6033, A => n6808, ZN => n6801);
   U6512 : NOR4_X1 port map( A1 => n7251, A2 => n7252, A3 => n7253, A4 => n7254
                           , ZN => n7241);
   U6513 : OAI221_X1 port map( B1 => n53163, B2 => n61922, C1 => n61919, C2 => 
                           n3152, A => n7257, ZN => n7252);
   U6514 : OAI221_X1 port map( B1 => n3424, B2 => n61933, C1 => n3448, C2 => 
                           n61930, A => n7256, ZN => n7253);
   U6515 : OAI221_X1 port map( B1 => n52971, B2 => n61719, C1 => n52995, C2 => 
                           n61721, A => n1529, ZN => n7251);
   U6516 : NOR4_X1 port map( A1 => n7865, A2 => n7866, A3 => n7867, A4 => n7868
                           , ZN => n7841);
   U6517 : OAI221_X1 port map( B1 => n53171, B2 => n61923, C1 => n61919, C2 => 
                           n3160, A => n7874, ZN => n7866);
   U6518 : OAI221_X1 port map( B1 => n3432, B2 => n61933, C1 => n3456, C2 => 
                           n61930, A => n7871, ZN => n7867);
   U6519 : OAI221_X1 port map( B1 => n52979, B2 => n61719, C1 => n53003, C2 => 
                           n61721, A => n1545, ZN => n7865);
   U6520 : NOR4_X1 port map( A1 => n7776, A2 => n7777, A3 => n7778, A4 => n7779
                           , ZN => n7766);
   U6521 : OAI221_X1 port map( B1 => n53170, B2 => n61923, C1 => n61920, C2 => 
                           n3159, A => n7782, ZN => n7777);
   U6522 : OAI221_X1 port map( B1 => n3431, B2 => n61933, C1 => n3455, C2 => 
                           n61930, A => n7781, ZN => n7778);
   U6523 : OAI221_X1 port map( B1 => n52978, B2 => n61719, C1 => n53002, C2 => 
                           n61721, A => n1543, ZN => n7776);
   U6524 : NOR4_X1 port map( A1 => n7701, A2 => n7702, A3 => n7703, A4 => n7704
                           , ZN => n7691);
   U6525 : OAI221_X1 port map( B1 => n53169, B2 => n61923, C1 => n61920, C2 => 
                           n3158, A => n7707, ZN => n7702);
   U6526 : OAI221_X1 port map( B1 => n3430, B2 => n61933, C1 => n3454, C2 => 
                           n61930, A => n7706, ZN => n7703);
   U6527 : OAI221_X1 port map( B1 => n52977, B2 => n61719, C1 => n53001, C2 => 
                           n61721, A => n1541, ZN => n7701);
   U6528 : NOR4_X1 port map( A1 => n7626, A2 => n7627, A3 => n7628, A4 => n7629
                           , ZN => n7616);
   U6529 : OAI221_X1 port map( B1 => n53168, B2 => n61923, C1 => n61920, C2 => 
                           n3157, A => n7632, ZN => n7627);
   U6530 : OAI221_X1 port map( B1 => n3429, B2 => n61933, C1 => n3453, C2 => 
                           n61930, A => n7631, ZN => n7628);
   U6531 : OAI221_X1 port map( B1 => n52976, B2 => n61719, C1 => n53000, C2 => 
                           n61721, A => n1539, ZN => n7626);
   U6532 : NOR4_X1 port map( A1 => n7551, A2 => n7552, A3 => n7553, A4 => n7554
                           , ZN => n7541);
   U6533 : OAI221_X1 port map( B1 => n53167, B2 => n61923, C1 => n61920, C2 => 
                           n3156, A => n7557, ZN => n7552);
   U6534 : OAI221_X1 port map( B1 => n3428, B2 => n61933, C1 => n3452, C2 => 
                           n61930, A => n7556, ZN => n7553);
   U6535 : OAI221_X1 port map( B1 => n52975, B2 => n61719, C1 => n52999, C2 => 
                           n61721, A => n1537, ZN => n7551);
   U6536 : NOR4_X1 port map( A1 => n7476, A2 => n7477, A3 => n7478, A4 => n7479
                           , ZN => n7466);
   U6537 : OAI221_X1 port map( B1 => n53166, B2 => n61923, C1 => n61920, C2 => 
                           n3155, A => n7482, ZN => n7477);
   U6538 : OAI221_X1 port map( B1 => n3427, B2 => n61933, C1 => n3451, C2 => 
                           n61930, A => n7481, ZN => n7478);
   U6539 : OAI221_X1 port map( B1 => n52974, B2 => n61719, C1 => n52998, C2 => 
                           n61721, A => n1535, ZN => n7476);
   U6540 : NOR4_X1 port map( A1 => n7401, A2 => n7402, A3 => n7403, A4 => n7404
                           , ZN => n7391);
   U6541 : OAI221_X1 port map( B1 => n53165, B2 => n61923, C1 => n61920, C2 => 
                           n3154, A => n7407, ZN => n7402);
   U6542 : OAI221_X1 port map( B1 => n3426, B2 => n61933, C1 => n3450, C2 => 
                           n61930, A => n7406, ZN => n7403);
   U6543 : OAI221_X1 port map( B1 => n52973, B2 => n61719, C1 => n52997, C2 => 
                           n61721, A => n1533, ZN => n7401);
   U6544 : NOR4_X1 port map( A1 => n7326, A2 => n7327, A3 => n7328, A4 => n7329
                           , ZN => n7316);
   U6545 : OAI221_X1 port map( B1 => n53164, B2 => n61922, C1 => n61920, C2 => 
                           n3153, A => n7332, ZN => n7327);
   U6546 : OAI221_X1 port map( B1 => n3425, B2 => n61933, C1 => n3449, C2 => 
                           n61930, A => n7331, ZN => n7328);
   U6547 : OAI221_X1 port map( B1 => n52972, B2 => n61719, C1 => n52996, C2 => 
                           n61721, A => n1531, ZN => n7326);
   U6548 : NOR4_X1 port map( A1 => n7176, A2 => n7177, A3 => n7178, A4 => n7179
                           , ZN => n7166);
   U6549 : OAI221_X1 port map( B1 => n53162, B2 => n61922, C1 => n61919, C2 => 
                           n3151, A => n7182, ZN => n7177);
   U6550 : OAI221_X1 port map( B1 => n3423, B2 => n61933, C1 => n3447, C2 => 
                           n61930, A => n7181, ZN => n7178);
   U6551 : OAI221_X1 port map( B1 => n52970, B2 => n61719, C1 => n52994, C2 => 
                           n61721, A => n1527, ZN => n7176);
   U6552 : NOR4_X1 port map( A1 => n6951, A2 => n6952, A3 => n6953, A4 => n6954
                           , ZN => n6941);
   U6553 : OAI221_X1 port map( B1 => n53159, B2 => n61922, C1 => n53183, C2 => 
                           n61918, A => n6957, ZN => n6952);
   U6554 : OAI221_X1 port map( B1 => n3420, B2 => n61934, C1 => n3444, C2 => 
                           n61931, A => n6956, ZN => n6953);
   U6555 : OAI221_X1 port map( B1 => n52967, B2 => n6034, C1 => n52991, C2 => 
                           n6033, A => n1521, ZN => n6951);
   U6556 : NOR4_X1 port map( A1 => n6079, A2 => n6080, A3 => n6081, A4 => n6082
                           , ZN => n6065);
   U6557 : OAI221_X1 port map( B1 => n61827, B2 => n260, C1 => n61824, C2 => 
                           n252, A => n6084, ZN => n6081);
   U6558 : OAI221_X1 port map( B1 => n5500, B2 => n4027, C1 => n5501, C2 => 
                           n4019, A => n6087, ZN => n6080);
   U6559 : OAI221_X1 port map( B1 => n52679, B2 => n5492, C1 => n5493, C2 => 
                           n268, A => n6083, ZN => n6082);
   U6560 : NOR4_X1 port map( A1 => n5981, A2 => n5982, A3 => n5983, A4 => n5984
                           , ZN => n5971);
   U6561 : OAI221_X1 port map( B1 => n61827, B2 => n259, C1 => n61824, C2 => 
                           n251, A => n5986, ZN => n5983);
   U6562 : OAI221_X1 port map( B1 => n5500, B2 => n4026, C1 => n5501, C2 => 
                           n4018, A => n5987, ZN => n5982);
   U6563 : OAI221_X1 port map( B1 => n52678, B2 => n5492, C1 => n5493, C2 => 
                           n267, A => n5985, ZN => n5984);
   U6564 : NOR4_X1 port map( A1 => n5906, A2 => n5907, A3 => n5908, A4 => n5909
                           , ZN => n5896);
   U6565 : OAI221_X1 port map( B1 => n61827, B2 => n258, C1 => n61824, C2 => 
                           n250, A => n5911, ZN => n5908);
   U6566 : OAI221_X1 port map( B1 => n5500, B2 => n4025, C1 => n5501, C2 => 
                           n4017, A => n5912, ZN => n5907);
   U6567 : OAI221_X1 port map( B1 => n52677, B2 => n5492, C1 => n5493, C2 => 
                           n266, A => n5910, ZN => n5909);
   U6568 : NOR4_X1 port map( A1 => n5831, A2 => n5832, A3 => n5833, A4 => n5834
                           , ZN => n5821);
   U6569 : OAI221_X1 port map( B1 => n61827, B2 => n257, C1 => n61824, C2 => 
                           n249, A => n5836, ZN => n5833);
   U6570 : OAI221_X1 port map( B1 => n5500, B2 => n4024, C1 => n5501, C2 => 
                           n4016, A => n5837, ZN => n5832);
   U6571 : OAI221_X1 port map( B1 => n52676, B2 => n5492, C1 => n5493, C2 => 
                           n265, A => n5835, ZN => n5834);
   U6572 : NOR4_X1 port map( A1 => n5756, A2 => n5757, A3 => n5758, A4 => n5759
                           , ZN => n5746);
   U6573 : OAI221_X1 port map( B1 => n61827, B2 => n256, C1 => n61824, C2 => 
                           n248, A => n5761, ZN => n5758);
   U6574 : OAI221_X1 port map( B1 => n5500, B2 => n4023, C1 => n5501, C2 => 
                           n4015, A => n5762, ZN => n5757);
   U6575 : OAI221_X1 port map( B1 => n52675, B2 => n5492, C1 => n5493, C2 => 
                           n264, A => n5760, ZN => n5759);
   U6576 : NOR4_X1 port map( A1 => n5681, A2 => n5682, A3 => n5683, A4 => n5684
                           , ZN => n5671);
   U6577 : OAI221_X1 port map( B1 => n61827, B2 => n255, C1 => n61824, C2 => 
                           n247, A => n5686, ZN => n5683);
   U6578 : OAI221_X1 port map( B1 => n5500, B2 => n4022, C1 => n5501, C2 => 
                           n4014, A => n5687, ZN => n5682);
   U6579 : OAI221_X1 port map( B1 => n52674, B2 => n5492, C1 => n5493, C2 => 
                           n263, A => n5685, ZN => n5684);
   U6580 : NOR4_X1 port map( A1 => n5606, A2 => n5607, A3 => n5608, A4 => n5609
                           , ZN => n5596);
   U6581 : OAI221_X1 port map( B1 => n61827, B2 => n254, C1 => n61824, C2 => 
                           n246, A => n5611, ZN => n5608);
   U6582 : OAI221_X1 port map( B1 => n5500, B2 => n4021, C1 => n5501, C2 => 
                           n4013, A => n5612, ZN => n5607);
   U6583 : OAI221_X1 port map( B1 => n52673, B2 => n5492, C1 => n5493, C2 => 
                           n262, A => n5610, ZN => n5609);
   U6584 : NOR4_X1 port map( A1 => n5488, A2 => n5489, A3 => n5490, A4 => n5491
                           , ZN => n5465);
   U6585 : OAI221_X1 port map( B1 => n61827, B2 => n253, C1 => n61824, C2 => 
                           n245, A => n5499, ZN => n5490);
   U6586 : OAI221_X1 port map( B1 => n5500, B2 => n4020, C1 => n5501, C2 => 
                           n4012, A => n5502, ZN => n5489);
   U6587 : OAI221_X1 port map( B1 => n52672, B2 => n5492, C1 => n5493, C2 => 
                           n261, A => n5494, ZN => n5491);
   U6588 : NOR4_X1 port map( A1 => n14380, A2 => n14381, A3 => n14382, A4 => 
                           n14383, ZN => n14370);
   U6589 : OAI221_X1 port map( B1 => n1608, B2 => n61589, C1 => n1530, C2 => 
                           n61586, A => n14386, ZN => n14381);
   U6590 : OAI221_X1 port map( B1 => n1580, B2 => n61601, C1 => n1720, C2 => 
                           n61598, A => n14385, ZN => n14382);
   U6591 : OAI221_X1 port map( B1 => n52971, B2 => n61613, C1 => n52995, C2 => 
                           n61610, A => n14384, ZN => n14383);
   U6592 : NOR4_X1 port map( A1 => n9889, A2 => n9890, A3 => n9891, A4 => n9892
                           , ZN => n9879);
   U6593 : OAI221_X1 port map( B1 => n1607, B2 => n61589, C1 => n1528, C2 => 
                           n61586, A => n9895, ZN => n9890);
   U6594 : OAI221_X1 port map( B1 => n1579, B2 => n61601, C1 => n1719, C2 => 
                           n61598, A => n9894, ZN => n9891);
   U6595 : OAI221_X1 port map( B1 => n52970, B2 => n61613, C1 => n52994, C2 => 
                           n61610, A => n9893, ZN => n9892);
   U6596 : NOR4_X1 port map( A1 => n9814, A2 => n9815, A3 => n9816, A4 => n9817
                           , ZN => n9740);
   U6597 : OAI221_X1 port map( B1 => n1590, B2 => n61589, C1 => n1526, C2 => 
                           n61586, A => n9820, ZN => n9815);
   U6598 : OAI221_X1 port map( B1 => n1578, B2 => n61601, C1 => n1718, C2 => 
                           n61598, A => n9819, ZN => n9816);
   U6599 : OAI221_X1 port map( B1 => n52969, B2 => n61613, C1 => n52993, C2 => 
                           n61610, A => n9818, ZN => n9817);
   U6600 : NOR4_X1 port map( A1 => n9675, A2 => n9676, A3 => n9677, A4 => n9678
                           , ZN => n9665);
   U6601 : OAI221_X1 port map( B1 => n1589, B2 => n61589, C1 => n1524, C2 => 
                           n61586, A => n9681, ZN => n9676);
   U6602 : OAI221_X1 port map( B1 => n1577, B2 => n61601, C1 => n1717, C2 => 
                           n61598, A => n9680, ZN => n9677);
   U6603 : OAI221_X1 port map( B1 => n52968, B2 => n61613, C1 => n52992, C2 => 
                           n61610, A => n9679, ZN => n9678);
   U6604 : NOR4_X1 port map( A1 => n9584, A2 => n9585, A3 => n9586, A4 => n9587
                           , ZN => n9574);
   U6605 : OAI221_X1 port map( B1 => n1558, B2 => n61590, C1 => n1522, C2 => 
                           n61587, A => n9590, ZN => n9585);
   U6606 : OAI221_X1 port map( B1 => n1576, B2 => n61602, C1 => n1716, C2 => 
                           n61599, A => n9589, ZN => n9586);
   U6607 : OAI221_X1 port map( B1 => n52967, B2 => n61614, C1 => n52991, C2 => 
                           n61611, A => n9588, ZN => n9587);
   U6608 : NOR4_X1 port map( A1 => n9509, A2 => n9510, A3 => n9511, A4 => n9512
                           , ZN => n9499);
   U6609 : OAI221_X1 port map( B1 => n1557, B2 => n61590, C1 => n1520, C2 => 
                           n61587, A => n9515, ZN => n9510);
   U6610 : OAI221_X1 port map( B1 => n1575, B2 => n61602, C1 => n1715, C2 => 
                           n61599, A => n9514, ZN => n9511);
   U6611 : OAI221_X1 port map( B1 => n52966, B2 => n61614, C1 => n52990, C2 => 
                           n61611, A => n9513, ZN => n9512);
   U6612 : NOR4_X1 port map( A1 => n9434, A2 => n9435, A3 => n9436, A4 => n9437
                           , ZN => n9424);
   U6613 : OAI221_X1 port map( B1 => n1556, B2 => n61590, C1 => n1517, C2 => 
                           n61587, A => n9440, ZN => n9435);
   U6614 : OAI221_X1 port map( B1 => n1738, B2 => n61602, C1 => n1714, C2 => 
                           n61599, A => n9439, ZN => n9436);
   U6615 : OAI221_X1 port map( B1 => n52965, B2 => n61614, C1 => n52989, C2 => 
                           n61611, A => n9438, ZN => n9437);
   U6616 : NOR4_X1 port map( A1 => n9359, A2 => n9360, A3 => n9361, A4 => n9362
                           , ZN => n9349);
   U6617 : OAI221_X1 port map( B1 => n1555, B2 => n61590, C1 => n1516, C2 => 
                           n61587, A => n9365, ZN => n9360);
   U6618 : OAI221_X1 port map( B1 => n1737, B2 => n61602, C1 => n1713, C2 => 
                           n61599, A => n9364, ZN => n9361);
   U6619 : OAI221_X1 port map( B1 => n52964, B2 => n61614, C1 => n52988, C2 => 
                           n61611, A => n9363, ZN => n9362);
   U6620 : NOR4_X1 port map( A1 => n9220, A2 => n9221, A3 => n9222, A4 => n9223
                           , ZN => n9210);
   U6621 : OAI221_X1 port map( B1 => n1554, B2 => n61590, C1 => n1515, C2 => 
                           n61587, A => n9226, ZN => n9221);
   U6622 : OAI221_X1 port map( B1 => n1736, B2 => n61602, C1 => n1712, C2 => 
                           n61599, A => n9225, ZN => n9222);
   U6623 : OAI221_X1 port map( B1 => n52963, B2 => n61614, C1 => n52987, C2 => 
                           n61611, A => n9224, ZN => n9223);
   U6624 : NOR4_X1 port map( A1 => n9145, A2 => n9146, A3 => n9147, A4 => n9148
                           , ZN => n9135);
   U6625 : OAI221_X1 port map( B1 => n1553, B2 => n61590, C1 => n1514, C2 => 
                           n61587, A => n9151, ZN => n9146);
   U6626 : OAI221_X1 port map( B1 => n1735, B2 => n61602, C1 => n1711, C2 => 
                           n61599, A => n9150, ZN => n9147);
   U6627 : OAI221_X1 port map( B1 => n52962, B2 => n61614, C1 => n52986, C2 => 
                           n61611, A => n9149, ZN => n9148);
   U6628 : NOR4_X1 port map( A1 => n9181, A2 => n9182, A3 => n9183, A4 => n9184
                           , ZN => n9171);
   U6629 : OAI221_X1 port map( B1 => n1908, B2 => n61398, C1 => n1932, C2 => 
                           n61395, A => n9186, ZN => n9183);
   U6630 : OAI221_X1 port map( B1 => n2028, B2 => n61410, C1 => n1980, C2 => 
                           n61407, A => n9185, ZN => n9184);
   U6631 : OAI221_X1 port map( B1 => n1836, B2 => n61386, C1 => n2651, C2 => 
                           n61383, A => n9187, ZN => n9182);
   U6632 : NOR4_X1 port map( A1 => n9070, A2 => n9071, A3 => n9072, A4 => n9073
                           , ZN => n9060);
   U6633 : OAI221_X1 port map( B1 => n1552, B2 => n61590, C1 => n1513, C2 => 
                           n61587, A => n9076, ZN => n9071);
   U6634 : OAI221_X1 port map( B1 => n1734, B2 => n61602, C1 => n1710, C2 => 
                           n61599, A => n9075, ZN => n9072);
   U6635 : OAI221_X1 port map( B1 => n52961, B2 => n61614, C1 => n52985, C2 => 
                           n61611, A => n9074, ZN => n9073);
   U6636 : NOR4_X1 port map( A1 => n9106, A2 => n9107, A3 => n9108, A4 => n9109
                           , ZN => n9096);
   U6637 : OAI221_X1 port map( B1 => n1907, B2 => n61398, C1 => n1931, C2 => 
                           n61395, A => n9111, ZN => n9108);
   U6638 : OAI221_X1 port map( B1 => n2027, B2 => n61410, C1 => n1979, C2 => 
                           n61407, A => n9110, ZN => n9109);
   U6639 : OAI221_X1 port map( B1 => n1835, B2 => n61386, C1 => n2650, C2 => 
                           n61383, A => n9112, ZN => n9107);
   U6640 : NOR4_X1 port map( A1 => n8995, A2 => n8996, A3 => n8997, A4 => n8998
                           , ZN => n8985);
   U6641 : OAI221_X1 port map( B1 => n1551, B2 => n61590, C1 => n1512, C2 => 
                           n61587, A => n9001, ZN => n8996);
   U6642 : OAI221_X1 port map( B1 => n1733, B2 => n61602, C1 => n1709, C2 => 
                           n61599, A => n9000, ZN => n8997);
   U6643 : OAI221_X1 port map( B1 => n52960, B2 => n61614, C1 => n52984, C2 => 
                           n61611, A => n8999, ZN => n8998);
   U6644 : NOR4_X1 port map( A1 => n9031, A2 => n9032, A3 => n9033, A4 => n9034
                           , ZN => n9021);
   U6645 : OAI221_X1 port map( B1 => n1906, B2 => n61398, C1 => n1930, C2 => 
                           n61395, A => n9036, ZN => n9033);
   U6646 : OAI221_X1 port map( B1 => n2026, B2 => n61410, C1 => n1978, C2 => 
                           n61407, A => n9035, ZN => n9034);
   U6647 : OAI221_X1 port map( B1 => n1834, B2 => n61386, C1 => n2649, C2 => 
                           n61383, A => n9037, ZN => n9032);
   U6648 : NOR4_X1 port map( A1 => n8920, A2 => n8921, A3 => n8922, A4 => n8923
                           , ZN => n8910);
   U6649 : OAI221_X1 port map( B1 => n1550, B2 => n61590, C1 => n1511, C2 => 
                           n61587, A => n8926, ZN => n8921);
   U6650 : OAI221_X1 port map( B1 => n1732, B2 => n61602, C1 => n1708, C2 => 
                           n61599, A => n8925, ZN => n8922);
   U6651 : OAI221_X1 port map( B1 => n52959, B2 => n61614, C1 => n52983, C2 => 
                           n61611, A => n8924, ZN => n8923);
   U6652 : NOR4_X1 port map( A1 => n8956, A2 => n8957, A3 => n8958, A4 => n8959
                           , ZN => n8946);
   U6653 : OAI221_X1 port map( B1 => n1905, B2 => n61398, C1 => n1929, C2 => 
                           n61395, A => n8961, ZN => n8958);
   U6654 : OAI221_X1 port map( B1 => n2025, B2 => n61410, C1 => n1977, C2 => 
                           n61407, A => n8960, ZN => n8959);
   U6655 : OAI221_X1 port map( B1 => n1833, B2 => n61386, C1 => n2648, C2 => 
                           n61383, A => n8962, ZN => n8957);
   U6656 : NOR4_X1 port map( A1 => n8845, A2 => n8846, A3 => n8847, A4 => n8848
                           , ZN => n8835);
   U6657 : OAI221_X1 port map( B1 => n1549, B2 => n61590, C1 => n1510, C2 => 
                           n61587, A => n8851, ZN => n8846);
   U6658 : OAI221_X1 port map( B1 => n1731, B2 => n61602, C1 => n1707, C2 => 
                           n61599, A => n8850, ZN => n8847);
   U6659 : OAI221_X1 port map( B1 => n52958, B2 => n61614, C1 => n52982, C2 => 
                           n61611, A => n8849, ZN => n8848);
   U6660 : NOR4_X1 port map( A1 => n8881, A2 => n8882, A3 => n8883, A4 => n8884
                           , ZN => n8871);
   U6661 : OAI221_X1 port map( B1 => n1904, B2 => n61398, C1 => n1928, C2 => 
                           n61395, A => n8886, ZN => n8883);
   U6662 : OAI221_X1 port map( B1 => n2024, B2 => n61410, C1 => n1976, C2 => 
                           n61407, A => n8885, ZN => n8884);
   U6663 : OAI221_X1 port map( B1 => n1832, B2 => n61386, C1 => n2647, C2 => 
                           n61383, A => n8887, ZN => n8882);
   U6664 : NOR4_X1 port map( A1 => n8770, A2 => n8771, A3 => n8772, A4 => n8773
                           , ZN => n8760);
   U6665 : OAI221_X1 port map( B1 => n1548, B2 => n61590, C1 => n1509, C2 => 
                           n61587, A => n8776, ZN => n8771);
   U6666 : OAI221_X1 port map( B1 => n1730, B2 => n61602, C1 => n1706, C2 => 
                           n61599, A => n8775, ZN => n8772);
   U6667 : OAI221_X1 port map( B1 => n52957, B2 => n61614, C1 => n52981, C2 => 
                           n61611, A => n8774, ZN => n8773);
   U6668 : NOR4_X1 port map( A1 => n8806, A2 => n8807, A3 => n8808, A4 => n8809
                           , ZN => n8796);
   U6669 : OAI221_X1 port map( B1 => n1903, B2 => n61398, C1 => n1927, C2 => 
                           n61395, A => n8811, ZN => n8808);
   U6670 : OAI221_X1 port map( B1 => n2023, B2 => n61410, C1 => n1975, C2 => 
                           n61407, A => n8810, ZN => n8809);
   U6671 : OAI221_X1 port map( B1 => n1831, B2 => n61386, C1 => n2646, C2 => 
                           n61383, A => n8812, ZN => n8807);
   U6672 : NOR4_X1 port map( A1 => n8695, A2 => n8696, A3 => n8697, A4 => n8698
                           , ZN => n8685);
   U6673 : OAI221_X1 port map( B1 => n1547, B2 => n61590, C1 => n1508, C2 => 
                           n61587, A => n8701, ZN => n8696);
   U6674 : OAI221_X1 port map( B1 => n1729, B2 => n61602, C1 => n1705, C2 => 
                           n61599, A => n8700, ZN => n8697);
   U6675 : OAI221_X1 port map( B1 => n52956, B2 => n61614, C1 => n52980, C2 => 
                           n61611, A => n8699, ZN => n8698);
   U6676 : NOR4_X1 port map( A1 => n8731, A2 => n8732, A3 => n8733, A4 => n8734
                           , ZN => n8721);
   U6677 : OAI221_X1 port map( B1 => n1902, B2 => n61398, C1 => n1926, C2 => 
                           n61395, A => n8736, ZN => n8733);
   U6678 : OAI221_X1 port map( B1 => n1998, B2 => n61410, C1 => n1974, C2 => 
                           n61407, A => n8735, ZN => n8734);
   U6679 : OAI221_X1 port map( B1 => n1830, B2 => n61386, C1 => n2645, C2 => 
                           n61383, A => n8737, ZN => n8732);
   U6680 : NOR4_X1 port map( A1 => n14994, A2 => n14995, A3 => n14996, A4 => 
                           n14997, ZN => n14970);
   U6681 : OAI221_X1 port map( B1 => n1616, B2 => n61589, C1 => n1546, C2 => 
                           n61586, A => n15002, ZN => n14995);
   U6682 : OAI221_X1 port map( B1 => n1588, B2 => n61601, C1 => n1728, C2 => 
                           n61598, A => n14999, ZN => n14996);
   U6683 : OAI221_X1 port map( B1 => n52979, B2 => n61613, C1 => n53003, C2 => 
                           n61610, A => n14998, ZN => n14997);
   U6684 : NOR4_X1 port map( A1 => n15042, A2 => n15043, A3 => n15044, A4 => 
                           n15045, ZN => n15029);
   U6685 : OAI221_X1 port map( B1 => n1925, B2 => n61397, C1 => n1949, C2 => 
                           n61394, A => n15048, ZN => n15044);
   U6686 : OAI221_X1 port map( B1 => n2045, B2 => n61409, C1 => n1997, C2 => 
                           n61406, A => n15046, ZN => n15045);
   U6687 : OAI221_X1 port map( B1 => n164, B2 => n61385, C1 => n1829, C2 => 
                           n61382, A => n15049, ZN => n15043);
   U6688 : NOR4_X1 port map( A1 => n14905, A2 => n14906, A3 => n14907, A4 => 
                           n14908, ZN => n14895);
   U6689 : OAI221_X1 port map( B1 => n1615, B2 => n61589, C1 => n1544, C2 => 
                           n61586, A => n14911, ZN => n14906);
   U6690 : OAI221_X1 port map( B1 => n1587, B2 => n61601, C1 => n1727, C2 => 
                           n61598, A => n14910, ZN => n14907);
   U6691 : OAI221_X1 port map( B1 => n52978, B2 => n61613, C1 => n53002, C2 => 
                           n61610, A => n14909, ZN => n14908);
   U6692 : NOR4_X1 port map( A1 => n14941, A2 => n14942, A3 => n14943, A4 => 
                           n14944, ZN => n14931);
   U6693 : OAI221_X1 port map( B1 => n1924, B2 => n61397, C1 => n1948, C2 => 
                           n61394, A => n14946, ZN => n14943);
   U6694 : OAI221_X1 port map( B1 => n2044, B2 => n61409, C1 => n1996, C2 => 
                           n61406, A => n14945, ZN => n14944);
   U6695 : OAI221_X1 port map( B1 => n163, B2 => n61385, C1 => n1828, C2 => 
                           n61382, A => n14947, ZN => n14942);
   U6696 : NOR4_X1 port map( A1 => n14830, A2 => n14831, A3 => n14832, A4 => 
                           n14833, ZN => n14820);
   U6697 : OAI221_X1 port map( B1 => n1614, B2 => n61589, C1 => n1542, C2 => 
                           n61586, A => n14836, ZN => n14831);
   U6698 : OAI221_X1 port map( B1 => n1586, B2 => n61601, C1 => n1726, C2 => 
                           n61598, A => n14835, ZN => n14832);
   U6699 : OAI221_X1 port map( B1 => n52977, B2 => n61613, C1 => n53001, C2 => 
                           n61610, A => n14834, ZN => n14833);
   U6700 : NOR4_X1 port map( A1 => n14866, A2 => n14867, A3 => n14868, A4 => 
                           n14869, ZN => n14856);
   U6701 : OAI221_X1 port map( B1 => n1923, B2 => n61397, C1 => n1947, C2 => 
                           n61394, A => n14871, ZN => n14868);
   U6702 : OAI221_X1 port map( B1 => n2043, B2 => n61409, C1 => n1995, C2 => 
                           n61406, A => n14870, ZN => n14869);
   U6703 : OAI221_X1 port map( B1 => n162, B2 => n61385, C1 => n1827, C2 => 
                           n61382, A => n14872, ZN => n14867);
   U6704 : NOR4_X1 port map( A1 => n14755, A2 => n14756, A3 => n14757, A4 => 
                           n14758, ZN => n14745);
   U6705 : OAI221_X1 port map( B1 => n1613, B2 => n61589, C1 => n1540, C2 => 
                           n61586, A => n14761, ZN => n14756);
   U6706 : OAI221_X1 port map( B1 => n1585, B2 => n61601, C1 => n1725, C2 => 
                           n61598, A => n14760, ZN => n14757);
   U6707 : OAI221_X1 port map( B1 => n52976, B2 => n61613, C1 => n53000, C2 => 
                           n61610, A => n14759, ZN => n14758);
   U6708 : NOR4_X1 port map( A1 => n14791, A2 => n14792, A3 => n14793, A4 => 
                           n14794, ZN => n14781);
   U6709 : OAI221_X1 port map( B1 => n1922, B2 => n61397, C1 => n1946, C2 => 
                           n61394, A => n14796, ZN => n14793);
   U6710 : OAI221_X1 port map( B1 => n2042, B2 => n61409, C1 => n1994, C2 => 
                           n61406, A => n14795, ZN => n14794);
   U6711 : OAI221_X1 port map( B1 => n161, B2 => n61385, C1 => n1826, C2 => 
                           n61382, A => n14797, ZN => n14792);
   U6712 : NOR4_X1 port map( A1 => n14680, A2 => n14681, A3 => n14682, A4 => 
                           n14683, ZN => n14670);
   U6713 : OAI221_X1 port map( B1 => n1612, B2 => n61589, C1 => n1538, C2 => 
                           n61586, A => n14686, ZN => n14681);
   U6714 : OAI221_X1 port map( B1 => n1584, B2 => n61601, C1 => n1724, C2 => 
                           n61598, A => n14685, ZN => n14682);
   U6715 : OAI221_X1 port map( B1 => n52975, B2 => n61613, C1 => n52999, C2 => 
                           n61610, A => n14684, ZN => n14683);
   U6716 : NOR4_X1 port map( A1 => n14716, A2 => n14717, A3 => n14718, A4 => 
                           n14719, ZN => n14706);
   U6717 : OAI221_X1 port map( B1 => n1921, B2 => n61397, C1 => n1945, C2 => 
                           n61394, A => n14721, ZN => n14718);
   U6718 : OAI221_X1 port map( B1 => n2041, B2 => n61409, C1 => n1993, C2 => 
                           n61406, A => n14720, ZN => n14719);
   U6719 : OAI221_X1 port map( B1 => n160, B2 => n61385, C1 => n1825, C2 => 
                           n61382, A => n14722, ZN => n14717);
   U6720 : NOR4_X1 port map( A1 => n14605, A2 => n14606, A3 => n14607, A4 => 
                           n14608, ZN => n14595);
   U6721 : OAI221_X1 port map( B1 => n1611, B2 => n61589, C1 => n1536, C2 => 
                           n61586, A => n14611, ZN => n14606);
   U6722 : OAI221_X1 port map( B1 => n1583, B2 => n61601, C1 => n1723, C2 => 
                           n61598, A => n14610, ZN => n14607);
   U6723 : OAI221_X1 port map( B1 => n52974, B2 => n61613, C1 => n52998, C2 => 
                           n61610, A => n14609, ZN => n14608);
   U6724 : NOR4_X1 port map( A1 => n14530, A2 => n14531, A3 => n14532, A4 => 
                           n14533, ZN => n14520);
   U6725 : OAI221_X1 port map( B1 => n1610, B2 => n61589, C1 => n1534, C2 => 
                           n61586, A => n14536, ZN => n14531);
   U6726 : OAI221_X1 port map( B1 => n1582, B2 => n61601, C1 => n1722, C2 => 
                           n61598, A => n14535, ZN => n14532);
   U6727 : OAI221_X1 port map( B1 => n52973, B2 => n61613, C1 => n52997, C2 => 
                           n61610, A => n14534, ZN => n14533);
   U6728 : NOR4_X1 port map( A1 => n14455, A2 => n14456, A3 => n14457, A4 => 
                           n14458, ZN => n14445);
   U6729 : OAI221_X1 port map( B1 => n1609, B2 => n61589, C1 => n1532, C2 => 
                           n61586, A => n14461, ZN => n14456);
   U6730 : OAI221_X1 port map( B1 => n1581, B2 => n61601, C1 => n1721, C2 => 
                           n61598, A => n14460, ZN => n14457);
   U6731 : OAI221_X1 port map( B1 => n52972, B2 => n61613, C1 => n52996, C2 => 
                           n61610, A => n14459, ZN => n14458);
   U6732 : NOR4_X1 port map( A1 => n8620, A2 => n8621, A3 => n8622, A4 => n8623
                           , ZN => n8610);
   U6733 : OAI221_X1 port map( B1 => n67, B2 => n61591, C1 => n59, C2 => n61588
                           , A => n8626, ZN => n8621);
   U6734 : OAI221_X1 port map( B1 => n831, B2 => n61603, C1 => n823, C2 => 
                           n61600, A => n8625, ZN => n8622);
   U6735 : OAI221_X1 port map( B1 => n4003, B2 => n61615, C1 => n4011, C2 => 
                           n61612, A => n8624, ZN => n8623);
   U6736 : NOR4_X1 port map( A1 => n8545, A2 => n8546, A3 => n8547, A4 => n8548
                           , ZN => n8535);
   U6737 : OAI221_X1 port map( B1 => n66, B2 => n61591, C1 => n58, C2 => n61588
                           , A => n8551, ZN => n8546);
   U6738 : OAI221_X1 port map( B1 => n830, B2 => n61603, C1 => n822, C2 => 
                           n61600, A => n8550, ZN => n8547);
   U6739 : OAI221_X1 port map( B1 => n4002, B2 => n61615, C1 => n4010, C2 => 
                           n61612, A => n8549, ZN => n8548);
   U6740 : NOR4_X1 port map( A1 => n8470, A2 => n8471, A3 => n8472, A4 => n8473
                           , ZN => n8460);
   U6741 : OAI221_X1 port map( B1 => n65, B2 => n61591, C1 => n57, C2 => n61588
                           , A => n8476, ZN => n8471);
   U6742 : OAI221_X1 port map( B1 => n829, B2 => n61603, C1 => n821, C2 => 
                           n61600, A => n8475, ZN => n8472);
   U6743 : OAI221_X1 port map( B1 => n4001, B2 => n61615, C1 => n4009, C2 => 
                           n61612, A => n8474, ZN => n8473);
   U6744 : NOR4_X1 port map( A1 => n8395, A2 => n8396, A3 => n8397, A4 => n8398
                           , ZN => n8385);
   U6745 : OAI221_X1 port map( B1 => n64, B2 => n61591, C1 => n56, C2 => n61588
                           , A => n8401, ZN => n8396);
   U6746 : OAI221_X1 port map( B1 => n828, B2 => n61603, C1 => n820, C2 => 
                           n61600, A => n8400, ZN => n8397);
   U6747 : OAI221_X1 port map( B1 => n4000, B2 => n61615, C1 => n4008, C2 => 
                           n61612, A => n8399, ZN => n8398);
   U6748 : NOR4_X1 port map( A1 => n8320, A2 => n8321, A3 => n8322, A4 => n8323
                           , ZN => n8310);
   U6749 : OAI221_X1 port map( B1 => n63, B2 => n61591, C1 => n55, C2 => n61588
                           , A => n8326, ZN => n8321);
   U6750 : OAI221_X1 port map( B1 => n827, B2 => n61603, C1 => n819, C2 => 
                           n61600, A => n8325, ZN => n8322);
   U6751 : OAI221_X1 port map( B1 => n3999, B2 => n61615, C1 => n4007, C2 => 
                           n61612, A => n8324, ZN => n8323);
   U6752 : NOR4_X1 port map( A1 => n8245, A2 => n8246, A3 => n8247, A4 => n8248
                           , ZN => n8235);
   U6753 : OAI221_X1 port map( B1 => n62, B2 => n61591, C1 => n54, C2 => n61588
                           , A => n8251, ZN => n8246);
   U6754 : OAI221_X1 port map( B1 => n826, B2 => n61603, C1 => n818, C2 => 
                           n61600, A => n8250, ZN => n8247);
   U6755 : OAI221_X1 port map( B1 => n3998, B2 => n61615, C1 => n4006, C2 => 
                           n61612, A => n8249, ZN => n8248);
   U6756 : NOR4_X1 port map( A1 => n8170, A2 => n8171, A3 => n8172, A4 => n8173
                           , ZN => n8160);
   U6757 : OAI221_X1 port map( B1 => n61, B2 => n61591, C1 => n53, C2 => n61588
                           , A => n8176, ZN => n8171);
   U6758 : OAI221_X1 port map( B1 => n825, B2 => n61603, C1 => n817, C2 => 
                           n61600, A => n8175, ZN => n8172);
   U6759 : OAI221_X1 port map( B1 => n3997, B2 => n61615, C1 => n4005, C2 => 
                           n61612, A => n8174, ZN => n8173);
   U6760 : NOR4_X1 port map( A1 => n7976, A2 => n7977, A3 => n7978, A4 => n7979
                           , ZN => n7949);
   U6761 : OAI221_X1 port map( B1 => n60, B2 => n61591, C1 => n52, C2 => n61588
                           , A => n7992, ZN => n7977);
   U6762 : OAI221_X1 port map( B1 => n824, B2 => n61603, C1 => n816, C2 => 
                           n61600, A => n7987, ZN => n7978);
   U6763 : OAI221_X1 port map( B1 => n3996, B2 => n61615, C1 => n4004, C2 => 
                           n61612, A => n7982, ZN => n7979);
   U6764 : NOR4_X1 port map( A1 => n6026, A2 => n6027, A3 => n6028, A4 => n6029
                           , ZN => n6010);
   U6765 : OAI221_X1 port map( B1 => n59744, B2 => n67, C1 => n59739, C2 => n59
                           , A => n6032, ZN => n6027);
   U6766 : OAI221_X1 port map( B1 => n61921, B2 => n974, C1 => n61919, C2 => 
                           n982, A => n6031, ZN => n6028);
   U6767 : OAI221_X1 port map( B1 => n2916, B2 => n61935, C1 => n2924, C2 => 
                           n61932, A => n6030, ZN => n6029);
   U6768 : NOR4_X1 port map( A1 => n5945, A2 => n5946, A3 => n5947, A4 => n5948
                           , ZN => n5935);
   U6769 : OAI221_X1 port map( B1 => n59745, B2 => n66, C1 => n59739, C2 => n58
                           , A => n5951, ZN => n5946);
   U6770 : OAI221_X1 port map( B1 => n61921, B2 => n973, C1 => n61919, C2 => 
                           n981, A => n5950, ZN => n5947);
   U6771 : OAI221_X1 port map( B1 => n2915, B2 => n61935, C1 => n2923, C2 => 
                           n61932, A => n5949, ZN => n5948);
   U6772 : NOR4_X1 port map( A1 => n5870, A2 => n5871, A3 => n5872, A4 => n5873
                           , ZN => n5860);
   U6773 : OAI221_X1 port map( B1 => n59744, B2 => n65, C1 => n59737, C2 => n57
                           , A => n5876, ZN => n5871);
   U6774 : OAI221_X1 port map( B1 => n61921, B2 => n972, C1 => n61919, C2 => 
                           n980, A => n5875, ZN => n5872);
   U6775 : OAI221_X1 port map( B1 => n2914, B2 => n61935, C1 => n2922, C2 => 
                           n61932, A => n5874, ZN => n5873);
   U6776 : NOR4_X1 port map( A1 => n5795, A2 => n5796, A3 => n5797, A4 => n5798
                           , ZN => n5785);
   U6777 : OAI221_X1 port map( B1 => n59745, B2 => n64, C1 => n59737, C2 => n56
                           , A => n5801, ZN => n5796);
   U6778 : OAI221_X1 port map( B1 => n61921, B2 => n815, C1 => n61919, C2 => 
                           n979, A => n5800, ZN => n5797);
   U6779 : OAI221_X1 port map( B1 => n2913, B2 => n61935, C1 => n2921, C2 => 
                           n61932, A => n5799, ZN => n5798);
   U6780 : NOR4_X1 port map( A1 => n5720, A2 => n5721, A3 => n5722, A4 => n5723
                           , ZN => n5710);
   U6781 : OAI221_X1 port map( B1 => n59746, B2 => n63, C1 => n59738, C2 => n55
                           , A => n5726, ZN => n5721);
   U6782 : OAI221_X1 port map( B1 => n61921, B2 => n814, C1 => n61919, C2 => 
                           n978, A => n5725, ZN => n5722);
   U6783 : OAI221_X1 port map( B1 => n2912, B2 => n61935, C1 => n2920, C2 => 
                           n61932, A => n5724, ZN => n5723);
   U6784 : NOR4_X1 port map( A1 => n5645, A2 => n5646, A3 => n5647, A4 => n5648
                           , ZN => n5635);
   U6785 : OAI221_X1 port map( B1 => n59747, B2 => n62, C1 => n59739, C2 => n54
                           , A => n5651, ZN => n5646);
   U6786 : OAI221_X1 port map( B1 => n61921, B2 => n813, C1 => n61919, C2 => 
                           n977, A => n5650, ZN => n5647);
   U6787 : OAI221_X1 port map( B1 => n2911, B2 => n61935, C1 => n2919, C2 => 
                           n61932, A => n5649, ZN => n5648);
   U6788 : NOR4_X1 port map( A1 => n5570, A2 => n5571, A3 => n5572, A4 => n5573
                           , ZN => n5560);
   U6789 : OAI221_X1 port map( B1 => n59746, B2 => n61, C1 => n59738, C2 => n53
                           , A => n5576, ZN => n5571);
   U6790 : OAI221_X1 port map( B1 => n61921, B2 => n812, C1 => n61919, C2 => 
                           n976, A => n5575, ZN => n5572);
   U6791 : OAI221_X1 port map( B1 => n2910, B2 => n61935, C1 => n2918, C2 => 
                           n61932, A => n5574, ZN => n5573);
   U6792 : NOR4_X1 port map( A1 => n5401, A2 => n5402, A3 => n5403, A4 => n5404
                           , ZN => n5380);
   U6793 : OAI221_X1 port map( B1 => n59747, B2 => n60, C1 => n59737, C2 => n52
                           , A => n5417, ZN => n5402);
   U6794 : OAI221_X1 port map( B1 => n61921, B2 => n811, C1 => n61919, C2 => 
                           n975, A => n5412, ZN => n5403);
   U6795 : OAI221_X1 port map( B1 => n2909, B2 => n61935, C1 => n2917, C2 => 
                           n61932, A => n5407, ZN => n5404);
   U6796 : NOR4_X1 port map( A1 => n6734, A2 => n6735, A3 => n6736, A4 => n6737
                           , ZN => n6715);
   U6797 : OAI221_X1 port map( B1 => n61900, B2 => n2685, C1 => n61898, C2 => 
                           n2709, A => n6739, ZN => n6736);
   U6798 : OAI221_X1 port map( B1 => n2007, B2 => n6044, C1 => n3629, C2 => 
                           n61716, A => n6740, ZN => n6735);
   U6799 : OAI221_X1 port map( B1 => n6062, B2 => n3039, C1 => n53036, C2 => 
                           n61700, A => n6738, ZN => n6737);
   U6800 : NOR4_X1 port map( A1 => n6659, A2 => n6660, A3 => n6661, A4 => n6662
                           , ZN => n6640);
   U6801 : OAI221_X1 port map( B1 => n61900, B2 => n2684, C1 => n61898, C2 => 
                           n2708, A => n6664, ZN => n6661);
   U6802 : OAI221_X1 port map( B1 => n2006, B2 => n6044, C1 => n3628, C2 => 
                           n61716, A => n6665, ZN => n6660);
   U6803 : OAI221_X1 port map( B1 => n6062, B2 => n3038, C1 => n53035, C2 => 
                           n61700, A => n6663, ZN => n6662);
   U6804 : NOR4_X1 port map( A1 => n6584, A2 => n6585, A3 => n6586, A4 => n6587
                           , ZN => n6565);
   U6805 : OAI221_X1 port map( B1 => n61900, B2 => n2683, C1 => n61898, C2 => 
                           n2707, A => n6589, ZN => n6586);
   U6806 : OAI221_X1 port map( B1 => n2005, B2 => n6044, C1 => n3627, C2 => 
                           n61716, A => n6590, ZN => n6585);
   U6807 : OAI221_X1 port map( B1 => n6062, B2 => n3037, C1 => n53034, C2 => 
                           n61700, A => n6588, ZN => n6587);
   U6808 : NOR4_X1 port map( A1 => n6509, A2 => n6510, A3 => n6511, A4 => n6512
                           , ZN => n6490);
   U6809 : OAI221_X1 port map( B1 => n61900, B2 => n2682, C1 => n61898, C2 => 
                           n2706, A => n6514, ZN => n6511);
   U6810 : OAI221_X1 port map( B1 => n2004, B2 => n6044, C1 => n3626, C2 => 
                           n61716, A => n6515, ZN => n6510);
   U6811 : OAI221_X1 port map( B1 => n6062, B2 => n3036, C1 => n53033, C2 => 
                           n61700, A => n6513, ZN => n6512);
   U6812 : NOR4_X1 port map( A1 => n6434, A2 => n6435, A3 => n6436, A4 => n6437
                           , ZN => n6415);
   U6813 : OAI221_X1 port map( B1 => n61900, B2 => n2681, C1 => n61898, C2 => 
                           n2705, A => n6439, ZN => n6436);
   U6814 : OAI221_X1 port map( B1 => n2003, B2 => n6044, C1 => n3625, C2 => 
                           n61716, A => n6440, ZN => n6435);
   U6815 : OAI221_X1 port map( B1 => n6062, B2 => n3035, C1 => n53032, C2 => 
                           n61700, A => n6438, ZN => n6437);
   U6816 : NOR4_X1 port map( A1 => n6359, A2 => n6360, A3 => n6361, A4 => n6362
                           , ZN => n6340);
   U6817 : OAI221_X1 port map( B1 => n61900, B2 => n2680, C1 => n61897, C2 => 
                           n2704, A => n6364, ZN => n6361);
   U6818 : OAI221_X1 port map( B1 => n2002, B2 => n6044, C1 => n3624, C2 => 
                           n61716, A => n6365, ZN => n6360);
   U6819 : OAI221_X1 port map( B1 => n6062, B2 => n3034, C1 => n53031, C2 => 
                           n61700, A => n6363, ZN => n6362);
   U6820 : NOR4_X1 port map( A1 => n6284, A2 => n6285, A3 => n6286, A4 => n6287
                           , ZN => n6265);
   U6821 : OAI221_X1 port map( B1 => n61900, B2 => n2679, C1 => n61897, C2 => 
                           n2703, A => n6289, ZN => n6286);
   U6822 : OAI221_X1 port map( B1 => n2001, B2 => n6044, C1 => n3623, C2 => 
                           n61716, A => n6290, ZN => n6285);
   U6823 : OAI221_X1 port map( B1 => n6062, B2 => n3033, C1 => n53030, C2 => 
                           n61700, A => n6288, ZN => n6287);
   U6824 : NOR4_X1 port map( A1 => n6209, A2 => n6210, A3 => n6211, A4 => n6212
                           , ZN => n6190);
   U6825 : OAI221_X1 port map( B1 => n61900, B2 => n2678, C1 => n61897, C2 => 
                           n2702, A => n6214, ZN => n6211);
   U6826 : OAI221_X1 port map( B1 => n2000, B2 => n6044, C1 => n3622, C2 => 
                           n61716, A => n6215, ZN => n6210);
   U6827 : OAI221_X1 port map( B1 => n6062, B2 => n3032, C1 => n53029, C2 => 
                           n61700, A => n6213, ZN => n6212);
   U6828 : NOR4_X1 port map( A1 => n6134, A2 => n6135, A3 => n6136, A4 => n6137
                           , ZN => n6115);
   U6829 : OAI221_X1 port map( B1 => n61900, B2 => n2677, C1 => n61897, C2 => 
                           n2701, A => n6139, ZN => n6136);
   U6830 : OAI221_X1 port map( B1 => n1999, B2 => n6044, C1 => n3621, C2 => 
                           n61716, A => n6140, ZN => n6135);
   U6831 : OAI221_X1 port map( B1 => n6062, B2 => n3031, C1 => n53028, C2 => 
                           n61700, A => n6138, ZN => n6137);
   U6832 : NOR4_X1 port map( A1 => n7109, A2 => n7110, A3 => n7111, A4 => n7112
                           , ZN => n7090);
   U6833 : OAI221_X1 port map( B1 => n81, B2 => n61901, C1 => n61898, C2 => 
                           n2714, A => n7114, ZN => n7111);
   U6834 : OAI221_X1 port map( B1 => n2012, B2 => n61713, C1 => n3634, C2 => 
                           n61715, A => n7115, ZN => n7110);
   U6835 : OAI221_X1 port map( B1 => n61697, B2 => n3044, C1 => n53041, C2 => 
                           n61699, A => n7113, ZN => n7112);
   U6836 : NOR4_X1 port map( A1 => n7034, A2 => n7035, A3 => n7036, A4 => n7037
                           , ZN => n7015);
   U6837 : OAI221_X1 port map( B1 => n80, B2 => n61901, C1 => n61898, C2 => 
                           n2713, A => n7039, ZN => n7036);
   U6838 : OAI221_X1 port map( B1 => n2011, B2 => n61713, C1 => n3633, C2 => 
                           n61715, A => n7040, ZN => n7035);
   U6839 : OAI221_X1 port map( B1 => n61697, B2 => n3043, C1 => n53040, C2 => 
                           n61699, A => n7038, ZN => n7037);
   U6840 : NOR4_X1 port map( A1 => n6884, A2 => n6885, A3 => n6886, A4 => n6887
                           , ZN => n6865);
   U6841 : OAI221_X1 port map( B1 => n61900, B2 => n2687, C1 => n61898, C2 => 
                           n2711, A => n6889, ZN => n6886);
   U6842 : OAI221_X1 port map( B1 => n2009, B2 => n6044, C1 => n3631, C2 => 
                           n61716, A => n6890, ZN => n6885);
   U6843 : OAI221_X1 port map( B1 => n6062, B2 => n3041, C1 => n53038, C2 => 
                           n61700, A => n6888, ZN => n6887);
   U6844 : NOR4_X1 port map( A1 => n6809, A2 => n6810, A3 => n6811, A4 => n6812
                           , ZN => n6790);
   U6845 : OAI221_X1 port map( B1 => n61900, B2 => n2686, C1 => n61898, C2 => 
                           n2710, A => n6814, ZN => n6811);
   U6846 : OAI221_X1 port map( B1 => n2008, B2 => n6044, C1 => n3630, C2 => 
                           n61716, A => n6815, ZN => n6810);
   U6847 : OAI221_X1 port map( B1 => n6062, B2 => n3040, C1 => n53037, C2 => 
                           n61700, A => n6813, ZN => n6812);
   U6848 : NOR4_X1 port map( A1 => n7259, A2 => n7260, A3 => n7261, A4 => n7262
                           , ZN => n7240);
   U6849 : OAI221_X1 port map( B1 => n83, B2 => n61901, C1 => n61898, C2 => 
                           n2716, A => n7264, ZN => n7261);
   U6850 : OAI221_X1 port map( B1 => n2014, B2 => n61713, C1 => n3636, C2 => 
                           n61715, A => n7265, ZN => n7260);
   U6851 : OAI221_X1 port map( B1 => n61697, B2 => n3046, C1 => n53043, C2 => 
                           n61699, A => n7263, ZN => n7262);
   U6852 : NOR4_X1 port map( A1 => n7878, A2 => n7879, A3 => n7880, A4 => n7881
                           , ZN => n7840);
   U6853 : OAI221_X1 port map( B1 => n91, B2 => n61901, C1 => n61899, C2 => 
                           n2724, A => n7884, ZN => n7880);
   U6854 : OAI221_X1 port map( B1 => n2022, B2 => n61713, C1 => n3644, C2 => 
                           n61715, A => n7887, ZN => n7879);
   U6855 : OAI221_X1 port map( B1 => n61697, B2 => n3054, C1 => n53051, C2 => 
                           n61699, A => n7882, ZN => n7881);
   U6856 : NOR4_X1 port map( A1 => n7784, A2 => n7785, A3 => n7786, A4 => n7787
                           , ZN => n7765);
   U6857 : OAI221_X1 port map( B1 => n90, B2 => n61902, C1 => n61899, C2 => 
                           n2723, A => n7789, ZN => n7786);
   U6858 : OAI221_X1 port map( B1 => n2021, B2 => n61713, C1 => n3643, C2 => 
                           n61715, A => n7790, ZN => n7785);
   U6859 : OAI221_X1 port map( B1 => n61697, B2 => n3053, C1 => n53050, C2 => 
                           n61699, A => n7788, ZN => n7787);
   U6860 : NOR4_X1 port map( A1 => n7709, A2 => n7710, A3 => n7711, A4 => n7712
                           , ZN => n7690);
   U6861 : OAI221_X1 port map( B1 => n89, B2 => n61902, C1 => n61899, C2 => 
                           n2722, A => n7714, ZN => n7711);
   U6862 : OAI221_X1 port map( B1 => n2020, B2 => n61713, C1 => n3642, C2 => 
                           n61715, A => n7715, ZN => n7710);
   U6863 : OAI221_X1 port map( B1 => n61697, B2 => n3052, C1 => n53049, C2 => 
                           n61699, A => n7713, ZN => n7712);
   U6864 : NOR4_X1 port map( A1 => n7634, A2 => n7635, A3 => n7636, A4 => n7637
                           , ZN => n7615);
   U6865 : OAI221_X1 port map( B1 => n88, B2 => n61902, C1 => n61899, C2 => 
                           n2721, A => n7639, ZN => n7636);
   U6866 : OAI221_X1 port map( B1 => n2019, B2 => n61713, C1 => n3641, C2 => 
                           n61715, A => n7640, ZN => n7635);
   U6867 : OAI221_X1 port map( B1 => n61697, B2 => n3051, C1 => n53048, C2 => 
                           n61699, A => n7638, ZN => n7637);
   U6868 : NOR4_X1 port map( A1 => n7559, A2 => n7560, A3 => n7561, A4 => n7562
                           , ZN => n7540);
   U6869 : OAI221_X1 port map( B1 => n87, B2 => n61902, C1 => n61899, C2 => 
                           n2720, A => n7564, ZN => n7561);
   U6870 : OAI221_X1 port map( B1 => n2018, B2 => n61713, C1 => n3640, C2 => 
                           n61715, A => n7565, ZN => n7560);
   U6871 : OAI221_X1 port map( B1 => n61697, B2 => n3050, C1 => n53047, C2 => 
                           n61699, A => n7563, ZN => n7562);
   U6872 : NOR4_X1 port map( A1 => n7484, A2 => n7485, A3 => n7486, A4 => n7487
                           , ZN => n7465);
   U6873 : OAI221_X1 port map( B1 => n86, B2 => n61902, C1 => n61899, C2 => 
                           n2719, A => n7489, ZN => n7486);
   U6874 : OAI221_X1 port map( B1 => n2017, B2 => n61713, C1 => n3639, C2 => 
                           n61715, A => n7490, ZN => n7485);
   U6875 : OAI221_X1 port map( B1 => n61697, B2 => n3049, C1 => n53046, C2 => 
                           n61699, A => n7488, ZN => n7487);
   U6876 : NOR4_X1 port map( A1 => n7409, A2 => n7410, A3 => n7411, A4 => n7412
                           , ZN => n7390);
   U6877 : OAI221_X1 port map( B1 => n85, B2 => n61902, C1 => n61899, C2 => 
                           n2718, A => n7414, ZN => n7411);
   U6878 : OAI221_X1 port map( B1 => n2016, B2 => n61713, C1 => n3638, C2 => 
                           n61715, A => n7415, ZN => n7410);
   U6879 : OAI221_X1 port map( B1 => n61697, B2 => n3048, C1 => n53045, C2 => 
                           n61699, A => n7413, ZN => n7412);
   U6880 : NOR4_X1 port map( A1 => n7334, A2 => n7335, A3 => n7336, A4 => n7337
                           , ZN => n7315);
   U6881 : OAI221_X1 port map( B1 => n84, B2 => n61902, C1 => n61898, C2 => 
                           n2717, A => n7339, ZN => n7336);
   U6882 : OAI221_X1 port map( B1 => n2015, B2 => n61713, C1 => n3637, C2 => 
                           n61715, A => n7340, ZN => n7335);
   U6883 : OAI221_X1 port map( B1 => n61697, B2 => n3047, C1 => n53044, C2 => 
                           n61699, A => n7338, ZN => n7337);
   U6884 : NOR4_X1 port map( A1 => n7184, A2 => n7185, A3 => n7186, A4 => n7187
                           , ZN => n7165);
   U6885 : OAI221_X1 port map( B1 => n82, B2 => n61901, C1 => n61898, C2 => 
                           n2715, A => n7189, ZN => n7186);
   U6886 : OAI221_X1 port map( B1 => n2013, B2 => n61713, C1 => n3635, C2 => 
                           n61715, A => n7190, ZN => n7185);
   U6887 : OAI221_X1 port map( B1 => n61697, B2 => n3045, C1 => n53042, C2 => 
                           n61699, A => n7188, ZN => n7187);
   U6888 : NOR4_X1 port map( A1 => n6959, A2 => n6960, A3 => n6961, A4 => n6962
                           , ZN => n6940);
   U6889 : OAI221_X1 port map( B1 => n61900, B2 => n2688, C1 => n61898, C2 => 
                           n2712, A => n6964, ZN => n6961);
   U6890 : OAI221_X1 port map( B1 => n2010, B2 => n6044, C1 => n3632, C2 => 
                           n61716, A => n6965, ZN => n6960);
   U6891 : OAI221_X1 port map( B1 => n6062, B2 => n3042, C1 => n53039, C2 => 
                           n61700, A => n6963, ZN => n6962);
   U6892 : NOR4_X1 port map( A1 => n6037, A2 => n6038, A3 => n6039, A4 => n6040
                           , ZN => n6009);
   U6893 : OAI221_X1 port map( B1 => n61890, B2 => n1005, C1 => n61887, C2 => 
                           n1013, A => n6042, ZN => n6039);
   U6894 : OAI221_X1 port map( B1 => n52743, B2 => n61901, C1 => n52751, C2 => 
                           n61897, A => n6041, ZN => n6040);
   U6895 : OAI221_X1 port map( B1 => n5440, B2 => n4240, C1 => n9754, C2 => 
                           n5441, A => n6046, ZN => n6037);
   U6896 : NOR4_X1 port map( A1 => n5953, A2 => n5954, A3 => n5955, A4 => n5956
                           , ZN => n5934);
   U6897 : OAI221_X1 port map( B1 => n61890, B2 => n1004, C1 => n61887, C2 => 
                           n1012, A => n5958, ZN => n5955);
   U6898 : OAI221_X1 port map( B1 => n52742, B2 => n61901, C1 => n52750, C2 => 
                           n61897, A => n5957, ZN => n5956);
   U6899 : OAI221_X1 port map( B1 => n5440, B2 => n4239, C1 => n9753, C2 => 
                           n5441, A => n5960, ZN => n5953);
   U6900 : NOR4_X1 port map( A1 => n5878, A2 => n5879, A3 => n5880, A4 => n5881
                           , ZN => n5859);
   U6901 : OAI221_X1 port map( B1 => n61890, B2 => n1003, C1 => n61887, C2 => 
                           n1011, A => n5883, ZN => n5880);
   U6902 : OAI221_X1 port map( B1 => n52741, B2 => n61901, C1 => n52749, C2 => 
                           n61897, A => n5882, ZN => n5881);
   U6903 : OAI221_X1 port map( B1 => n5440, B2 => n4238, C1 => n9752, C2 => 
                           n5441, A => n5885, ZN => n5878);
   U6904 : NOR4_X1 port map( A1 => n5803, A2 => n5804, A3 => n5805, A4 => n5806
                           , ZN => n5784);
   U6905 : OAI221_X1 port map( B1 => n61890, B2 => n1002, C1 => n61887, C2 => 
                           n1010, A => n5808, ZN => n5805);
   U6906 : OAI221_X1 port map( B1 => n52740, B2 => n61901, C1 => n52748, C2 => 
                           n61897, A => n5807, ZN => n5806);
   U6907 : OAI221_X1 port map( B1 => n5440, B2 => n4237, C1 => n9751, C2 => 
                           n5441, A => n5810, ZN => n5803);
   U6908 : NOR4_X1 port map( A1 => n5728, A2 => n5729, A3 => n5730, A4 => n5731
                           , ZN => n5709);
   U6909 : OAI221_X1 port map( B1 => n61890, B2 => n1001, C1 => n61887, C2 => 
                           n1009, A => n5733, ZN => n5730);
   U6910 : OAI221_X1 port map( B1 => n52739, B2 => n61901, C1 => n52747, C2 => 
                           n61897, A => n5732, ZN => n5731);
   U6911 : OAI221_X1 port map( B1 => n5440, B2 => n4236, C1 => n9750, C2 => 
                           n5441, A => n5735, ZN => n5728);
   U6912 : NOR4_X1 port map( A1 => n5653, A2 => n5654, A3 => n5655, A4 => n5656
                           , ZN => n5634);
   U6913 : OAI221_X1 port map( B1 => n61890, B2 => n1000, C1 => n61887, C2 => 
                           n1008, A => n5658, ZN => n5655);
   U6914 : OAI221_X1 port map( B1 => n52738, B2 => n61901, C1 => n52746, C2 => 
                           n61897, A => n5657, ZN => n5656);
   U6915 : OAI221_X1 port map( B1 => n5440, B2 => n985, C1 => n9749, C2 => 
                           n5441, A => n5660, ZN => n5653);
   U6916 : NOR4_X1 port map( A1 => n5578, A2 => n5579, A3 => n5580, A4 => n5581
                           , ZN => n5559);
   U6917 : OAI221_X1 port map( B1 => n61890, B2 => n995, C1 => n61887, C2 => 
                           n1007, A => n5583, ZN => n5580);
   U6918 : OAI221_X1 port map( B1 => n52737, B2 => n61901, C1 => n52745, C2 => 
                           n61897, A => n5582, ZN => n5581);
   U6919 : OAI221_X1 port map( B1 => n5440, B2 => n984, C1 => n9748, C2 => 
                           n5441, A => n5585, ZN => n5578);
   U6920 : NOR4_X1 port map( A1 => n5423, A2 => n5424, A3 => n5425, A4 => n5426
                           , ZN => n5379);
   U6921 : OAI221_X1 port map( B1 => n61890, B2 => n994, C1 => n61887, C2 => 
                           n1006, A => n5434, ZN => n5425);
   U6922 : OAI221_X1 port map( B1 => n52736, B2 => n61901, C1 => n52744, C2 => 
                           n61897, A => n5429, ZN => n5426);
   U6923 : OAI221_X1 port map( B1 => n5440, B2 => n983, C1 => n9747, C2 => 
                           n5441, A => n5442, ZN => n5423);
   U6924 : NOR4_X1 port map( A1 => n14388, A2 => n14389, A3 => n14390, A4 => 
                           n14391, ZN => n14369);
   U6925 : OAI221_X1 port map( B1 => n3190, B2 => n61538, C1 => n3200, C2 => 
                           n61535, A => n14394, ZN => n14389);
   U6926 : OAI221_X1 port map( B1 => n3224, B2 => n61550, C1 => n3248, C2 => 
                           n61547, A => n14393, ZN => n14390);
   U6927 : OAI221_X1 port map( B1 => n3636, B2 => n61562, C1 => n2014, C2 => 
                           n61559, A => n14392, ZN => n14391);
   U6928 : NOR4_X1 port map( A1 => n14424, A2 => n14425, A3 => n14426, A4 => 
                           n14427, ZN => n14405);
   U6929 : OAI221_X1 port map( B1 => n3564, B2 => n61334, C1 => n3588, C2 => 
                           n61331, A => n14430, ZN => n14425);
   U6930 : OAI221_X1 port map( B1 => n2502, B2 => n61346, C1 => n3982, C2 => 
                           n61343, A => n14429, ZN => n14426);
   U6931 : OAI221_X1 port map( B1 => n3694, B2 => n61358, C1 => n3718, C2 => 
                           n61355, A => n14428, ZN => n14427);
   U6932 : NOR4_X1 port map( A1 => n9897, A2 => n9898, A3 => n9899, A4 => n9900
                           , ZN => n9878);
   U6933 : OAI221_X1 port map( B1 => n3189, B2 => n61538, C1 => n3199, C2 => 
                           n61535, A => n9903, ZN => n9898);
   U6934 : OAI221_X1 port map( B1 => n3223, B2 => n61550, C1 => n3247, C2 => 
                           n61547, A => n9902, ZN => n9899);
   U6935 : OAI221_X1 port map( B1 => n3635, B2 => n61562, C1 => n2013, C2 => 
                           n61559, A => n9901, ZN => n9900);
   U6936 : NOR4_X1 port map( A1 => n14349, A2 => n14350, A3 => n14351, A4 => 
                           n14352, ZN => n9914);
   U6937 : OAI221_X1 port map( B1 => n3563, B2 => n61334, C1 => n3587, C2 => 
                           n61331, A => n14355, ZN => n14350);
   U6938 : OAI221_X1 port map( B1 => n2501, B2 => n61346, C1 => n3981, C2 => 
                           n61343, A => n14354, ZN => n14351);
   U6939 : OAI221_X1 port map( B1 => n3693, B2 => n61358, C1 => n3717, C2 => 
                           n61355, A => n14353, ZN => n14352);
   U6940 : NOR4_X1 port map( A1 => n9822, A2 => n9823, A3 => n9824, A4 => n9825
                           , ZN => n9739);
   U6941 : OAI221_X1 port map( B1 => n3188, B2 => n61538, C1 => n53257, C2 => 
                           n61535, A => n9828, ZN => n9823);
   U6942 : OAI221_X1 port map( B1 => n3222, B2 => n61550, C1 => n3246, C2 => 
                           n61547, A => n9827, ZN => n9824);
   U6943 : OAI221_X1 port map( B1 => n3634, B2 => n61562, C1 => n2012, C2 => 
                           n61559, A => n9826, ZN => n9825);
   U6944 : NOR4_X1 port map( A1 => n9858, A2 => n9859, A3 => n9860, A4 => n9861
                           , ZN => n9839);
   U6945 : OAI221_X1 port map( B1 => n3562, B2 => n61334, C1 => n3586, C2 => 
                           n61331, A => n9864, ZN => n9859);
   U6946 : OAI221_X1 port map( B1 => n2500, B2 => n61346, C1 => n3980, C2 => 
                           n61343, A => n9863, ZN => n9860);
   U6947 : OAI221_X1 port map( B1 => n3692, B2 => n61358, C1 => n3716, C2 => 
                           n61355, A => n9862, ZN => n9861);
   U6948 : NOR4_X1 port map( A1 => n9683, A2 => n9684, A3 => n9685, A4 => n9686
                           , ZN => n9664);
   U6949 : OAI221_X1 port map( B1 => n3187, B2 => n61538, C1 => n53256, C2 => 
                           n61535, A => n9689, ZN => n9684);
   U6950 : OAI221_X1 port map( B1 => n3221, B2 => n61550, C1 => n3245, C2 => 
                           n61547, A => n9688, ZN => n9685);
   U6951 : OAI221_X1 port map( B1 => n3633, B2 => n61562, C1 => n2011, C2 => 
                           n61559, A => n9687, ZN => n9686);
   U6952 : NOR4_X1 port map( A1 => n9719, A2 => n9720, A3 => n9721, A4 => n9722
                           , ZN => n9700);
   U6953 : OAI221_X1 port map( B1 => n3561, B2 => n61334, C1 => n3585, C2 => 
                           n61331, A => n9725, ZN => n9720);
   U6954 : OAI221_X1 port map( B1 => n2499, B2 => n61346, C1 => n3979, C2 => 
                           n61343, A => n9724, ZN => n9721);
   U6955 : OAI221_X1 port map( B1 => n3691, B2 => n61358, C1 => n3715, C2 => 
                           n61355, A => n9723, ZN => n9722);
   U6956 : NOR4_X1 port map( A1 => n9592, A2 => n9593, A3 => n9594, A4 => n9595
                           , ZN => n9573);
   U6957 : OAI221_X1 port map( B1 => n3186, B2 => n61539, C1 => n53255, C2 => 
                           n61536, A => n9598, ZN => n9593);
   U6958 : OAI221_X1 port map( B1 => n3220, B2 => n61551, C1 => n3244, C2 => 
                           n61548, A => n9597, ZN => n9594);
   U6959 : OAI221_X1 port map( B1 => n3632, B2 => n61563, C1 => n2010, C2 => 
                           n61560, A => n9596, ZN => n9595);
   U6960 : NOR4_X1 port map( A1 => n9644, A2 => n9645, A3 => n9646, A4 => n9647
                           , ZN => n9625);
   U6961 : OAI221_X1 port map( B1 => n3560, B2 => n61335, C1 => n3584, C2 => 
                           n61332, A => n9650, ZN => n9645);
   U6962 : OAI221_X1 port map( B1 => n2498, B2 => n61347, C1 => n3978, C2 => 
                           n61344, A => n9649, ZN => n9646);
   U6963 : OAI221_X1 port map( B1 => n3690, B2 => n61359, C1 => n3714, C2 => 
                           n61356, A => n9648, ZN => n9647);
   U6964 : NOR4_X1 port map( A1 => n9517, A2 => n9518, A3 => n9519, A4 => n9520
                           , ZN => n9498);
   U6965 : OAI221_X1 port map( B1 => n3185, B2 => n61539, C1 => n53254, C2 => 
                           n61536, A => n9523, ZN => n9518);
   U6966 : OAI221_X1 port map( B1 => n3219, B2 => n61551, C1 => n3243, C2 => 
                           n61548, A => n9522, ZN => n9519);
   U6967 : OAI221_X1 port map( B1 => n3631, B2 => n61563, C1 => n2009, C2 => 
                           n61560, A => n9521, ZN => n9520);
   U6968 : NOR4_X1 port map( A1 => n9553, A2 => n9554, A3 => n9555, A4 => n9556
                           , ZN => n9534);
   U6969 : OAI221_X1 port map( B1 => n3559, B2 => n61335, C1 => n3583, C2 => 
                           n61332, A => n9559, ZN => n9554);
   U6970 : OAI221_X1 port map( B1 => n2497, B2 => n61347, C1 => n3977, C2 => 
                           n61344, A => n9558, ZN => n9555);
   U6971 : OAI221_X1 port map( B1 => n3689, B2 => n61359, C1 => n3713, C2 => 
                           n61356, A => n9557, ZN => n9556);
   U6972 : NOR4_X1 port map( A1 => n9442, A2 => n9443, A3 => n9444, A4 => n9445
                           , ZN => n9423);
   U6973 : OAI221_X1 port map( B1 => n3184, B2 => n61539, C1 => n53253, C2 => 
                           n61536, A => n9448, ZN => n9443);
   U6974 : OAI221_X1 port map( B1 => n3218, B2 => n61551, C1 => n3242, C2 => 
                           n61548, A => n9447, ZN => n9444);
   U6975 : OAI221_X1 port map( B1 => n3630, B2 => n61563, C1 => n2008, C2 => 
                           n61560, A => n9446, ZN => n9445);
   U6976 : NOR4_X1 port map( A1 => n9478, A2 => n9479, A3 => n9480, A4 => n9481
                           , ZN => n9459);
   U6977 : OAI221_X1 port map( B1 => n3558, B2 => n61335, C1 => n3582, C2 => 
                           n61332, A => n9484, ZN => n9479);
   U6978 : OAI221_X1 port map( B1 => n2496, B2 => n61347, C1 => n3976, C2 => 
                           n61344, A => n9483, ZN => n9480);
   U6979 : OAI221_X1 port map( B1 => n3688, B2 => n61359, C1 => n3712, C2 => 
                           n61356, A => n9482, ZN => n9481);
   U6980 : NOR4_X1 port map( A1 => n9367, A2 => n9368, A3 => n9369, A4 => n9370
                           , ZN => n9348);
   U6981 : OAI221_X1 port map( B1 => n3183, B2 => n61539, C1 => n53252, C2 => 
                           n61536, A => n9373, ZN => n9368);
   U6982 : OAI221_X1 port map( B1 => n3217, B2 => n61551, C1 => n3241, C2 => 
                           n61548, A => n9372, ZN => n9369);
   U6983 : OAI221_X1 port map( B1 => n3629, B2 => n61563, C1 => n2007, C2 => 
                           n61560, A => n9371, ZN => n9370);
   U6984 : NOR4_X1 port map( A1 => n9403, A2 => n9404, A3 => n9405, A4 => n9406
                           , ZN => n9384);
   U6985 : OAI221_X1 port map( B1 => n3557, B2 => n61335, C1 => n3581, C2 => 
                           n61332, A => n9409, ZN => n9404);
   U6986 : OAI221_X1 port map( B1 => n2495, B2 => n61347, C1 => n3975, C2 => 
                           n61344, A => n9408, ZN => n9405);
   U6987 : OAI221_X1 port map( B1 => n3687, B2 => n61359, C1 => n3711, C2 => 
                           n61356, A => n9407, ZN => n9406);
   U6988 : NOR4_X1 port map( A1 => n9228, A2 => n9229, A3 => n9230, A4 => n9231
                           , ZN => n9209);
   U6989 : OAI221_X1 port map( B1 => n3182, B2 => n61539, C1 => n53251, C2 => 
                           n61536, A => n9234, ZN => n9229);
   U6990 : OAI221_X1 port map( B1 => n3216, B2 => n61551, C1 => n3240, C2 => 
                           n61548, A => n9233, ZN => n9230);
   U6991 : OAI221_X1 port map( B1 => n3628, B2 => n61563, C1 => n2006, C2 => 
                           n61560, A => n9232, ZN => n9231);
   U6992 : NOR4_X1 port map( A1 => n9264, A2 => n9265, A3 => n9266, A4 => n9267
                           , ZN => n9245);
   U6993 : OAI221_X1 port map( B1 => n3556, B2 => n61335, C1 => n3580, C2 => 
                           n61332, A => n9270, ZN => n9265);
   U6994 : OAI221_X1 port map( B1 => n2494, B2 => n61347, C1 => n3974, C2 => 
                           n61344, A => n9269, ZN => n9266);
   U6995 : OAI221_X1 port map( B1 => n3686, B2 => n61359, C1 => n3710, C2 => 
                           n61356, A => n9268, ZN => n9267);
   U6996 : NOR4_X1 port map( A1 => n9153, A2 => n9154, A3 => n9155, A4 => n9156
                           , ZN => n9134);
   U6997 : OAI221_X1 port map( B1 => n3181, B2 => n61539, C1 => n53250, C2 => 
                           n61536, A => n9159, ZN => n9154);
   U6998 : OAI221_X1 port map( B1 => n3215, B2 => n61551, C1 => n3239, C2 => 
                           n61548, A => n9158, ZN => n9155);
   U6999 : OAI221_X1 port map( B1 => n3627, B2 => n61563, C1 => n2005, C2 => 
                           n61560, A => n9157, ZN => n9156);
   U7000 : NOR4_X1 port map( A1 => n9189, A2 => n9190, A3 => n9191, A4 => n9192
                           , ZN => n9170);
   U7001 : OAI221_X1 port map( B1 => n3555, B2 => n61335, C1 => n3579, C2 => 
                           n61332, A => n9195, ZN => n9190);
   U7002 : OAI221_X1 port map( B1 => n2493, B2 => n61347, C1 => n3973, C2 => 
                           n61344, A => n9194, ZN => n9191);
   U7003 : OAI221_X1 port map( B1 => n3685, B2 => n61359, C1 => n3709, C2 => 
                           n61356, A => n9193, ZN => n9192);
   U7004 : NOR4_X1 port map( A1 => n9078, A2 => n9079, A3 => n9080, A4 => n9081
                           , ZN => n9059);
   U7005 : OAI221_X1 port map( B1 => n3180, B2 => n61539, C1 => n53249, C2 => 
                           n61536, A => n9084, ZN => n9079);
   U7006 : OAI221_X1 port map( B1 => n3214, B2 => n61551, C1 => n3238, C2 => 
                           n61548, A => n9083, ZN => n9080);
   U7007 : OAI221_X1 port map( B1 => n3626, B2 => n61563, C1 => n2004, C2 => 
                           n61560, A => n9082, ZN => n9081);
   U7008 : NOR4_X1 port map( A1 => n9114, A2 => n9115, A3 => n9116, A4 => n9117
                           , ZN => n9095);
   U7009 : OAI221_X1 port map( B1 => n3554, B2 => n61335, C1 => n3578, C2 => 
                           n61332, A => n9120, ZN => n9115);
   U7010 : OAI221_X1 port map( B1 => n2492, B2 => n61347, C1 => n3972, C2 => 
                           n61344, A => n9119, ZN => n9116);
   U7011 : OAI221_X1 port map( B1 => n3684, B2 => n61359, C1 => n3708, C2 => 
                           n61356, A => n9118, ZN => n9117);
   U7012 : NOR4_X1 port map( A1 => n9003, A2 => n9004, A3 => n9005, A4 => n9006
                           , ZN => n8984);
   U7013 : OAI221_X1 port map( B1 => n3179, B2 => n61539, C1 => n53248, C2 => 
                           n61536, A => n9009, ZN => n9004);
   U7014 : OAI221_X1 port map( B1 => n3213, B2 => n61551, C1 => n3237, C2 => 
                           n61548, A => n9008, ZN => n9005);
   U7015 : OAI221_X1 port map( B1 => n3625, B2 => n61563, C1 => n2003, C2 => 
                           n61560, A => n9007, ZN => n9006);
   U7016 : NOR4_X1 port map( A1 => n9039, A2 => n9040, A3 => n9041, A4 => n9042
                           , ZN => n9020);
   U7017 : OAI221_X1 port map( B1 => n3553, B2 => n61335, C1 => n3577, C2 => 
                           n61332, A => n9045, ZN => n9040);
   U7018 : OAI221_X1 port map( B1 => n2491, B2 => n61347, C1 => n3971, C2 => 
                           n61344, A => n9044, ZN => n9041);
   U7019 : OAI221_X1 port map( B1 => n3683, B2 => n61359, C1 => n3707, C2 => 
                           n61356, A => n9043, ZN => n9042);
   U7020 : NOR4_X1 port map( A1 => n8928, A2 => n8929, A3 => n8930, A4 => n8931
                           , ZN => n8909);
   U7021 : OAI221_X1 port map( B1 => n3178, B2 => n61539, C1 => n53247, C2 => 
                           n61536, A => n8934, ZN => n8929);
   U7022 : OAI221_X1 port map( B1 => n3212, B2 => n61551, C1 => n3236, C2 => 
                           n61548, A => n8933, ZN => n8930);
   U7023 : OAI221_X1 port map( B1 => n3624, B2 => n61563, C1 => n2002, C2 => 
                           n61560, A => n8932, ZN => n8931);
   U7024 : NOR4_X1 port map( A1 => n8964, A2 => n8965, A3 => n8966, A4 => n8967
                           , ZN => n8945);
   U7025 : OAI221_X1 port map( B1 => n3552, B2 => n61335, C1 => n3576, C2 => 
                           n61332, A => n8970, ZN => n8965);
   U7026 : OAI221_X1 port map( B1 => n2490, B2 => n61347, C1 => n3970, C2 => 
                           n61344, A => n8969, ZN => n8966);
   U7027 : OAI221_X1 port map( B1 => n3682, B2 => n61359, C1 => n3706, C2 => 
                           n61356, A => n8968, ZN => n8967);
   U7028 : NOR4_X1 port map( A1 => n8853, A2 => n8854, A3 => n8855, A4 => n8856
                           , ZN => n8834);
   U7029 : OAI221_X1 port map( B1 => n3177, B2 => n61539, C1 => n53246, C2 => 
                           n61536, A => n8859, ZN => n8854);
   U7030 : OAI221_X1 port map( B1 => n3211, B2 => n61551, C1 => n3235, C2 => 
                           n61548, A => n8858, ZN => n8855);
   U7031 : OAI221_X1 port map( B1 => n3623, B2 => n61563, C1 => n2001, C2 => 
                           n61560, A => n8857, ZN => n8856);
   U7032 : NOR4_X1 port map( A1 => n8889, A2 => n8890, A3 => n8891, A4 => n8892
                           , ZN => n8870);
   U7033 : OAI221_X1 port map( B1 => n3551, B2 => n61335, C1 => n3575, C2 => 
                           n61332, A => n8895, ZN => n8890);
   U7034 : OAI221_X1 port map( B1 => n2489, B2 => n61347, C1 => n3969, C2 => 
                           n61344, A => n8894, ZN => n8891);
   U7035 : OAI221_X1 port map( B1 => n3681, B2 => n61359, C1 => n3705, C2 => 
                           n61356, A => n8893, ZN => n8892);
   U7036 : NOR4_X1 port map( A1 => n8778, A2 => n8779, A3 => n8780, A4 => n8781
                           , ZN => n8759);
   U7037 : OAI221_X1 port map( B1 => n3176, B2 => n61539, C1 => n53245, C2 => 
                           n61536, A => n8784, ZN => n8779);
   U7038 : OAI221_X1 port map( B1 => n3210, B2 => n61551, C1 => n3234, C2 => 
                           n61548, A => n8783, ZN => n8780);
   U7039 : OAI221_X1 port map( B1 => n3622, B2 => n61563, C1 => n2000, C2 => 
                           n61560, A => n8782, ZN => n8781);
   U7040 : NOR4_X1 port map( A1 => n8814, A2 => n8815, A3 => n8816, A4 => n8817
                           , ZN => n8795);
   U7041 : OAI221_X1 port map( B1 => n3550, B2 => n61335, C1 => n3574, C2 => 
                           n61332, A => n8820, ZN => n8815);
   U7042 : OAI221_X1 port map( B1 => n2488, B2 => n61347, C1 => n3968, C2 => 
                           n61344, A => n8819, ZN => n8816);
   U7043 : OAI221_X1 port map( B1 => n3680, B2 => n61359, C1 => n3704, C2 => 
                           n61356, A => n8818, ZN => n8817);
   U7044 : NOR4_X1 port map( A1 => n8703, A2 => n8704, A3 => n8705, A4 => n8706
                           , ZN => n8684);
   U7045 : OAI221_X1 port map( B1 => n3175, B2 => n61539, C1 => n53244, C2 => 
                           n61536, A => n8709, ZN => n8704);
   U7046 : OAI221_X1 port map( B1 => n3209, B2 => n61551, C1 => n3233, C2 => 
                           n61548, A => n8708, ZN => n8705);
   U7047 : OAI221_X1 port map( B1 => n3621, B2 => n61563, C1 => n1999, C2 => 
                           n61560, A => n8707, ZN => n8706);
   U7048 : NOR4_X1 port map( A1 => n8739, A2 => n8740, A3 => n8741, A4 => n8742
                           , ZN => n8720);
   U7049 : OAI221_X1 port map( B1 => n3549, B2 => n61335, C1 => n3573, C2 => 
                           n61332, A => n8745, ZN => n8740);
   U7050 : OAI221_X1 port map( B1 => n2487, B2 => n61347, C1 => n3967, C2 => 
                           n61344, A => n8744, ZN => n8741);
   U7051 : OAI221_X1 port map( B1 => n3679, B2 => n61359, C1 => n3703, C2 => 
                           n61356, A => n8743, ZN => n8742);
   U7052 : NOR4_X1 port map( A1 => n15006, A2 => n15007, A3 => n15008, A4 => 
                           n15009, ZN => n14969);
   U7053 : OAI221_X1 port map( B1 => n3198, B2 => n61538, C1 => n3208, C2 => 
                           n61535, A => n15014, ZN => n15007);
   U7054 : OAI221_X1 port map( B1 => n3232, B2 => n61550, C1 => n3256, C2 => 
                           n61547, A => n15011, ZN => n15008);
   U7055 : OAI221_X1 port map( B1 => n3644, B2 => n61562, C1 => n2022, C2 => 
                           n61559, A => n15010, ZN => n15009);
   U7056 : NOR4_X1 port map( A1 => n15052, A2 => n15053, A3 => n15054, A4 => 
                           n15055, ZN => n15028);
   U7057 : OAI221_X1 port map( B1 => n3572, B2 => n61334, C1 => n3596, C2 => 
                           n61331, A => n15060, ZN => n15053);
   U7058 : OAI221_X1 port map( B1 => n2510, B2 => n61346, C1 => n3990, C2 => 
                           n61343, A => n15059, ZN => n15054);
   U7059 : OAI221_X1 port map( B1 => n3702, B2 => n61358, C1 => n3726, C2 => 
                           n61355, A => n15056, ZN => n15055);
   U7060 : NOR4_X1 port map( A1 => n14913, A2 => n14914, A3 => n14915, A4 => 
                           n14916, ZN => n14894);
   U7061 : OAI221_X1 port map( B1 => n3197, B2 => n61538, C1 => n3207, C2 => 
                           n61535, A => n14919, ZN => n14914);
   U7062 : OAI221_X1 port map( B1 => n3231, B2 => n61550, C1 => n3255, C2 => 
                           n61547, A => n14918, ZN => n14915);
   U7063 : OAI221_X1 port map( B1 => n3643, B2 => n61562, C1 => n2021, C2 => 
                           n61559, A => n14917, ZN => n14916);
   U7064 : NOR4_X1 port map( A1 => n14949, A2 => n14950, A3 => n14951, A4 => 
                           n14952, ZN => n14930);
   U7065 : OAI221_X1 port map( B1 => n3571, B2 => n61334, C1 => n3595, C2 => 
                           n61331, A => n14955, ZN => n14950);
   U7066 : OAI221_X1 port map( B1 => n2509, B2 => n61346, C1 => n3989, C2 => 
                           n61343, A => n14954, ZN => n14951);
   U7067 : OAI221_X1 port map( B1 => n3701, B2 => n61358, C1 => n3725, C2 => 
                           n61355, A => n14953, ZN => n14952);
   U7068 : NOR4_X1 port map( A1 => n14838, A2 => n14839, A3 => n14840, A4 => 
                           n14841, ZN => n14819);
   U7069 : OAI221_X1 port map( B1 => n3196, B2 => n61538, C1 => n3206, C2 => 
                           n61535, A => n14844, ZN => n14839);
   U7070 : OAI221_X1 port map( B1 => n3230, B2 => n61550, C1 => n3254, C2 => 
                           n61547, A => n14843, ZN => n14840);
   U7071 : OAI221_X1 port map( B1 => n3642, B2 => n61562, C1 => n2020, C2 => 
                           n61559, A => n14842, ZN => n14841);
   U7072 : NOR4_X1 port map( A1 => n14874, A2 => n14875, A3 => n14876, A4 => 
                           n14877, ZN => n14855);
   U7073 : OAI221_X1 port map( B1 => n3570, B2 => n61334, C1 => n3594, C2 => 
                           n61331, A => n14880, ZN => n14875);
   U7074 : OAI221_X1 port map( B1 => n2508, B2 => n61346, C1 => n3988, C2 => 
                           n61343, A => n14879, ZN => n14876);
   U7075 : OAI221_X1 port map( B1 => n3700, B2 => n61358, C1 => n3724, C2 => 
                           n61355, A => n14878, ZN => n14877);
   U7076 : NOR4_X1 port map( A1 => n14763, A2 => n14764, A3 => n14765, A4 => 
                           n14766, ZN => n14744);
   U7077 : OAI221_X1 port map( B1 => n3195, B2 => n61538, C1 => n3205, C2 => 
                           n61535, A => n14769, ZN => n14764);
   U7078 : OAI221_X1 port map( B1 => n3229, B2 => n61550, C1 => n3253, C2 => 
                           n61547, A => n14768, ZN => n14765);
   U7079 : OAI221_X1 port map( B1 => n3641, B2 => n61562, C1 => n2019, C2 => 
                           n61559, A => n14767, ZN => n14766);
   U7080 : NOR4_X1 port map( A1 => n14799, A2 => n14800, A3 => n14801, A4 => 
                           n14802, ZN => n14780);
   U7081 : OAI221_X1 port map( B1 => n3569, B2 => n61334, C1 => n3593, C2 => 
                           n61331, A => n14805, ZN => n14800);
   U7082 : OAI221_X1 port map( B1 => n2507, B2 => n61346, C1 => n3987, C2 => 
                           n61343, A => n14804, ZN => n14801);
   U7083 : OAI221_X1 port map( B1 => n3699, B2 => n61358, C1 => n3723, C2 => 
                           n61355, A => n14803, ZN => n14802);
   U7084 : NOR4_X1 port map( A1 => n14688, A2 => n14689, A3 => n14690, A4 => 
                           n14691, ZN => n14669);
   U7085 : OAI221_X1 port map( B1 => n3194, B2 => n61538, C1 => n3204, C2 => 
                           n61535, A => n14694, ZN => n14689);
   U7086 : OAI221_X1 port map( B1 => n3228, B2 => n61550, C1 => n3252, C2 => 
                           n61547, A => n14693, ZN => n14690);
   U7087 : OAI221_X1 port map( B1 => n3640, B2 => n61562, C1 => n2018, C2 => 
                           n61559, A => n14692, ZN => n14691);
   U7088 : NOR4_X1 port map( A1 => n14724, A2 => n14725, A3 => n14726, A4 => 
                           n14727, ZN => n14705);
   U7089 : OAI221_X1 port map( B1 => n3568, B2 => n61334, C1 => n3592, C2 => 
                           n61331, A => n14730, ZN => n14725);
   U7090 : OAI221_X1 port map( B1 => n2506, B2 => n61346, C1 => n3986, C2 => 
                           n61343, A => n14729, ZN => n14726);
   U7091 : OAI221_X1 port map( B1 => n3698, B2 => n61358, C1 => n3722, C2 => 
                           n61355, A => n14728, ZN => n14727);
   U7092 : NOR4_X1 port map( A1 => n14613, A2 => n14614, A3 => n14615, A4 => 
                           n14616, ZN => n14594);
   U7093 : OAI221_X1 port map( B1 => n3193, B2 => n61538, C1 => n3203, C2 => 
                           n61535, A => n14619, ZN => n14614);
   U7094 : OAI221_X1 port map( B1 => n3227, B2 => n61550, C1 => n3251, C2 => 
                           n61547, A => n14618, ZN => n14615);
   U7095 : OAI221_X1 port map( B1 => n3639, B2 => n61562, C1 => n2017, C2 => 
                           n61559, A => n14617, ZN => n14616);
   U7096 : NOR4_X1 port map( A1 => n14649, A2 => n14650, A3 => n14651, A4 => 
                           n14652, ZN => n14630);
   U7097 : OAI221_X1 port map( B1 => n3567, B2 => n61334, C1 => n3591, C2 => 
                           n61331, A => n14655, ZN => n14650);
   U7098 : OAI221_X1 port map( B1 => n2505, B2 => n61346, C1 => n3985, C2 => 
                           n61343, A => n14654, ZN => n14651);
   U7099 : OAI221_X1 port map( B1 => n3697, B2 => n61358, C1 => n3721, C2 => 
                           n61355, A => n14653, ZN => n14652);
   U7100 : NOR4_X1 port map( A1 => n14538, A2 => n14539, A3 => n14540, A4 => 
                           n14541, ZN => n14519);
   U7101 : OAI221_X1 port map( B1 => n3192, B2 => n61538, C1 => n3202, C2 => 
                           n61535, A => n14544, ZN => n14539);
   U7102 : OAI221_X1 port map( B1 => n3226, B2 => n61550, C1 => n3250, C2 => 
                           n61547, A => n14543, ZN => n14540);
   U7103 : OAI221_X1 port map( B1 => n3638, B2 => n61562, C1 => n2016, C2 => 
                           n61559, A => n14542, ZN => n14541);
   U7104 : NOR4_X1 port map( A1 => n14574, A2 => n14575, A3 => n14576, A4 => 
                           n14577, ZN => n14555);
   U7105 : OAI221_X1 port map( B1 => n3566, B2 => n61334, C1 => n3590, C2 => 
                           n61331, A => n14580, ZN => n14575);
   U7106 : OAI221_X1 port map( B1 => n2504, B2 => n61346, C1 => n3984, C2 => 
                           n61343, A => n14579, ZN => n14576);
   U7107 : OAI221_X1 port map( B1 => n3696, B2 => n61358, C1 => n3720, C2 => 
                           n61355, A => n14578, ZN => n14577);
   U7108 : NOR4_X1 port map( A1 => n14463, A2 => n14464, A3 => n14465, A4 => 
                           n14466, ZN => n14444);
   U7109 : OAI221_X1 port map( B1 => n3191, B2 => n61538, C1 => n3201, C2 => 
                           n61535, A => n14469, ZN => n14464);
   U7110 : OAI221_X1 port map( B1 => n3225, B2 => n61550, C1 => n3249, C2 => 
                           n61547, A => n14468, ZN => n14465);
   U7111 : OAI221_X1 port map( B1 => n3637, B2 => n61562, C1 => n2015, C2 => 
                           n61559, A => n14467, ZN => n14466);
   U7112 : NOR4_X1 port map( A1 => n14499, A2 => n14500, A3 => n14501, A4 => 
                           n14502, ZN => n14480);
   U7113 : OAI221_X1 port map( B1 => n3565, B2 => n61334, C1 => n3589, C2 => 
                           n61331, A => n14505, ZN => n14500);
   U7114 : OAI221_X1 port map( B1 => n2503, B2 => n61346, C1 => n3983, C2 => 
                           n61343, A => n14504, ZN => n14501);
   U7115 : OAI221_X1 port map( B1 => n3695, B2 => n61358, C1 => n3719, C2 => 
                           n61355, A => n14503, ZN => n14502);
   U7116 : NOR4_X1 port map( A1 => n6742, A2 => n6743, A3 => n6744, A4 => n6745
                           , ZN => n6714);
   U7117 : OAI221_X1 port map( B1 => n53252, B2 => n6048, C1 => n61711, C2 => 
                           n3135, A => n6747, ZN => n6744);
   U7118 : OAI221_X1 port map( B1 => n6056, B2 => n2883, C1 => n61708, C2 => 
                           n2943, A => n6748, ZN => n6743);
   U7119 : OAI221_X1 port map( B1 => n61945, B2 => n2757, C1 => n53582, C2 => 
                           n61949, A => n6746, ZN => n6745);
   U7120 : NOR4_X1 port map( A1 => n6667, A2 => n6668, A3 => n6669, A4 => n6670
                           , ZN => n6639);
   U7121 : OAI221_X1 port map( B1 => n53251, B2 => n6048, C1 => n6047, C2 => 
                           n3134, A => n6672, ZN => n6669);
   U7122 : OAI221_X1 port map( B1 => n6056, B2 => n2882, C1 => n61708, C2 => 
                           n2942, A => n6673, ZN => n6668);
   U7123 : OAI221_X1 port map( B1 => n61945, B2 => n2756, C1 => n53581, C2 => 
                           n61949, A => n6671, ZN => n6670);
   U7124 : NOR4_X1 port map( A1 => n6592, A2 => n6593, A3 => n6594, A4 => n6595
                           , ZN => n6564);
   U7125 : OAI221_X1 port map( B1 => n53250, B2 => n6048, C1 => n6047, C2 => 
                           n3133, A => n6597, ZN => n6594);
   U7126 : OAI221_X1 port map( B1 => n6056, B2 => n2881, C1 => n61708, C2 => 
                           n2941, A => n6598, ZN => n6593);
   U7127 : OAI221_X1 port map( B1 => n61945, B2 => n2755, C1 => n53580, C2 => 
                           n61949, A => n6596, ZN => n6595);
   U7128 : NOR4_X1 port map( A1 => n6517, A2 => n6518, A3 => n6519, A4 => n6520
                           , ZN => n6489);
   U7129 : OAI221_X1 port map( B1 => n53249, B2 => n6048, C1 => n6047, C2 => 
                           n3132, A => n6522, ZN => n6519);
   U7130 : OAI221_X1 port map( B1 => n6056, B2 => n2880, C1 => n61708, C2 => 
                           n2940, A => n6523, ZN => n6518);
   U7131 : OAI221_X1 port map( B1 => n61945, B2 => n2754, C1 => n53579, C2 => 
                           n61949, A => n6521, ZN => n6520);
   U7132 : NOR4_X1 port map( A1 => n6442, A2 => n6443, A3 => n6444, A4 => n6445
                           , ZN => n6414);
   U7133 : OAI221_X1 port map( B1 => n53248, B2 => n6048, C1 => n6047, C2 => 
                           n3131, A => n6447, ZN => n6444);
   U7134 : OAI221_X1 port map( B1 => n6056, B2 => n2879, C1 => n61708, C2 => 
                           n2939, A => n6448, ZN => n6443);
   U7135 : OAI221_X1 port map( B1 => n61945, B2 => n2753, C1 => n53578, C2 => 
                           n61949, A => n6446, ZN => n6445);
   U7136 : NOR4_X1 port map( A1 => n6367, A2 => n6368, A3 => n6369, A4 => n6370
                           , ZN => n6339);
   U7137 : OAI221_X1 port map( B1 => n53247, B2 => n6048, C1 => n6047, C2 => 
                           n3130, A => n6372, ZN => n6369);
   U7138 : OAI221_X1 port map( B1 => n6056, B2 => n2878, C1 => n61708, C2 => 
                           n2938, A => n6373, ZN => n6368);
   U7139 : OAI221_X1 port map( B1 => n61945, B2 => n2752, C1 => n53577, C2 => 
                           n61948, A => n6371, ZN => n6370);
   U7140 : NOR4_X1 port map( A1 => n6292, A2 => n6293, A3 => n6294, A4 => n6295
                           , ZN => n6264);
   U7141 : OAI221_X1 port map( B1 => n53246, B2 => n6048, C1 => n6047, C2 => 
                           n3129, A => n6297, ZN => n6294);
   U7142 : OAI221_X1 port map( B1 => n6056, B2 => n2877, C1 => n61708, C2 => 
                           n2937, A => n6298, ZN => n6293);
   U7143 : OAI221_X1 port map( B1 => n61945, B2 => n2751, C1 => n53576, C2 => 
                           n61948, A => n6296, ZN => n6295);
   U7144 : NOR4_X1 port map( A1 => n6217, A2 => n6218, A3 => n6219, A4 => n6220
                           , ZN => n6189);
   U7145 : OAI221_X1 port map( B1 => n53245, B2 => n6048, C1 => n6047, C2 => 
                           n3128, A => n6222, ZN => n6219);
   U7146 : OAI221_X1 port map( B1 => n6056, B2 => n2876, C1 => n61708, C2 => 
                           n2936, A => n6223, ZN => n6218);
   U7147 : OAI221_X1 port map( B1 => n957, B2 => n61949, C1 => n61946, C2 => 
                           n2750, A => n6221, ZN => n6220);
   U7148 : NOR4_X1 port map( A1 => n6142, A2 => n6143, A3 => n6144, A4 => n6145
                           , ZN => n6114);
   U7149 : OAI221_X1 port map( B1 => n53244, B2 => n6048, C1 => n6047, C2 => 
                           n3127, A => n6147, ZN => n6144);
   U7150 : OAI221_X1 port map( B1 => n6056, B2 => n2875, C1 => n61708, C2 => 
                           n2935, A => n6148, ZN => n6143);
   U7151 : OAI221_X1 port map( B1 => n61945, B2 => n2749, C1 => n53575, C2 => 
                           n61948, A => n6146, ZN => n6145);
   U7152 : NOR4_X1 port map( A1 => n7117, A2 => n7118, A3 => n7119, A4 => n7120
                           , ZN => n7089);
   U7153 : OAI221_X1 port map( B1 => n53257, B2 => n61709, C1 => n61711, C2 => 
                           n3140, A => n7122, ZN => n7119);
   U7154 : OAI221_X1 port map( B1 => n61705, B2 => n2908, C1 => n61707, C2 => 
                           n2948, A => n7123, ZN => n7118);
   U7155 : OAI221_X1 port map( B1 => n961, B2 => n61949, C1 => n61946, C2 => 
                           n2762, A => n7121, ZN => n7120);
   U7156 : NOR4_X1 port map( A1 => n7042, A2 => n7043, A3 => n7044, A4 => n7045
                           , ZN => n7014);
   U7157 : OAI221_X1 port map( B1 => n53256, B2 => n61709, C1 => n61711, C2 => 
                           n3139, A => n7047, ZN => n7044);
   U7158 : OAI221_X1 port map( B1 => n61705, B2 => n2907, C1 => n61707, C2 => 
                           n2947, A => n7048, ZN => n7043);
   U7159 : OAI221_X1 port map( B1 => n960, B2 => n61949, C1 => n61946, C2 => 
                           n2761, A => n7046, ZN => n7045);
   U7160 : NOR4_X1 port map( A1 => n6892, A2 => n6893, A3 => n6894, A4 => n6895
                           , ZN => n6864);
   U7161 : OAI221_X1 port map( B1 => n53254, B2 => n6048, C1 => n6047, C2 => 
                           n3137, A => n6897, ZN => n6894);
   U7162 : OAI221_X1 port map( B1 => n6056, B2 => n2885, C1 => n61708, C2 => 
                           n2945, A => n6898, ZN => n6893);
   U7163 : OAI221_X1 port map( B1 => n958, B2 => n61949, C1 => n61946, C2 => 
                           n2759, A => n6896, ZN => n6895);
   U7164 : NOR4_X1 port map( A1 => n6817, A2 => n6818, A3 => n6819, A4 => n6820
                           , ZN => n6789);
   U7165 : OAI221_X1 port map( B1 => n53253, B2 => n6048, C1 => n6047, C2 => 
                           n3136, A => n6822, ZN => n6819);
   U7166 : OAI221_X1 port map( B1 => n6056, B2 => n2884, C1 => n61708, C2 => 
                           n2944, A => n6823, ZN => n6818);
   U7167 : OAI221_X1 port map( B1 => n61945, B2 => n2758, C1 => n53583, C2 => 
                           n61949, A => n6821, ZN => n6820);
   U7168 : NOR4_X1 port map( A1 => n7891, A2 => n7892, A3 => n7893, A4 => n7894
                           , ZN => n7839);
   U7169 : OAI221_X1 port map( B1 => n61709, B2 => n3208, C1 => n61711, C2 => 
                           n3150, A => n7897, ZN => n7893);
   U7170 : OAI221_X1 port map( B1 => n61705, B2 => n2934, C1 => n61707, C2 => 
                           n2958, A => n7898, ZN => n7892);
   U7171 : OAI221_X1 port map( B1 => n61948, B2 => n2778, C1 => n53574, C2 => 
                           n61945, A => n7895, ZN => n7894);
   U7172 : NOR4_X1 port map( A1 => n7792, A2 => n7793, A3 => n7794, A4 => n7795
                           , ZN => n7764);
   U7173 : OAI221_X1 port map( B1 => n61709, B2 => n3207, C1 => n61711, C2 => 
                           n3149, A => n7797, ZN => n7794);
   U7174 : OAI221_X1 port map( B1 => n61705, B2 => n2933, C1 => n61707, C2 => 
                           n2957, A => n7798, ZN => n7793);
   U7175 : OAI221_X1 port map( B1 => n61948, B2 => n2777, C1 => n53573, C2 => 
                           n61946, A => n7796, ZN => n7795);
   U7176 : NOR4_X1 port map( A1 => n7717, A2 => n7718, A3 => n7719, A4 => n7720
                           , ZN => n7689);
   U7177 : OAI221_X1 port map( B1 => n61709, B2 => n3206, C1 => n61711, C2 => 
                           n3148, A => n7722, ZN => n7719);
   U7178 : OAI221_X1 port map( B1 => n61705, B2 => n2932, C1 => n61707, C2 => 
                           n2956, A => n7723, ZN => n7718);
   U7179 : OAI221_X1 port map( B1 => n61948, B2 => n2776, C1 => n53572, C2 => 
                           n61946, A => n7721, ZN => n7720);
   U7180 : NOR4_X1 port map( A1 => n7192, A2 => n7193, A3 => n7194, A4 => n7195
                           , ZN => n7164);
   U7181 : OAI221_X1 port map( B1 => n61709, B2 => n3199, C1 => n61711, C2 => 
                           n3141, A => n7197, ZN => n7194);
   U7182 : OAI221_X1 port map( B1 => n61705, B2 => n2925, C1 => n61707, C2 => 
                           n2949, A => n7198, ZN => n7193);
   U7183 : OAI221_X1 port map( B1 => n962, B2 => n61950, C1 => n61946, C2 => 
                           n2763, A => n7196, ZN => n7195);
   U7184 : NOR4_X1 port map( A1 => n6967, A2 => n6968, A3 => n6969, A4 => n6970
                           , ZN => n6939);
   U7185 : OAI221_X1 port map( B1 => n53255, B2 => n6048, C1 => n6047, C2 => 
                           n3138, A => n6972, ZN => n6969);
   U7186 : OAI221_X1 port map( B1 => n6056, B2 => n2886, C1 => n61708, C2 => 
                           n2946, A => n6973, ZN => n6968);
   U7187 : OAI221_X1 port map( B1 => n959, B2 => n61949, C1 => n61947, C2 => 
                           n2760, A => n6971, ZN => n6970);
   U7188 : NOR4_X1 port map( A1 => n6049, A2 => n6050, A3 => n6051, A4 => n6052
                           , ZN => n6008);
   U7189 : OAI221_X1 port map( B1 => n5456, B2 => n794, C1 => n5457, C2 => n802
                           , A => n6057, ZN => n6050);
   U7190 : OAI221_X1 port map( B1 => n546, B2 => n5453, C1 => n5454, C2 => 
                           n4219, A => n6054, ZN => n6051);
   U7191 : OAI221_X1 port map( B1 => n5459, B2 => n562, C1 => n52735, C2 => 
                           n5460, A => n6060, ZN => n6049);
   U7192 : NOR4_X1 port map( A1 => n5961, A2 => n5962, A3 => n5963, A4 => n5964
                           , ZN => n5933);
   U7193 : OAI221_X1 port map( B1 => n5456, B2 => n793, C1 => n5457, C2 => n801
                           , A => n5967, ZN => n5962);
   U7194 : OAI221_X1 port map( B1 => n545, B2 => n5453, C1 => n5454, C2 => 
                           n4218, A => n5966, ZN => n5963);
   U7195 : OAI221_X1 port map( B1 => n5459, B2 => n561, C1 => n52734, C2 => 
                           n5460, A => n5968, ZN => n5961);
   U7196 : NOR4_X1 port map( A1 => n5886, A2 => n5887, A3 => n5888, A4 => n5889
                           , ZN => n5858);
   U7197 : OAI221_X1 port map( B1 => n5456, B2 => n792, C1 => n5457, C2 => n800
                           , A => n5892, ZN => n5887);
   U7198 : OAI221_X1 port map( B1 => n544, B2 => n5453, C1 => n5454, C2 => 
                           n4217, A => n5891, ZN => n5888);
   U7199 : OAI221_X1 port map( B1 => n5459, B2 => n560, C1 => n52733, C2 => 
                           n5460, A => n5893, ZN => n5886);
   U7200 : NOR4_X1 port map( A1 => n5811, A2 => n5812, A3 => n5813, A4 => n5814
                           , ZN => n5783);
   U7201 : OAI221_X1 port map( B1 => n5456, B2 => n791, C1 => n5457, C2 => n799
                           , A => n5817, ZN => n5812);
   U7202 : OAI221_X1 port map( B1 => n543, B2 => n5453, C1 => n5454, C2 => 
                           n4216, A => n5816, ZN => n5813);
   U7203 : OAI221_X1 port map( B1 => n5459, B2 => n499, C1 => n52732, C2 => 
                           n5460, A => n5818, ZN => n5811);
   U7204 : NOR4_X1 port map( A1 => n5736, A2 => n5737, A3 => n5738, A4 => n5739
                           , ZN => n5708);
   U7205 : OAI221_X1 port map( B1 => n5456, B2 => n790, C1 => n5457, C2 => n798
                           , A => n5742, ZN => n5737);
   U7206 : OAI221_X1 port map( B1 => n542, B2 => n5453, C1 => n5454, C2 => 
                           n4215, A => n5741, ZN => n5738);
   U7207 : OAI221_X1 port map( B1 => n5459, B2 => n498, C1 => n52731, C2 => 
                           n5460, A => n5743, ZN => n5736);
   U7208 : NOR4_X1 port map( A1 => n5661, A2 => n5662, A3 => n5663, A4 => n5664
                           , ZN => n5633);
   U7209 : OAI221_X1 port map( B1 => n5456, B2 => n789, C1 => n5457, C2 => n797
                           , A => n5667, ZN => n5662);
   U7210 : OAI221_X1 port map( B1 => n541, B2 => n5453, C1 => n5454, C2 => 
                           n4214, A => n5666, ZN => n5663);
   U7211 : OAI221_X1 port map( B1 => n5459, B2 => n497, C1 => n52730, C2 => 
                           n5460, A => n5668, ZN => n5661);
   U7212 : NOR4_X1 port map( A1 => n5586, A2 => n5587, A3 => n5588, A4 => n5589
                           , ZN => n5558);
   U7213 : OAI221_X1 port map( B1 => n5456, B2 => n788, C1 => n5457, C2 => n796
                           , A => n5592, ZN => n5587);
   U7214 : OAI221_X1 port map( B1 => n540, B2 => n5453, C1 => n5454, C2 => 
                           n4213, A => n5591, ZN => n5588);
   U7215 : OAI221_X1 port map( B1 => n5459, B2 => n496, C1 => n52729, C2 => 
                           n5460, A => n5593, ZN => n5586);
   U7216 : NOR4_X1 port map( A1 => n5444, A2 => n5445, A3 => n5446, A4 => n5447
                           , ZN => n5378);
   U7217 : OAI221_X1 port map( B1 => n5456, B2 => n787, C1 => n5457, C2 => n795
                           , A => n5458, ZN => n5445);
   U7218 : OAI221_X1 port map( B1 => n539, B2 => n5453, C1 => n5454, C2 => 
                           n4212, A => n5455, ZN => n5446);
   U7219 : OAI221_X1 port map( B1 => n5459, B2 => n495, C1 => n52728, C2 => 
                           n5460, A => n5461, ZN => n5444);
   U7220 : NOR4_X1 port map( A1 => n14396, A2 => n14397, A3 => n14398, A4 => 
                           n14399, ZN => n14368);
   U7221 : OAI221_X1 port map( B1 => n1684, B2 => n61475, C1 => n428, C2 => 
                           n61472, A => n14403, ZN => n14396);
   U7222 : OAI221_X1 port map( B1 => n4729, B2 => n61487, C1 => n53043, C2 => 
                           n61484, A => n14402, ZN => n14397);
   U7223 : OAI221_X1 port map( B1 => n2950, B2 => n61499, C1 => n2926, C2 => 
                           n61496, A => n14401, ZN => n14398);
   U7224 : NOR4_X1 port map( A1 => n9905, A2 => n9906, A3 => n9907, A4 => n9908
                           , ZN => n9877);
   U7225 : OAI221_X1 port map( B1 => n1683, B2 => n61475, C1 => n427, C2 => 
                           n61472, A => n9912, ZN => n9905);
   U7226 : OAI221_X1 port map( B1 => n4728, B2 => n61487, C1 => n53042, C2 => 
                           n61484, A => n9911, ZN => n9906);
   U7227 : OAI221_X1 port map( B1 => n2949, B2 => n61499, C1 => n2925, C2 => 
                           n61496, A => n9910, ZN => n9907);
   U7228 : NOR4_X1 port map( A1 => n9830, A2 => n9831, A3 => n9832, A4 => n9833
                           , ZN => n9738);
   U7229 : OAI221_X1 port map( B1 => n1682, B2 => n61475, C1 => n426, C2 => 
                           n61472, A => n9837, ZN => n9830);
   U7230 : OAI221_X1 port map( B1 => n4727, B2 => n61487, C1 => n53041, C2 => 
                           n61484, A => n9836, ZN => n9831);
   U7231 : OAI221_X1 port map( B1 => n2948, B2 => n61499, C1 => n2908, C2 => 
                           n61496, A => n9835, ZN => n9832);
   U7232 : NOR4_X1 port map( A1 => n9691, A2 => n9692, A3 => n9693, A4 => n9694
                           , ZN => n9663);
   U7233 : OAI221_X1 port map( B1 => n1681, B2 => n61475, C1 => n425, C2 => 
                           n61472, A => n9698, ZN => n9691);
   U7234 : OAI221_X1 port map( B1 => n4726, B2 => n61487, C1 => n53040, C2 => 
                           n61484, A => n9697, ZN => n9692);
   U7235 : OAI221_X1 port map( B1 => n2947, B2 => n61499, C1 => n2907, C2 => 
                           n61496, A => n9696, ZN => n9693);
   U7236 : NOR4_X1 port map( A1 => n9600, A2 => n9601, A3 => n9602, A4 => n9619
                           , ZN => n9572);
   U7237 : OAI221_X1 port map( B1 => n1680, B2 => n61476, C1 => n424, C2 => 
                           n61473, A => n9623, ZN => n9600);
   U7238 : OAI221_X1 port map( B1 => n4725, B2 => n61488, C1 => n53039, C2 => 
                           n61485, A => n9622, ZN => n9601);
   U7239 : OAI221_X1 port map( B1 => n2946, B2 => n61500, C1 => n2886, C2 => 
                           n61497, A => n9621, ZN => n9602);
   U7240 : NOR4_X1 port map( A1 => n9525, A2 => n9526, A3 => n9527, A4 => n9528
                           , ZN => n9497);
   U7241 : OAI221_X1 port map( B1 => n1679, B2 => n61476, C1 => n423, C2 => 
                           n61473, A => n9532, ZN => n9525);
   U7242 : OAI221_X1 port map( B1 => n4724, B2 => n61488, C1 => n53038, C2 => 
                           n61485, A => n9531, ZN => n9526);
   U7243 : OAI221_X1 port map( B1 => n2945, B2 => n61500, C1 => n2885, C2 => 
                           n61497, A => n9530, ZN => n9527);
   U7244 : NOR4_X1 port map( A1 => n9450, A2 => n9451, A3 => n9452, A4 => n9453
                           , ZN => n9422);
   U7245 : OAI221_X1 port map( B1 => n1678, B2 => n61476, C1 => n422, C2 => 
                           n61473, A => n9457, ZN => n9450);
   U7246 : OAI221_X1 port map( B1 => n4723, B2 => n61488, C1 => n53037, C2 => 
                           n61485, A => n9456, ZN => n9451);
   U7247 : OAI221_X1 port map( B1 => n2944, B2 => n61500, C1 => n2884, C2 => 
                           n61497, A => n9455, ZN => n9452);
   U7248 : NOR4_X1 port map( A1 => n9375, A2 => n9376, A3 => n9377, A4 => n9378
                           , ZN => n9347);
   U7249 : OAI221_X1 port map( B1 => n1677, B2 => n61476, C1 => n421, C2 => 
                           n61473, A => n9382, ZN => n9375);
   U7250 : OAI221_X1 port map( B1 => n4722, B2 => n61488, C1 => n53036, C2 => 
                           n61485, A => n9381, ZN => n9376);
   U7251 : OAI221_X1 port map( B1 => n2943, B2 => n61500, C1 => n2883, C2 => 
                           n61497, A => n9380, ZN => n9377);
   U7252 : NOR4_X1 port map( A1 => n9236, A2 => n9237, A3 => n9238, A4 => n9239
                           , ZN => n9208);
   U7253 : OAI221_X1 port map( B1 => n1676, B2 => n61476, C1 => n420, C2 => 
                           n61473, A => n9243, ZN => n9236);
   U7254 : OAI221_X1 port map( B1 => n4721, B2 => n61488, C1 => n53035, C2 => 
                           n61485, A => n9242, ZN => n9237);
   U7255 : OAI221_X1 port map( B1 => n2942, B2 => n61500, C1 => n2882, C2 => 
                           n61497, A => n9241, ZN => n9238);
   U7256 : NOR4_X1 port map( A1 => n9161, A2 => n9162, A3 => n9163, A4 => n9164
                           , ZN => n9133);
   U7257 : OAI221_X1 port map( B1 => n1675, B2 => n61476, C1 => n419, C2 => 
                           n61473, A => n9168, ZN => n9161);
   U7258 : OAI221_X1 port map( B1 => n4720, B2 => n61488, C1 => n53034, C2 => 
                           n61485, A => n9167, ZN => n9162);
   U7259 : OAI221_X1 port map( B1 => n2941, B2 => n61500, C1 => n2881, C2 => 
                           n61497, A => n9166, ZN => n9163);
   U7260 : NOR4_X1 port map( A1 => n9086, A2 => n9087, A3 => n9088, A4 => n9089
                           , ZN => n9058);
   U7261 : OAI221_X1 port map( B1 => n1674, B2 => n61476, C1 => n418, C2 => 
                           n61473, A => n9093, ZN => n9086);
   U7262 : OAI221_X1 port map( B1 => n4719, B2 => n61488, C1 => n53033, C2 => 
                           n61485, A => n9092, ZN => n9087);
   U7263 : OAI221_X1 port map( B1 => n2940, B2 => n61500, C1 => n2880, C2 => 
                           n61497, A => n9091, ZN => n9088);
   U7264 : NOR4_X1 port map( A1 => n9011, A2 => n9012, A3 => n9013, A4 => n9014
                           , ZN => n8983);
   U7265 : OAI221_X1 port map( B1 => n1673, B2 => n61476, C1 => n417, C2 => 
                           n61473, A => n9018, ZN => n9011);
   U7266 : OAI221_X1 port map( B1 => n4718, B2 => n61488, C1 => n53032, C2 => 
                           n61485, A => n9017, ZN => n9012);
   U7267 : OAI221_X1 port map( B1 => n2939, B2 => n61500, C1 => n2879, C2 => 
                           n61497, A => n9016, ZN => n9013);
   U7268 : NOR4_X1 port map( A1 => n8936, A2 => n8937, A3 => n8938, A4 => n8939
                           , ZN => n8908);
   U7269 : OAI221_X1 port map( B1 => n1672, B2 => n61476, C1 => n416, C2 => 
                           n61473, A => n8943, ZN => n8936);
   U7270 : OAI221_X1 port map( B1 => n4717, B2 => n61488, C1 => n53031, C2 => 
                           n61485, A => n8942, ZN => n8937);
   U7271 : OAI221_X1 port map( B1 => n2938, B2 => n61500, C1 => n2878, C2 => 
                           n61497, A => n8941, ZN => n8938);
   U7272 : NOR4_X1 port map( A1 => n8861, A2 => n8862, A3 => n8863, A4 => n8864
                           , ZN => n8833);
   U7273 : OAI221_X1 port map( B1 => n1671, B2 => n61476, C1 => n415, C2 => 
                           n61473, A => n8868, ZN => n8861);
   U7274 : OAI221_X1 port map( B1 => n4716, B2 => n61488, C1 => n53030, C2 => 
                           n61485, A => n8867, ZN => n8862);
   U7275 : OAI221_X1 port map( B1 => n2937, B2 => n61500, C1 => n2877, C2 => 
                           n61497, A => n8866, ZN => n8863);
   U7276 : NOR4_X1 port map( A1 => n8786, A2 => n8787, A3 => n8788, A4 => n8789
                           , ZN => n8758);
   U7277 : OAI221_X1 port map( B1 => n1670, B2 => n61476, C1 => n414, C2 => 
                           n61473, A => n8793, ZN => n8786);
   U7278 : OAI221_X1 port map( B1 => n4715, B2 => n61488, C1 => n53029, C2 => 
                           n61485, A => n8792, ZN => n8787);
   U7279 : OAI221_X1 port map( B1 => n2936, B2 => n61500, C1 => n2876, C2 => 
                           n61497, A => n8791, ZN => n8788);
   U7280 : NOR4_X1 port map( A1 => n8711, A2 => n8712, A3 => n8713, A4 => n8714
                           , ZN => n8683);
   U7281 : OAI221_X1 port map( B1 => n1669, B2 => n61476, C1 => n413, C2 => 
                           n61473, A => n8718, ZN => n8711);
   U7282 : OAI221_X1 port map( B1 => n4714, B2 => n61488, C1 => n53028, C2 => 
                           n61485, A => n8717, ZN => n8712);
   U7283 : OAI221_X1 port map( B1 => n2935, B2 => n61500, C1 => n2875, C2 => 
                           n61497, A => n8716, ZN => n8713);
   U7284 : NOR4_X1 port map( A1 => n15017, A2 => n15018, A3 => n15019, A4 => 
                           n15020, ZN => n14968);
   U7285 : OAI221_X1 port map( B1 => n1692, B2 => n61475, C1 => n452, C2 => 
                           n61472, A => n15025, ZN => n15017);
   U7286 : OAI221_X1 port map( B1 => n4737, B2 => n61487, C1 => n53051, C2 => 
                           n61484, A => n15024, ZN => n15018);
   U7287 : OAI221_X1 port map( B1 => n2958, B2 => n61499, C1 => n2934, C2 => 
                           n61496, A => n15022, ZN => n15019);
   U7288 : NOR4_X1 port map( A1 => n14921, A2 => n14922, A3 => n14923, A4 => 
                           n14924, ZN => n14893);
   U7289 : OAI221_X1 port map( B1 => n1691, B2 => n61475, C1 => n435, C2 => 
                           n61472, A => n14928, ZN => n14921);
   U7290 : OAI221_X1 port map( B1 => n4736, B2 => n61487, C1 => n53050, C2 => 
                           n61484, A => n14927, ZN => n14922);
   U7291 : OAI221_X1 port map( B1 => n2957, B2 => n61499, C1 => n2933, C2 => 
                           n61496, A => n14926, ZN => n14923);
   U7292 : NOR4_X1 port map( A1 => n14846, A2 => n14847, A3 => n14848, A4 => 
                           n14849, ZN => n14818);
   U7293 : OAI221_X1 port map( B1 => n1690, B2 => n61475, C1 => n434, C2 => 
                           n61472, A => n14853, ZN => n14846);
   U7294 : OAI221_X1 port map( B1 => n4735, B2 => n61487, C1 => n53049, C2 => 
                           n61484, A => n14852, ZN => n14847);
   U7295 : OAI221_X1 port map( B1 => n2956, B2 => n61499, C1 => n2932, C2 => 
                           n61496, A => n14851, ZN => n14848);
   U7296 : NOR4_X1 port map( A1 => n14771, A2 => n14772, A3 => n14773, A4 => 
                           n14774, ZN => n14743);
   U7297 : OAI221_X1 port map( B1 => n1689, B2 => n61475, C1 => n433, C2 => 
                           n61472, A => n14778, ZN => n14771);
   U7298 : OAI221_X1 port map( B1 => n4734, B2 => n61487, C1 => n53048, C2 => 
                           n61484, A => n14777, ZN => n14772);
   U7299 : OAI221_X1 port map( B1 => n2955, B2 => n61499, C1 => n2931, C2 => 
                           n61496, A => n14776, ZN => n14773);
   U7300 : NOR4_X1 port map( A1 => n14696, A2 => n14697, A3 => n14698, A4 => 
                           n14699, ZN => n14668);
   U7301 : OAI221_X1 port map( B1 => n1688, B2 => n61475, C1 => n432, C2 => 
                           n61472, A => n14703, ZN => n14696);
   U7302 : OAI221_X1 port map( B1 => n4733, B2 => n61487, C1 => n53047, C2 => 
                           n61484, A => n14702, ZN => n14697);
   U7303 : OAI221_X1 port map( B1 => n2954, B2 => n61499, C1 => n2930, C2 => 
                           n61496, A => n14701, ZN => n14698);
   U7304 : NOR4_X1 port map( A1 => n14621, A2 => n14622, A3 => n14623, A4 => 
                           n14624, ZN => n14593);
   U7305 : OAI221_X1 port map( B1 => n1687, B2 => n61475, C1 => n431, C2 => 
                           n61472, A => n14628, ZN => n14621);
   U7306 : OAI221_X1 port map( B1 => n4732, B2 => n61487, C1 => n53046, C2 => 
                           n61484, A => n14627, ZN => n14622);
   U7307 : OAI221_X1 port map( B1 => n2953, B2 => n61499, C1 => n2929, C2 => 
                           n61496, A => n14626, ZN => n14623);
   U7308 : NOR4_X1 port map( A1 => n14546, A2 => n14547, A3 => n14548, A4 => 
                           n14549, ZN => n14518);
   U7309 : OAI221_X1 port map( B1 => n1686, B2 => n61475, C1 => n430, C2 => 
                           n61472, A => n14553, ZN => n14546);
   U7310 : OAI221_X1 port map( B1 => n4731, B2 => n61487, C1 => n53045, C2 => 
                           n61484, A => n14552, ZN => n14547);
   U7311 : OAI221_X1 port map( B1 => n2952, B2 => n61499, C1 => n2928, C2 => 
                           n61496, A => n14551, ZN => n14548);
   U7312 : NOR4_X1 port map( A1 => n14471, A2 => n14472, A3 => n14473, A4 => 
                           n14474, ZN => n14443);
   U7313 : OAI221_X1 port map( B1 => n1685, B2 => n61475, C1 => n429, C2 => 
                           n61472, A => n14478, ZN => n14471);
   U7314 : OAI221_X1 port map( B1 => n4730, B2 => n61487, C1 => n53044, C2 => 
                           n61484, A => n14477, ZN => n14472);
   U7315 : OAI221_X1 port map( B1 => n2951, B2 => n61499, C1 => n2927, C2 => 
                           n61496, A => n14476, ZN => n14473);
   U7316 : NOR4_X1 port map( A1 => n8636, A2 => n8637, A3 => n8638, A4 => n8639
                           , ZN => n8608);
   U7317 : OAI221_X1 port map( B1 => n505, B2 => n61477, C1 => n388, C2 => 
                           n61474, A => n8643, ZN => n8636);
   U7318 : OAI221_X1 port map( B1 => n562, B2 => n61489, C1 => n494, C2 => 
                           n61486, A => n8642, ZN => n8637);
   U7319 : OAI221_X1 port map( B1 => n770, B2 => n61501, C1 => n762, C2 => 
                           n61498, A => n8641, ZN => n8638);
   U7320 : NOR4_X1 port map( A1 => n8561, A2 => n8562, A3 => n8563, A4 => n8564
                           , ZN => n8533);
   U7321 : OAI221_X1 port map( B1 => n504, B2 => n61477, C1 => n371, C2 => 
                           n61474, A => n8568, ZN => n8561);
   U7322 : OAI221_X1 port map( B1 => n561, B2 => n61489, C1 => n493, C2 => 
                           n61486, A => n8567, ZN => n8562);
   U7323 : OAI221_X1 port map( B1 => n769, B2 => n61501, C1 => n761, C2 => 
                           n61498, A => n8566, ZN => n8563);
   U7324 : NOR4_X1 port map( A1 => n8486, A2 => n8487, A3 => n8488, A4 => n8489
                           , ZN => n8458);
   U7325 : OAI221_X1 port map( B1 => n503, B2 => n61477, C1 => n370, C2 => 
                           n61474, A => n8493, ZN => n8486);
   U7326 : OAI221_X1 port map( B1 => n560, B2 => n61489, C1 => n492, C2 => 
                           n61486, A => n8492, ZN => n8487);
   U7327 : OAI221_X1 port map( B1 => n768, B2 => n61501, C1 => n760, C2 => 
                           n61498, A => n8491, ZN => n8488);
   U7328 : NOR4_X1 port map( A1 => n8411, A2 => n8412, A3 => n8413, A4 => n8414
                           , ZN => n8383);
   U7329 : OAI221_X1 port map( B1 => n502, B2 => n61477, C1 => n369, C2 => 
                           n61474, A => n8418, ZN => n8411);
   U7330 : OAI221_X1 port map( B1 => n499, B2 => n61489, C1 => n491, C2 => 
                           n61486, A => n8417, ZN => n8412);
   U7331 : OAI221_X1 port map( B1 => n767, B2 => n61501, C1 => n567, C2 => 
                           n61498, A => n8416, ZN => n8413);
   U7332 : NOR4_X1 port map( A1 => n8336, A2 => n8337, A3 => n8338, A4 => n8339
                           , ZN => n8308);
   U7333 : OAI221_X1 port map( B1 => n501, B2 => n61477, C1 => n368, C2 => 
                           n61474, A => n8343, ZN => n8336);
   U7334 : OAI221_X1 port map( B1 => n498, B2 => n61489, C1 => n490, C2 => 
                           n61486, A => n8342, ZN => n8337);
   U7335 : OAI221_X1 port map( B1 => n766, B2 => n61501, C1 => n566, C2 => 
                           n61498, A => n8341, ZN => n8338);
   U7336 : NOR4_X1 port map( A1 => n8261, A2 => n8262, A3 => n8263, A4 => n8264
                           , ZN => n8233);
   U7337 : OAI221_X1 port map( B1 => n500, B2 => n61477, C1 => n367, C2 => 
                           n61474, A => n8268, ZN => n8261);
   U7338 : OAI221_X1 port map( B1 => n497, B2 => n61489, C1 => n489, C2 => 
                           n61486, A => n8267, ZN => n8262);
   U7339 : OAI221_X1 port map( B1 => n765, B2 => n61501, C1 => n565, C2 => 
                           n61498, A => n8266, ZN => n8263);
   U7340 : NOR4_X1 port map( A1 => n8186, A2 => n8187, A3 => n8188, A4 => n8189
                           , ZN => n8158);
   U7341 : OAI221_X1 port map( B1 => n475, B2 => n61477, C1 => n366, C2 => 
                           n61474, A => n8193, ZN => n8186);
   U7342 : OAI221_X1 port map( B1 => n496, B2 => n61489, C1 => n488, C2 => 
                           n61486, A => n8192, ZN => n8187);
   U7343 : OAI221_X1 port map( B1 => n764, B2 => n61501, C1 => n564, C2 => 
                           n61498, A => n8191, ZN => n8188);
   U7344 : NOR4_X1 port map( A1 => n8026, A2 => n8027, A3 => n8028, A4 => n8029
                           , ZN => n7947);
   U7345 : OAI221_X1 port map( B1 => n474, B2 => n61477, C1 => n365, C2 => 
                           n61474, A => n8047, ZN => n8026);
   U7346 : OAI221_X1 port map( B1 => n495, B2 => n61489, C1 => n487, C2 => 
                           n61486, A => n8042, ZN => n8027);
   U7347 : OAI221_X1 port map( B1 => n763, B2 => n61501, C1 => n563, C2 => 
                           n61498, A => n8037, ZN => n8028);
   U7348 : OAI221_X1 port map( B1 => n5435, B2 => n4288, C1 => n5436, C2 => 
                           n4280, A => n6045, ZN => n6038);
   U7349 : AOI22_X1 port map( A1 => n16437, A2 => n61884, B1 => n16445, B2 => 
                           n61881, ZN => n6045);
   U7350 : OAI221_X1 port map( B1 => n5435, B2 => n4287, C1 => n5436, C2 => 
                           n4279, A => n5959, ZN => n5954);
   U7351 : AOI22_X1 port map( A1 => n16438, A2 => n61884, B1 => n16446, B2 => 
                           n61881, ZN => n5959);
   U7352 : OAI221_X1 port map( B1 => n5435, B2 => n4286, C1 => n5436, C2 => 
                           n4278, A => n5884, ZN => n5879);
   U7353 : AOI22_X1 port map( A1 => n16439, A2 => n61884, B1 => n16447, B2 => 
                           n61881, ZN => n5884);
   U7354 : OAI221_X1 port map( B1 => n5435, B2 => n4285, C1 => n5436, C2 => 
                           n4277, A => n5809, ZN => n5804);
   U7355 : AOI22_X1 port map( A1 => n16440, A2 => n61884, B1 => n16448, B2 => 
                           n61881, ZN => n5809);
   U7356 : OAI221_X1 port map( B1 => n5435, B2 => n4284, C1 => n5436, C2 => 
                           n4276, A => n5734, ZN => n5729);
   U7357 : AOI22_X1 port map( A1 => n16441, A2 => n61884, B1 => n16449, B2 => 
                           n61881, ZN => n5734);
   U7358 : OAI221_X1 port map( B1 => n5435, B2 => n4283, C1 => n5436, C2 => 
                           n4275, A => n5659, ZN => n5654);
   U7359 : AOI22_X1 port map( A1 => n16442, A2 => n61884, B1 => n16450, B2 => 
                           n61881, ZN => n5659);
   U7360 : OAI221_X1 port map( B1 => n5435, B2 => n4282, C1 => n5436, C2 => 
                           n4274, A => n5584, ZN => n5579);
   U7361 : AOI22_X1 port map( A1 => n16443, A2 => n61884, B1 => n16451, B2 => 
                           n61881, ZN => n5584);
   U7362 : OAI221_X1 port map( B1 => n5435, B2 => n4281, C1 => n5436, C2 => 
                           n4273, A => n5437, ZN => n5424);
   U7363 : AOI22_X1 port map( A1 => n16444, A2 => n61884, B1 => n16452, B2 => 
                           n61881, ZN => n5437);
   U7364 : OAI221_X1 port map( B1 => n5397, B2 => n4147, C1 => n5398, C2 => 
                           n468, A => n6023, ZN => n6012);
   U7365 : AOI222_X1 port map( A1 => n51655, A2 => n61936, B1 => n16413, B2 => 
                           n61724, C1 => n51607, C2 => n59646, ZN => n6023);
   U7366 : OAI221_X1 port map( B1 => n5397, B2 => n4146, C1 => n5398, C2 => 
                           n467, A => n5944, ZN => n5937);
   U7367 : AOI222_X1 port map( A1 => n51654, A2 => n61936, B1 => n16414, B2 => 
                           n61724, C1 => n51606, C2 => n59646, ZN => n5944);
   U7368 : OAI221_X1 port map( B1 => n5397, B2 => n4145, C1 => n5398, C2 => 
                           n466, A => n5869, ZN => n5862);
   U7369 : AOI222_X1 port map( A1 => n51653, A2 => n61936, B1 => n16415, B2 => 
                           n61724, C1 => n51605, C2 => n59646, ZN => n5869);
   U7370 : OAI221_X1 port map( B1 => n5397, B2 => n4144, C1 => n5398, C2 => 
                           n465, A => n5794, ZN => n5787);
   U7371 : AOI222_X1 port map( A1 => n51652, A2 => n61936, B1 => n16416, B2 => 
                           n61724, C1 => n51604, C2 => n59646, ZN => n5794);
   U7372 : OAI221_X1 port map( B1 => n5397, B2 => n4143, C1 => n5398, C2 => 
                           n464, A => n5719, ZN => n5712);
   U7373 : AOI222_X1 port map( A1 => n51651, A2 => n61936, B1 => n16417, B2 => 
                           n61724, C1 => n51603, C2 => n59646, ZN => n5719);
   U7374 : OAI221_X1 port map( B1 => n5397, B2 => n4142, C1 => n5398, C2 => 
                           n463, A => n5644, ZN => n5637);
   U7375 : AOI222_X1 port map( A1 => n51650, A2 => n61936, B1 => n16418, B2 => 
                           n61724, C1 => n51602, C2 => n59646, ZN => n5644);
   U7376 : OAI221_X1 port map( B1 => n5397, B2 => n4141, C1 => n5398, C2 => 
                           n462, A => n5569, ZN => n5562);
   U7377 : AOI222_X1 port map( A1 => n51649, A2 => n61936, B1 => n16419, B2 => 
                           n61724, C1 => n51601, C2 => n59646, ZN => n5569);
   U7378 : OAI221_X1 port map( B1 => n5397, B2 => n4140, C1 => n5398, C2 => 
                           n461, A => n5399, ZN => n5382);
   U7379 : AOI222_X1 port map( A1 => n51648, A2 => n61936, B1 => n16420, B2 => 
                           n61724, C1 => n51600, C2 => n59646, ZN => n5399);
   U7380 : OAI221_X1 port map( B1 => n5503, B2 => n1242, C1 => n5504, C2 => 
                           n159, A => n6090, ZN => n6079);
   U7381 : AOI222_X1 port map( A1 => n15363, A2 => n61820, B1 => n1574, B2 => 
                           n61678, C1 => n52599, C2 => n59647, ZN => n6090);
   U7382 : OAI221_X1 port map( B1 => n5503, B2 => n1241, C1 => n5504, C2 => 
                           n158, A => n5988, ZN => n5981);
   U7383 : AOI222_X1 port map( A1 => n15364, A2 => n61820, B1 => n1573, B2 => 
                           n61678, C1 => n52598, C2 => n59647, ZN => n5988);
   U7384 : OAI221_X1 port map( B1 => n5503, B2 => n1240, C1 => n5504, C2 => 
                           n157, A => n5913, ZN => n5906);
   U7385 : AOI222_X1 port map( A1 => n15365, A2 => n61820, B1 => n1572, B2 => 
                           n61678, C1 => n52597, C2 => n59647, ZN => n5913);
   U7386 : OAI221_X1 port map( B1 => n5503, B2 => n1239, C1 => n5504, C2 => 
                           n156, A => n5838, ZN => n5831);
   U7387 : AOI222_X1 port map( A1 => n15366, A2 => n61820, B1 => n1571, B2 => 
                           n61678, C1 => n52596, C2 => n59647, ZN => n5838);
   U7388 : OAI221_X1 port map( B1 => n5503, B2 => n1238, C1 => n5504, C2 => 
                           n155, A => n5763, ZN => n5756);
   U7389 : AOI222_X1 port map( A1 => n15367, A2 => n61820, B1 => n1570, B2 => 
                           n61678, C1 => n52595, C2 => n59647, ZN => n5763);
   U7390 : OAI221_X1 port map( B1 => n5503, B2 => n1237, C1 => n5504, C2 => 
                           n154, A => n5688, ZN => n5681);
   U7391 : AOI222_X1 port map( A1 => n15368, A2 => n61820, B1 => n1569, B2 => 
                           n61678, C1 => n52594, C2 => n59647, ZN => n5688);
   U7392 : OAI221_X1 port map( B1 => n5503, B2 => n1236, C1 => n5504, C2 => 
                           n153, A => n5613, ZN => n5606);
   U7393 : AOI222_X1 port map( A1 => n15369, A2 => n61821, B1 => n1568, B2 => 
                           n61678, C1 => n52593, C2 => n59647, ZN => n5613);
   U7394 : OAI221_X1 port map( B1 => n5503, B2 => n1235, C1 => n5504, C2 => 
                           n152, A => n5505, ZN => n5488);
   U7395 : AOI222_X1 port map( A1 => n15370, A2 => n61820, B1 => n1567, B2 => 
                           n61678, C1 => n52592, C2 => n59647, ZN => n5505);
   U7396 : OAI221_X1 port map( B1 => n15306, B2 => n5448, C1 => n15338, C2 => 
                           n5449, A => n6053, ZN => n6052);
   U7397 : AOI22_X1 port map( A1 => n16461, A2 => n61875, B1 => n16453, B2 => 
                           n61872, ZN => n6053);
   U7398 : OAI221_X1 port map( B1 => n15305, B2 => n5448, C1 => n15337, C2 => 
                           n5449, A => n5965, ZN => n5964);
   U7399 : AOI22_X1 port map( A1 => n16462, A2 => n61875, B1 => n16454, B2 => 
                           n61872, ZN => n5965);
   U7400 : OAI221_X1 port map( B1 => n15304, B2 => n5448, C1 => n15336, C2 => 
                           n5449, A => n5890, ZN => n5889);
   U7401 : AOI22_X1 port map( A1 => n16463, A2 => n61875, B1 => n16455, B2 => 
                           n61872, ZN => n5890);
   U7402 : OAI221_X1 port map( B1 => n15303, B2 => n5448, C1 => n15335, C2 => 
                           n5449, A => n5815, ZN => n5814);
   U7403 : AOI22_X1 port map( A1 => n16464, A2 => n61875, B1 => n16456, B2 => 
                           n61872, ZN => n5815);
   U7404 : OAI221_X1 port map( B1 => n15302, B2 => n5448, C1 => n15334, C2 => 
                           n5449, A => n5740, ZN => n5739);
   U7405 : AOI22_X1 port map( A1 => n16465, A2 => n61875, B1 => n16457, B2 => 
                           n61872, ZN => n5740);
   U7406 : OAI221_X1 port map( B1 => n15301, B2 => n5448, C1 => n15333, C2 => 
                           n5449, A => n5665, ZN => n5664);
   U7407 : AOI22_X1 port map( A1 => n16466, A2 => n61875, B1 => n16458, B2 => 
                           n61872, ZN => n5665);
   U7408 : OAI221_X1 port map( B1 => n15300, B2 => n5448, C1 => n15332, C2 => 
                           n5449, A => n5590, ZN => n5589);
   U7409 : AOI22_X1 port map( A1 => n16467, A2 => n61875, B1 => n16459, B2 => 
                           n61872, ZN => n5590);
   U7410 : OAI221_X1 port map( B1 => n15299, B2 => n5448, C1 => n15331, C2 => 
                           n5449, A => n5450, ZN => n5447);
   U7411 : AOI22_X1 port map( A1 => n16468, A2 => n61875, B1 => n16460, B2 => 
                           n61872, ZN => n5450);
   U7412 : OAI221_X1 port map( B1 => n61723, B2 => n4589, C1 => n581, C2 => 
                           n61725, A => n7105, ZN => n7104);
   U7413 : AOI22_X1 port map( A1 => n61877, A2 => n4919, B1 => n749, B2 => 
                           n62165, ZN => n7105);
   U7414 : OAI221_X1 port map( B1 => n61723, B2 => n4588, C1 => n580, C2 => 
                           n61725, A => n7030, ZN => n7029);
   U7415 : AOI22_X1 port map( A1 => n61877, A2 => n4918, B1 => n748, B2 => 
                           n62165, ZN => n7030);
   U7416 : OAI221_X1 port map( B1 => n61723, B2 => n4591, C1 => n583, C2 => 
                           n61725, A => n7255, ZN => n7254);
   U7417 : AOI22_X1 port map( A1 => n61877, A2 => n4921, B1 => n751, B2 => 
                           n62165, ZN => n7255);
   U7418 : OAI221_X1 port map( B1 => n61723, B2 => n4599, C1 => n591, C2 => 
                           n61725, A => n7869, ZN => n7868);
   U7419 : AOI22_X1 port map( A1 => n61878, A2 => n4929, B1 => n759, B2 => 
                           n62165, ZN => n7869);
   U7420 : OAI221_X1 port map( B1 => n61723, B2 => n4598, C1 => n590, C2 => 
                           n61725, A => n7780, ZN => n7779);
   U7421 : AOI22_X1 port map( A1 => n61878, A2 => n4928, B1 => n758, B2 => 
                           n62165, ZN => n7780);
   U7422 : OAI221_X1 port map( B1 => n61723, B2 => n4597, C1 => n589, C2 => 
                           n61725, A => n7705, ZN => n7704);
   U7423 : AOI22_X1 port map( A1 => n61878, A2 => n4927, B1 => n757, B2 => 
                           n62165, ZN => n7705);
   U7424 : OAI221_X1 port map( B1 => n61723, B2 => n4596, C1 => n588, C2 => 
                           n61725, A => n7630, ZN => n7629);
   U7425 : AOI22_X1 port map( A1 => n61878, A2 => n4926, B1 => n756, B2 => 
                           n62165, ZN => n7630);
   U7426 : OAI221_X1 port map( B1 => n61723, B2 => n4595, C1 => n587, C2 => 
                           n61725, A => n7555, ZN => n7554);
   U7427 : AOI22_X1 port map( A1 => n61878, A2 => n4925, B1 => n755, B2 => 
                           n62165, ZN => n7555);
   U7428 : OAI221_X1 port map( B1 => n61723, B2 => n4594, C1 => n586, C2 => 
                           n61725, A => n7480, ZN => n7479);
   U7429 : AOI22_X1 port map( A1 => n61878, A2 => n4924, B1 => n754, B2 => 
                           n62165, ZN => n7480);
   U7430 : OAI221_X1 port map( B1 => n61723, B2 => n4593, C1 => n585, C2 => 
                           n61725, A => n7405, ZN => n7404);
   U7431 : AOI22_X1 port map( A1 => n61878, A2 => n4923, B1 => n753, B2 => 
                           n62165, ZN => n7405);
   U7432 : OAI221_X1 port map( B1 => n61723, B2 => n4592, C1 => n584, C2 => 
                           n61725, A => n7330, ZN => n7329);
   U7433 : AOI22_X1 port map( A1 => n61878, A2 => n4922, B1 => n752, B2 => 
                           n62165, ZN => n7330);
   U7434 : OAI221_X1 port map( B1 => n61723, B2 => n4590, C1 => n582, C2 => 
                           n61725, A => n7180, ZN => n7179);
   U7435 : AOI22_X1 port map( A1 => n61877, A2 => n4920, B1 => n750, B2 => 
                           n62165, ZN => n7180);
   U7436 : OAI221_X1 port map( B1 => n421, B2 => n61865, C1 => n1677, C2 => 
                           n61862, A => n6758, ZN => n6757);
   U7437 : AOI22_X1 port map( A1 => n16781, A2 => n62174, B1 => n54380, B2 => 
                           n62126, ZN => n6758);
   U7438 : OAI221_X1 port map( B1 => n2351, B2 => n6107, C1 => n2375, C2 => 
                           n61676, A => n6782, ZN => n6781);
   U7439 : AOI22_X1 port map( A1 => n53736, A2 => n62150, B1 => n53688, B2 => 
                           n62148, ZN => n6782);
   U7440 : OAI221_X1 port map( B1 => n420, B2 => n61865, C1 => n1676, C2 => 
                           n61862, A => n6683, ZN => n6682);
   U7441 : AOI22_X1 port map( A1 => n16782, A2 => n62174, B1 => n54379, B2 => 
                           n62126, ZN => n6683);
   U7442 : OAI221_X1 port map( B1 => n2350, B2 => n6107, C1 => n2374, C2 => 
                           n61676, A => n6707, ZN => n6706);
   U7443 : AOI22_X1 port map( A1 => n53735, A2 => n62150, B1 => n53687, B2 => 
                           n62148, ZN => n6707);
   U7444 : OAI221_X1 port map( B1 => n419, B2 => n61865, C1 => n1675, C2 => 
                           n61862, A => n6608, ZN => n6607);
   U7445 : AOI22_X1 port map( A1 => n16783, A2 => n62174, B1 => n54378, B2 => 
                           n62126, ZN => n6608);
   U7446 : OAI221_X1 port map( B1 => n2349, B2 => n6107, C1 => n2373, C2 => 
                           n61676, A => n6632, ZN => n6631);
   U7447 : AOI22_X1 port map( A1 => n53734, A2 => n62150, B1 => n53686, B2 => 
                           n62148, ZN => n6632);
   U7448 : OAI221_X1 port map( B1 => n418, B2 => n61865, C1 => n1674, C2 => 
                           n61862, A => n6533, ZN => n6532);
   U7449 : AOI22_X1 port map( A1 => n16784, A2 => n62174, B1 => n54377, B2 => 
                           n62126, ZN => n6533);
   U7450 : OAI221_X1 port map( B1 => n2348, B2 => n6107, C1 => n2372, C2 => 
                           n61676, A => n6557, ZN => n6556);
   U7451 : AOI22_X1 port map( A1 => n53733, A2 => n62150, B1 => n53685, B2 => 
                           n62148, ZN => n6557);
   U7452 : OAI221_X1 port map( B1 => n417, B2 => n61865, C1 => n1673, C2 => 
                           n61862, A => n6458, ZN => n6457);
   U7453 : AOI22_X1 port map( A1 => n16785, A2 => n62174, B1 => n54376, B2 => 
                           n62126, ZN => n6458);
   U7454 : OAI221_X1 port map( B1 => n2347, B2 => n6107, C1 => n2371, C2 => 
                           n61676, A => n6482, ZN => n6481);
   U7455 : AOI22_X1 port map( A1 => n53732, A2 => n62150, B1 => n53684, B2 => 
                           n62148, ZN => n6482);
   U7456 : OAI221_X1 port map( B1 => n416, B2 => n61864, C1 => n1672, C2 => 
                           n61862, A => n6383, ZN => n6382);
   U7457 : AOI22_X1 port map( A1 => n16786, A2 => n62174, B1 => n54375, B2 => 
                           n62126, ZN => n6383);
   U7458 : OAI221_X1 port map( B1 => n2346, B2 => n6107, C1 => n2370, C2 => 
                           n61676, A => n6407, ZN => n6406);
   U7459 : AOI22_X1 port map( A1 => n53731, A2 => n62150, B1 => n53683, B2 => 
                           n62148, ZN => n6407);
   U7460 : OAI221_X1 port map( B1 => n415, B2 => n61864, C1 => n1671, C2 => 
                           n61862, A => n6308, ZN => n6307);
   U7461 : AOI22_X1 port map( A1 => n16787, A2 => n62174, B1 => n54374, B2 => 
                           n62126, ZN => n6308);
   U7462 : OAI221_X1 port map( B1 => n2345, B2 => n6107, C1 => n2369, C2 => 
                           n61676, A => n6332, ZN => n6331);
   U7463 : AOI22_X1 port map( A1 => n53730, A2 => n62150, B1 => n53682, B2 => 
                           n62148, ZN => n6332);
   U7464 : OAI221_X1 port map( B1 => n414, B2 => n61864, C1 => n1670, C2 => 
                           n61862, A => n6233, ZN => n6232);
   U7465 : AOI22_X1 port map( A1 => n16788, A2 => n62174, B1 => n54373, B2 => 
                           n62126, ZN => n6233);
   U7466 : OAI221_X1 port map( B1 => n2344, B2 => n6107, C1 => n2368, C2 => 
                           n61676, A => n6257, ZN => n6256);
   U7467 : AOI22_X1 port map( A1 => n53729, A2 => n62150, B1 => n53681, B2 => 
                           n62148, ZN => n6257);
   U7468 : OAI221_X1 port map( B1 => n413, B2 => n61864, C1 => n1669, C2 => 
                           n61862, A => n6158, ZN => n6157);
   U7469 : AOI22_X1 port map( A1 => n16789, A2 => n62174, B1 => n54372, B2 => 
                           n62126, ZN => n6158);
   U7470 : OAI221_X1 port map( B1 => n2343, B2 => n6107, C1 => n2367, C2 => 
                           n61676, A => n6182, ZN => n6181);
   U7471 : AOI22_X1 port map( A1 => n53728, A2 => n62150, B1 => n53680, B2 => 
                           n62148, ZN => n6182);
   U7472 : OAI221_X1 port map( B1 => n426, B2 => n61865, C1 => n1682, C2 => 
                           n61861, A => n7133, ZN => n7132);
   U7473 : AOI22_X1 port map( A1 => n16776, A2 => n62175, B1 => n54385, B2 => 
                           n62127, ZN => n7133);
   U7474 : OAI221_X1 port map( B1 => n2356, B2 => n61673, C1 => n2380, C2 => 
                           n61675, A => n7157, ZN => n7156);
   U7475 : AOI22_X1 port map( A1 => n53741, A2 => n62151, B1 => n53693, B2 => 
                           n62149, ZN => n7157);
   U7476 : OAI221_X1 port map( B1 => n425, B2 => n61865, C1 => n1681, C2 => 
                           n61861, A => n7058, ZN => n7057);
   U7477 : AOI22_X1 port map( A1 => n16777, A2 => n62175, B1 => n54384, B2 => 
                           n62127, ZN => n7058);
   U7478 : OAI221_X1 port map( B1 => n2355, B2 => n61673, C1 => n2379, C2 => 
                           n61675, A => n7082, ZN => n7081);
   U7479 : AOI22_X1 port map( A1 => n53740, A2 => n62151, B1 => n53692, B2 => 
                           n62149, ZN => n7082);
   U7480 : OAI221_X1 port map( B1 => n423, B2 => n61865, C1 => n1679, C2 => 
                           n61862, A => n6908, ZN => n6907);
   U7481 : AOI22_X1 port map( A1 => n16779, A2 => n62174, B1 => n54382, B2 => 
                           n62126, ZN => n6908);
   U7482 : OAI221_X1 port map( B1 => n2353, B2 => n6107, C1 => n2377, C2 => 
                           n61676, A => n6932, ZN => n6931);
   U7483 : AOI22_X1 port map( A1 => n53738, A2 => n62150, B1 => n53690, B2 => 
                           n62148, ZN => n6932);
   U7484 : OAI221_X1 port map( B1 => n422, B2 => n61865, C1 => n1678, C2 => 
                           n61862, A => n6833, ZN => n6832);
   U7485 : AOI22_X1 port map( A1 => n16780, A2 => n62174, B1 => n54381, B2 => 
                           n62126, ZN => n6833);
   U7486 : OAI221_X1 port map( B1 => n2352, B2 => n6107, C1 => n2376, C2 => 
                           n61676, A => n6857, ZN => n6856);
   U7487 : AOI22_X1 port map( A1 => n53737, A2 => n62150, B1 => n53689, B2 => 
                           n62148, ZN => n6857);
   U7488 : OAI221_X1 port map( B1 => n428, B2 => n61865, C1 => n1684, C2 => 
                           n61861, A => n7283, ZN => n7282);
   U7489 : AOI22_X1 port map( A1 => n16774, A2 => n62175, B1 => n54387, B2 => 
                           n62127, ZN => n7283);
   U7490 : OAI221_X1 port map( B1 => n2358, B2 => n61673, C1 => n2382, C2 => 
                           n61675, A => n7307, ZN => n7306);
   U7491 : AOI22_X1 port map( A1 => n53743, A2 => n62151, B1 => n53695, B2 => 
                           n62149, ZN => n7307);
   U7492 : OAI221_X1 port map( B1 => n452, B2 => n61866, C1 => n1692, C2 => 
                           n61861, A => n7908, ZN => n7907);
   U7493 : AOI22_X1 port map( A1 => n16766, A2 => n62175, B1 => n54395, B2 => 
                           n62127, ZN => n7908);
   U7494 : OAI221_X1 port map( B1 => n2366, B2 => n61673, C1 => n2390, C2 => 
                           n61675, A => n7939, ZN => n7938);
   U7495 : AOI22_X1 port map( A1 => n53751, A2 => n62151, B1 => n53703, B2 => 
                           n62149, ZN => n7939);
   U7496 : OAI221_X1 port map( B1 => n435, B2 => n61866, C1 => n1691, C2 => 
                           n61861, A => n7808, ZN => n7807);
   U7497 : AOI22_X1 port map( A1 => n16767, A2 => n62175, B1 => n54394, B2 => 
                           n62127, ZN => n7808);
   U7498 : OAI221_X1 port map( B1 => n2365, B2 => n61673, C1 => n2389, C2 => 
                           n61675, A => n7832, ZN => n7831);
   U7499 : AOI22_X1 port map( A1 => n53750, A2 => n62151, B1 => n53702, B2 => 
                           n62149, ZN => n7832);
   U7500 : OAI221_X1 port map( B1 => n434, B2 => n61866, C1 => n1690, C2 => 
                           n61861, A => n7733, ZN => n7732);
   U7501 : AOI22_X1 port map( A1 => n16768, A2 => n62175, B1 => n54393, B2 => 
                           n62127, ZN => n7733);
   U7502 : OAI221_X1 port map( B1 => n2364, B2 => n61673, C1 => n2388, C2 => 
                           n61675, A => n7757, ZN => n7756);
   U7503 : AOI22_X1 port map( A1 => n53749, A2 => n62151, B1 => n53701, B2 => 
                           n62149, ZN => n7757);
   U7504 : OAI221_X1 port map( B1 => n433, B2 => n61866, C1 => n1689, C2 => 
                           n61861, A => n7658, ZN => n7657);
   U7505 : AOI22_X1 port map( A1 => n16769, A2 => n62175, B1 => n54392, B2 => 
                           n62127, ZN => n7658);
   U7506 : OAI221_X1 port map( B1 => n2363, B2 => n61673, C1 => n2387, C2 => 
                           n61675, A => n7682, ZN => n7681);
   U7507 : AOI22_X1 port map( A1 => n53748, A2 => n62151, B1 => n53700, B2 => 
                           n62149, ZN => n7682);
   U7508 : OAI221_X1 port map( B1 => n432, B2 => n61866, C1 => n1688, C2 => 
                           n61861, A => n7583, ZN => n7582);
   U7509 : AOI22_X1 port map( A1 => n16770, A2 => n62175, B1 => n54391, B2 => 
                           n62127, ZN => n7583);
   U7510 : OAI221_X1 port map( B1 => n2362, B2 => n61673, C1 => n2386, C2 => 
                           n61675, A => n7607, ZN => n7606);
   U7511 : AOI22_X1 port map( A1 => n53747, A2 => n62151, B1 => n53699, B2 => 
                           n62149, ZN => n7607);
   U7512 : OAI221_X1 port map( B1 => n431, B2 => n61866, C1 => n1687, C2 => 
                           n61861, A => n7508, ZN => n7507);
   U7513 : AOI22_X1 port map( A1 => n16771, A2 => n62175, B1 => n54390, B2 => 
                           n62127, ZN => n7508);
   U7514 : OAI221_X1 port map( B1 => n2361, B2 => n61673, C1 => n2385, C2 => 
                           n61675, A => n7532, ZN => n7531);
   U7515 : AOI22_X1 port map( A1 => n53746, A2 => n62151, B1 => n53698, B2 => 
                           n62149, ZN => n7532);
   U7516 : OAI221_X1 port map( B1 => n430, B2 => n61866, C1 => n1686, C2 => 
                           n61861, A => n7433, ZN => n7432);
   U7517 : AOI22_X1 port map( A1 => n16772, A2 => n62175, B1 => n54389, B2 => 
                           n62127, ZN => n7433);
   U7518 : OAI221_X1 port map( B1 => n2360, B2 => n61673, C1 => n2384, C2 => 
                           n61675, A => n7457, ZN => n7456);
   U7519 : AOI22_X1 port map( A1 => n53745, A2 => n62151, B1 => n53697, B2 => 
                           n62149, ZN => n7457);
   U7520 : OAI221_X1 port map( B1 => n429, B2 => n61865, C1 => n1685, C2 => 
                           n61861, A => n7358, ZN => n7357);
   U7521 : AOI22_X1 port map( A1 => n16773, A2 => n62175, B1 => n54388, B2 => 
                           n62127, ZN => n7358);
   U7522 : OAI221_X1 port map( B1 => n2359, B2 => n61673, C1 => n2383, C2 => 
                           n61675, A => n7382, ZN => n7381);
   U7523 : AOI22_X1 port map( A1 => n53744, A2 => n62151, B1 => n53696, B2 => 
                           n62149, ZN => n7382);
   U7524 : OAI221_X1 port map( B1 => n427, B2 => n61865, C1 => n1683, C2 => 
                           n61861, A => n7208, ZN => n7207);
   U7525 : AOI22_X1 port map( A1 => n16775, A2 => n62175, B1 => n54386, B2 => 
                           n62127, ZN => n7208);
   U7526 : OAI221_X1 port map( B1 => n2357, B2 => n61673, C1 => n2381, C2 => 
                           n61675, A => n7232, ZN => n7231);
   U7527 : AOI22_X1 port map( A1 => n53742, A2 => n62151, B1 => n53694, B2 => 
                           n62149, ZN => n7232);
   U7528 : OAI221_X1 port map( B1 => n424, B2 => n61865, C1 => n1680, C2 => 
                           n61862, A => n6983, ZN => n6982);
   U7529 : AOI22_X1 port map( A1 => n16778, A2 => n62174, B1 => n54383, B2 => 
                           n62126, ZN => n6983);
   U7530 : OAI221_X1 port map( B1 => n2354, B2 => n6107, C1 => n2378, C2 => 
                           n61676, A => n7007, ZN => n7006);
   U7531 : AOI22_X1 port map( A1 => n53739, A2 => n62150, B1 => n53691, B2 => 
                           n62148, ZN => n7007);
   U7532 : OAI221_X1 port map( B1 => n2382, B2 => n61307, C1 => n2358, C2 => 
                           n61304, A => n14436, ZN => n14435);
   U7533 : AOI22_X1 port map( A1 => n61301, A2 => n53647, B1 => n61299, B2 => 
                           n53671, ZN => n14436);
   U7534 : OAI221_X1 port map( B1 => n2381, B2 => n61307, C1 => n2357, C2 => 
                           n61304, A => n14361, ZN => n14360);
   U7535 : AOI22_X1 port map( A1 => n61301, A2 => n53646, B1 => n61299, B2 => 
                           n53670, ZN => n14361);
   U7536 : OAI221_X1 port map( B1 => n2380, B2 => n61307, C1 => n2356, C2 => 
                           n61304, A => n9870, ZN => n9869);
   U7537 : AOI22_X1 port map( A1 => n61301, A2 => n53645, B1 => n61299, B2 => 
                           n53669, ZN => n9870);
   U7538 : OAI221_X1 port map( B1 => n2379, B2 => n61307, C1 => n2355, C2 => 
                           n61304, A => n9731, ZN => n9730);
   U7539 : AOI22_X1 port map( A1 => n61301, A2 => n53644, B1 => n61299, B2 => 
                           n53668, ZN => n9731);
   U7540 : OAI221_X1 port map( B1 => n2378, B2 => n61308, C1 => n2354, C2 => 
                           n61305, A => n9656, ZN => n9655);
   U7541 : AOI22_X1 port map( A1 => n61302, A2 => n53643, B1 => n61299, B2 => 
                           n53667, ZN => n9656);
   U7542 : OAI221_X1 port map( B1 => n2377, B2 => n61308, C1 => n2353, C2 => 
                           n61305, A => n9565, ZN => n9564);
   U7543 : AOI22_X1 port map( A1 => n61302, A2 => n53642, B1 => n61299, B2 => 
                           n53666, ZN => n9565);
   U7544 : OAI221_X1 port map( B1 => n2376, B2 => n61308, C1 => n2352, C2 => 
                           n61305, A => n9490, ZN => n9489);
   U7545 : AOI22_X1 port map( A1 => n61302, A2 => n53641, B1 => n61299, B2 => 
                           n53665, ZN => n9490);
   U7546 : OAI221_X1 port map( B1 => n2375, B2 => n61308, C1 => n2351, C2 => 
                           n61305, A => n9415, ZN => n9414);
   U7547 : AOI22_X1 port map( A1 => n61302, A2 => n53640, B1 => n61299, B2 => 
                           n53664, ZN => n9415);
   U7548 : OAI221_X1 port map( B1 => n2374, B2 => n61308, C1 => n2350, C2 => 
                           n61305, A => n9276, ZN => n9275);
   U7549 : AOI22_X1 port map( A1 => n61302, A2 => n53639, B1 => n61299, B2 => 
                           n53663, ZN => n9276);
   U7550 : OAI221_X1 port map( B1 => n2373, B2 => n61308, C1 => n2349, C2 => 
                           n61305, A => n9201, ZN => n9200);
   U7551 : AOI22_X1 port map( A1 => n61302, A2 => n53638, B1 => n61299, B2 => 
                           n53662, ZN => n9201);
   U7552 : OAI221_X1 port map( B1 => n2372, B2 => n61308, C1 => n2348, C2 => 
                           n61305, A => n9126, ZN => n9125);
   U7553 : AOI22_X1 port map( A1 => n61302, A2 => n53637, B1 => n61299, B2 => 
                           n53661, ZN => n9126);
   U7554 : OAI221_X1 port map( B1 => n2371, B2 => n61308, C1 => n2347, C2 => 
                           n61305, A => n9051, ZN => n9050);
   U7555 : AOI22_X1 port map( A1 => n61302, A2 => n53636, B1 => n61299, B2 => 
                           n53660, ZN => n9051);
   U7556 : OAI221_X1 port map( B1 => n2370, B2 => n61308, C1 => n2346, C2 => 
                           n61305, A => n8976, ZN => n8975);
   U7557 : AOI22_X1 port map( A1 => n61302, A2 => n53635, B1 => n61298, B2 => 
                           n53659, ZN => n8976);
   U7558 : OAI221_X1 port map( B1 => n2369, B2 => n61308, C1 => n2345, C2 => 
                           n61305, A => n8901, ZN => n8900);
   U7559 : AOI22_X1 port map( A1 => n61302, A2 => n53634, B1 => n61298, B2 => 
                           n53658, ZN => n8901);
   U7560 : OAI221_X1 port map( B1 => n2368, B2 => n61308, C1 => n2344, C2 => 
                           n61305, A => n8826, ZN => n8825);
   U7561 : AOI22_X1 port map( A1 => n61302, A2 => n53633, B1 => n61298, B2 => 
                           n53657, ZN => n8826);
   U7562 : OAI221_X1 port map( B1 => n2367, B2 => n61308, C1 => n2343, C2 => 
                           n61305, A => n8751, ZN => n8750);
   U7563 : AOI22_X1 port map( A1 => n61302, A2 => n53632, B1 => n61298, B2 => 
                           n53656, ZN => n8751);
   U7564 : OAI221_X1 port map( B1 => n2390, B2 => n61307, C1 => n2366, C2 => 
                           n61304, A => n15067, ZN => n15066);
   U7565 : AOI22_X1 port map( A1 => n61301, A2 => n53655, B1 => n61300, B2 => 
                           n53679, ZN => n15067);
   U7566 : OAI221_X1 port map( B1 => n2389, B2 => n61307, C1 => n2365, C2 => 
                           n61304, A => n14961, ZN => n14960);
   U7567 : AOI22_X1 port map( A1 => n61301, A2 => n53654, B1 => n61300, B2 => 
                           n53678, ZN => n14961);
   U7568 : OAI221_X1 port map( B1 => n2388, B2 => n61307, C1 => n2364, C2 => 
                           n61304, A => n14886, ZN => n14885);
   U7569 : AOI22_X1 port map( A1 => n61301, A2 => n53653, B1 => n61300, B2 => 
                           n53677, ZN => n14886);
   U7570 : OAI221_X1 port map( B1 => n2387, B2 => n61307, C1 => n2363, C2 => 
                           n61304, A => n14811, ZN => n14810);
   U7571 : AOI22_X1 port map( A1 => n61301, A2 => n53652, B1 => n61300, B2 => 
                           n53676, ZN => n14811);
   U7572 : OAI221_X1 port map( B1 => n2386, B2 => n61307, C1 => n2362, C2 => 
                           n61304, A => n14736, ZN => n14735);
   U7573 : AOI22_X1 port map( A1 => n61301, A2 => n53651, B1 => n61300, B2 => 
                           n53675, ZN => n14736);
   U7574 : OAI221_X1 port map( B1 => n2385, B2 => n61307, C1 => n2361, C2 => 
                           n61304, A => n14661, ZN => n14660);
   U7575 : AOI22_X1 port map( A1 => n61301, A2 => n53650, B1 => n61300, B2 => 
                           n53674, ZN => n14661);
   U7576 : OAI221_X1 port map( B1 => n2384, B2 => n61307, C1 => n2360, C2 => 
                           n61304, A => n14586, ZN => n14585);
   U7577 : AOI22_X1 port map( A1 => n61301, A2 => n53649, B1 => n61300, B2 => 
                           n53673, ZN => n14586);
   U7578 : OAI221_X1 port map( B1 => n2383, B2 => n61307, C1 => n2359, C2 => 
                           n61304, A => n14511, ZN => n14510);
   U7579 : AOI22_X1 port map( A1 => n61301, A2 => n53648, B1 => n61300, B2 => 
                           n53672, ZN => n14511);
   U7580 : OAI221_X1 port map( B1 => n802, B2 => n61513, C1 => n794, C2 => 
                           n61510, A => n8640, ZN => n8639);
   U7581 : AOI22_X1 port map( A1 => n61507, A2 => n786, B1 => n61502, B2 => 
                           n554, ZN => n8640);
   U7582 : OAI221_X1 port map( B1 => n1089, B2 => n61309, C1 => n1081, C2 => 
                           n61306, A => n8676, ZN => n8675);
   U7583 : AOI22_X1 port map( A1 => n61303, A2 => n4312, B1 => n61298, B2 => 
                           n52511, ZN => n8676);
   U7584 : OAI221_X1 port map( B1 => n801, B2 => n61513, C1 => n793, C2 => 
                           n61510, A => n8565, ZN => n8564);
   U7585 : AOI22_X1 port map( A1 => n61507, A2 => n785, B1 => n61502, B2 => 
                           n553, ZN => n8565);
   U7586 : OAI221_X1 port map( B1 => n1088, B2 => n61309, C1 => n1080, C2 => 
                           n61306, A => n8601, ZN => n8600);
   U7587 : AOI22_X1 port map( A1 => n61303, A2 => n4311, B1 => n61298, B2 => 
                           n52510, ZN => n8601);
   U7588 : OAI221_X1 port map( B1 => n800, B2 => n61513, C1 => n792, C2 => 
                           n61510, A => n8490, ZN => n8489);
   U7589 : AOI22_X1 port map( A1 => n61507, A2 => n784, B1 => n61502, B2 => 
                           n552, ZN => n8490);
   U7590 : OAI221_X1 port map( B1 => n1087, B2 => n61309, C1 => n1079, C2 => 
                           n61306, A => n8526, ZN => n8525);
   U7591 : AOI22_X1 port map( A1 => n61303, A2 => n4310, B1 => n61298, B2 => 
                           n52509, ZN => n8526);
   U7592 : OAI221_X1 port map( B1 => n799, B2 => n61513, C1 => n791, C2 => 
                           n61510, A => n8415, ZN => n8414);
   U7593 : AOI22_X1 port map( A1 => n61507, A2 => n775, B1 => n61502, B2 => 
                           n551, ZN => n8415);
   U7594 : OAI221_X1 port map( B1 => n1086, B2 => n61309, C1 => n1078, C2 => 
                           n61306, A => n8451, ZN => n8450);
   U7595 : AOI22_X1 port map( A1 => n61303, A2 => n4309, B1 => n61298, B2 => 
                           n52508, ZN => n8451);
   U7596 : OAI221_X1 port map( B1 => n798, B2 => n61513, C1 => n790, C2 => 
                           n61510, A => n8340, ZN => n8339);
   U7597 : AOI22_X1 port map( A1 => n61507, A2 => n774, B1 => n61502, B2 => 
                           n550, ZN => n8340);
   U7598 : OAI221_X1 port map( B1 => n1085, B2 => n61309, C1 => n1077, C2 => 
                           n61306, A => n8376, ZN => n8375);
   U7599 : AOI22_X1 port map( A1 => n61303, A2 => n4308, B1 => n61298, B2 => 
                           n4316, ZN => n8376);
   U7600 : OAI221_X1 port map( B1 => n797, B2 => n61513, C1 => n789, C2 => 
                           n61510, A => n8265, ZN => n8264);
   U7601 : AOI22_X1 port map( A1 => n61507, A2 => n773, B1 => n61502, B2 => 
                           n549, ZN => n8265);
   U7602 : OAI221_X1 port map( B1 => n1084, B2 => n61309, C1 => n1076, C2 => 
                           n61306, A => n8301, ZN => n8300);
   U7603 : AOI22_X1 port map( A1 => n61303, A2 => n4307, B1 => n61298, B2 => 
                           n4315, ZN => n8301);
   U7604 : OAI221_X1 port map( B1 => n796, B2 => n61513, C1 => n788, C2 => 
                           n61510, A => n8190, ZN => n8189);
   U7605 : AOI22_X1 port map( A1 => n61507, A2 => n772, B1 => n61502, B2 => 
                           n548, ZN => n8190);
   U7606 : OAI221_X1 port map( B1 => n1083, B2 => n61309, C1 => n1075, C2 => 
                           n61306, A => n8226, ZN => n8225);
   U7607 : AOI22_X1 port map( A1 => n61303, A2 => n4306, B1 => n61298, B2 => 
                           n4314, ZN => n8226);
   U7608 : OAI221_X1 port map( B1 => n795, B2 => n61513, C1 => n787, C2 => 
                           n61510, A => n8032, ZN => n8029);
   U7609 : AOI22_X1 port map( A1 => n61507, A2 => n771, B1 => n61502, B2 => 
                           n547, ZN => n8032);
   U7610 : OAI221_X1 port map( B1 => n1082, B2 => n61309, C1 => n1074, C2 => 
                           n61306, A => n8136, ZN => n8133);
   U7611 : AOI22_X1 port map( A1 => n61303, A2 => n4305, B1 => n61298, B2 => 
                           n4313, ZN => n8136);
   U7612 : OAI221_X1 port map( B1 => n6025, B2 => n4584, C1 => n576, C2 => 
                           n61726, A => n6730, ZN => n6729);
   U7613 : AOI22_X1 port map( A1 => n61877, A2 => n4914, B1 => n744, B2 => 
                           n62164, ZN => n6730);
   U7614 : OAI221_X1 port map( B1 => n6025, B2 => n4583, C1 => n575, C2 => 
                           n61726, A => n6655, ZN => n6654);
   U7615 : AOI22_X1 port map( A1 => n61877, A2 => n4913, B1 => n743, B2 => 
                           n62164, ZN => n6655);
   U7616 : OAI221_X1 port map( B1 => n6025, B2 => n4582, C1 => n574, C2 => 
                           n61726, A => n6580, ZN => n6579);
   U7617 : AOI22_X1 port map( A1 => n61877, A2 => n4912, B1 => n742, B2 => 
                           n62164, ZN => n6580);
   U7618 : OAI221_X1 port map( B1 => n6025, B2 => n4581, C1 => n573, C2 => 
                           n61726, A => n6505, ZN => n6504);
   U7619 : AOI22_X1 port map( A1 => n61877, A2 => n4911, B1 => n741, B2 => 
                           n62164, ZN => n6505);
   U7620 : OAI221_X1 port map( B1 => n6025, B2 => n4580, C1 => n572, C2 => 
                           n61726, A => n6430, ZN => n6429);
   U7621 : AOI22_X1 port map( A1 => n61877, A2 => n4910, B1 => n740, B2 => 
                           n62164, ZN => n6430);
   U7622 : OAI221_X1 port map( B1 => n6025, B2 => n4579, C1 => n571, C2 => 
                           n61726, A => n6355, ZN => n6354);
   U7623 : AOI22_X1 port map( A1 => n61876, A2 => n4909, B1 => n739, B2 => 
                           n62164, ZN => n6355);
   U7624 : OAI221_X1 port map( B1 => n6025, B2 => n4578, C1 => n570, C2 => 
                           n61726, A => n6280, ZN => n6279);
   U7625 : AOI22_X1 port map( A1 => n61876, A2 => n4908, B1 => n738, B2 => 
                           n62164, ZN => n6280);
   U7626 : OAI221_X1 port map( B1 => n6025, B2 => n4577, C1 => n569, C2 => 
                           n61726, A => n6205, ZN => n6204);
   U7627 : AOI22_X1 port map( A1 => n61876, A2 => n4907, B1 => n737, B2 => 
                           n62164, ZN => n6205);
   U7628 : OAI221_X1 port map( B1 => n6025, B2 => n4576, C1 => n568, C2 => 
                           n61726, A => n6130, ZN => n6129);
   U7629 : AOI22_X1 port map( A1 => n61876, A2 => n4906, B1 => n736, B2 => 
                           n62164, ZN => n6130);
   U7630 : OAI221_X1 port map( B1 => n6025, B2 => n4586, C1 => n578, C2 => 
                           n61726, A => n6880, ZN => n6879);
   U7631 : AOI22_X1 port map( A1 => n61877, A2 => n4916, B1 => n746, B2 => 
                           n62164, ZN => n6880);
   U7632 : OAI221_X1 port map( B1 => n6025, B2 => n4585, C1 => n577, C2 => 
                           n61726, A => n6805, ZN => n6804);
   U7633 : AOI22_X1 port map( A1 => n61877, A2 => n4915, B1 => n745, B2 => 
                           n62164, ZN => n6805);
   U7634 : OAI221_X1 port map( B1 => n6025, B2 => n4587, C1 => n579, C2 => 
                           n61726, A => n6955, ZN => n6954);
   U7635 : AOI22_X1 port map( A1 => n61877, A2 => n4917, B1 => n747, B2 => 
                           n62164, ZN => n6955);
   U7636 : OAI221_X1 port map( B1 => n4777, B2 => n61511, C1 => n4753, C2 => 
                           n61508, A => n14400, ZN => n14399);
   U7637 : AOI22_X1 port map( A1 => n61505, A2 => n703, B1 => n61503, B2 => 
                           n727, ZN => n14400);
   U7638 : OAI221_X1 port map( B1 => n4776, B2 => n61511, C1 => n4752, C2 => 
                           n61508, A => n9909, ZN => n9908);
   U7639 : AOI22_X1 port map( A1 => n61505, A2 => n702, B1 => n61503, B2 => 
                           n726, ZN => n9909);
   U7640 : OAI221_X1 port map( B1 => n4775, B2 => n61511, C1 => n4751, C2 => 
                           n61508, A => n9834, ZN => n9833);
   U7641 : AOI22_X1 port map( A1 => n61505, A2 => n701, B1 => n61503, B2 => 
                           n725, ZN => n9834);
   U7642 : OAI221_X1 port map( B1 => n4774, B2 => n61511, C1 => n4750, C2 => 
                           n61508, A => n9695, ZN => n9694);
   U7643 : AOI22_X1 port map( A1 => n61505, A2 => n700, B1 => n61503, B2 => 
                           n724, ZN => n9695);
   U7644 : OAI221_X1 port map( B1 => n4773, B2 => n61512, C1 => n4749, C2 => 
                           n61509, A => n9620, ZN => n9619);
   U7645 : AOI22_X1 port map( A1 => n61506, A2 => n699, B1 => n61503, B2 => 
                           n723, ZN => n9620);
   U7646 : OAI221_X1 port map( B1 => n4772, B2 => n61512, C1 => n4748, C2 => 
                           n61509, A => n9529, ZN => n9528);
   U7647 : AOI22_X1 port map( A1 => n61506, A2 => n698, B1 => n61503, B2 => 
                           n722, ZN => n9529);
   U7648 : OAI221_X1 port map( B1 => n4771, B2 => n61512, C1 => n4747, C2 => 
                           n61509, A => n9454, ZN => n9453);
   U7649 : AOI22_X1 port map( A1 => n61506, A2 => n697, B1 => n61503, B2 => 
                           n721, ZN => n9454);
   U7650 : OAI221_X1 port map( B1 => n4770, B2 => n61512, C1 => n4746, C2 => 
                           n61509, A => n9379, ZN => n9378);
   U7651 : AOI22_X1 port map( A1 => n61506, A2 => n696, B1 => n61503, B2 => 
                           n720, ZN => n9379);
   U7652 : OAI221_X1 port map( B1 => n4769, B2 => n61512, C1 => n4745, C2 => 
                           n61509, A => n9240, ZN => n9239);
   U7653 : AOI22_X1 port map( A1 => n61506, A2 => n695, B1 => n61503, B2 => 
                           n719, ZN => n9240);
   U7654 : OAI221_X1 port map( B1 => n4768, B2 => n61512, C1 => n4744, C2 => 
                           n61509, A => n9165, ZN => n9164);
   U7655 : AOI22_X1 port map( A1 => n61506, A2 => n694, B1 => n61503, B2 => 
                           n718, ZN => n9165);
   U7656 : OAI221_X1 port map( B1 => n4767, B2 => n61512, C1 => n4743, C2 => 
                           n61509, A => n9090, ZN => n9089);
   U7657 : AOI22_X1 port map( A1 => n61506, A2 => n693, B1 => n61503, B2 => 
                           n717, ZN => n9090);
   U7658 : OAI221_X1 port map( B1 => n4766, B2 => n61512, C1 => n4742, C2 => 
                           n61509, A => n9015, ZN => n9014);
   U7659 : AOI22_X1 port map( A1 => n61506, A2 => n692, B1 => n61503, B2 => 
                           n716, ZN => n9015);
   U7660 : OAI221_X1 port map( B1 => n4765, B2 => n61512, C1 => n4741, C2 => 
                           n61509, A => n8940, ZN => n8939);
   U7661 : AOI22_X1 port map( A1 => n61506, A2 => n691, B1 => n61502, B2 => 
                           n715, ZN => n8940);
   U7662 : OAI221_X1 port map( B1 => n4764, B2 => n61512, C1 => n4740, C2 => 
                           n61509, A => n8865, ZN => n8864);
   U7663 : AOI22_X1 port map( A1 => n61506, A2 => n690, B1 => n61502, B2 => 
                           n714, ZN => n8865);
   U7664 : OAI221_X1 port map( B1 => n4763, B2 => n61512, C1 => n4739, C2 => 
                           n61509, A => n8790, ZN => n8789);
   U7665 : AOI22_X1 port map( A1 => n61506, A2 => n689, B1 => n61502, B2 => 
                           n713, ZN => n8790);
   U7666 : OAI221_X1 port map( B1 => n4762, B2 => n61512, C1 => n4738, C2 => 
                           n61509, A => n8715, ZN => n8714);
   U7667 : AOI22_X1 port map( A1 => n61506, A2 => n688, B1 => n61502, B2 => 
                           n712, ZN => n8715);
   U7668 : OAI221_X1 port map( B1 => n4785, B2 => n61511, C1 => n4761, C2 => 
                           n61508, A => n15021, ZN => n15020);
   U7669 : AOI22_X1 port map( A1 => n61505, A2 => n711, B1 => n61504, B2 => 
                           n735, ZN => n15021);
   U7670 : OAI221_X1 port map( B1 => n4784, B2 => n61511, C1 => n4760, C2 => 
                           n61508, A => n14925, ZN => n14924);
   U7671 : AOI22_X1 port map( A1 => n61505, A2 => n710, B1 => n61504, B2 => 
                           n734, ZN => n14925);
   U7672 : OAI221_X1 port map( B1 => n4783, B2 => n61511, C1 => n4759, C2 => 
                           n61508, A => n14850, ZN => n14849);
   U7673 : AOI22_X1 port map( A1 => n61505, A2 => n709, B1 => n61504, B2 => 
                           n733, ZN => n14850);
   U7674 : OAI221_X1 port map( B1 => n4782, B2 => n61511, C1 => n4758, C2 => 
                           n61508, A => n14775, ZN => n14774);
   U7675 : AOI22_X1 port map( A1 => n61505, A2 => n708, B1 => n61504, B2 => 
                           n732, ZN => n14775);
   U7676 : OAI221_X1 port map( B1 => n4781, B2 => n61511, C1 => n4757, C2 => 
                           n61508, A => n14700, ZN => n14699);
   U7677 : AOI22_X1 port map( A1 => n61505, A2 => n707, B1 => n61504, B2 => 
                           n731, ZN => n14700);
   U7678 : OAI221_X1 port map( B1 => n4780, B2 => n61511, C1 => n4756, C2 => 
                           n61508, A => n14625, ZN => n14624);
   U7679 : AOI22_X1 port map( A1 => n61505, A2 => n706, B1 => n61504, B2 => 
                           n730, ZN => n14625);
   U7680 : OAI221_X1 port map( B1 => n4779, B2 => n61511, C1 => n4755, C2 => 
                           n61508, A => n14550, ZN => n14549);
   U7681 : AOI22_X1 port map( A1 => n61505, A2 => n705, B1 => n61504, B2 => 
                           n729, ZN => n14550);
   U7682 : OAI221_X1 port map( B1 => n4778, B2 => n61511, C1 => n4754, C2 => 
                           n61508, A => n14475, ZN => n14474);
   U7683 : AOI22_X1 port map( A1 => n61505, A2 => n704, B1 => n61504, B2 => 
                           n728, ZN => n14475);
   U7684 : OAI221_X1 port map( B1 => n61860, B2 => n324, C1 => n61857, C2 => 
                           n332, A => n6074, ZN => n6069);
   U7685 : AOI22_X1 port map( A1 => n51775, A2 => n61854, B1 => n51767, B2 => 
                           n61851, ZN => n6074);
   U7686 : OAI221_X1 port map( B1 => n61860, B2 => n323, C1 => n61857, C2 => 
                           n331, A => n5978, ZN => n5975);
   U7687 : AOI22_X1 port map( A1 => n51774, A2 => n61854, B1 => n51766, B2 => 
                           n61851, ZN => n5978);
   U7688 : OAI221_X1 port map( B1 => n61860, B2 => n322, C1 => n61857, C2 => 
                           n330, A => n5903, ZN => n5900);
   U7689 : AOI22_X1 port map( A1 => n51773, A2 => n61854, B1 => n51765, B2 => 
                           n61851, ZN => n5903);
   U7690 : OAI221_X1 port map( B1 => n61860, B2 => n321, C1 => n61857, C2 => 
                           n329, A => n5828, ZN => n5825);
   U7691 : AOI22_X1 port map( A1 => n51772, A2 => n61854, B1 => n51764, B2 => 
                           n61851, ZN => n5828);
   U7692 : OAI221_X1 port map( B1 => n61860, B2 => n320, C1 => n61857, C2 => 
                           n328, A => n5753, ZN => n5750);
   U7693 : AOI22_X1 port map( A1 => n51771, A2 => n61854, B1 => n51763, B2 => 
                           n61851, ZN => n5753);
   U7694 : OAI221_X1 port map( B1 => n61860, B2 => n319, C1 => n61857, C2 => 
                           n327, A => n5678, ZN => n5675);
   U7695 : AOI22_X1 port map( A1 => n51770, A2 => n61854, B1 => n51762, B2 => 
                           n61851, ZN => n5678);
   U7696 : OAI221_X1 port map( B1 => n61860, B2 => n318, C1 => n61857, C2 => 
                           n326, A => n5603, ZN => n5600);
   U7697 : AOI22_X1 port map( A1 => n51769, A2 => n61854, B1 => n51761, B2 => 
                           n61851, ZN => n5603);
   U7698 : OAI221_X1 port map( B1 => n61860, B2 => n317, C1 => n61857, C2 => 
                           n325, A => n5476, ZN => n5469);
   U7699 : AOI22_X1 port map( A1 => n51768, A2 => n61854, B1 => n51760, B2 => 
                           n61851, ZN => n5476);
   U7700 : OAI221_X1 port map( B1 => n61773, B2 => n1073, C1 => n52503, C2 => 
                           n61768, A => n6108, ZN => n6103);
   U7701 : AOI22_X1 port map( A1 => n51671, A2 => n61767, B1 => n51679, B2 => 
                           n61764, ZN => n6108);
   U7702 : OAI221_X1 port map( B1 => n61773, B2 => n1072, C1 => n52502, C2 => 
                           n61768, A => n6002, ZN => n5999);
   U7703 : AOI22_X1 port map( A1 => n51670, A2 => n61767, B1 => n51678, B2 => 
                           n61764, ZN => n6002);
   U7704 : OAI221_X1 port map( B1 => n61773, B2 => n1071, C1 => n52501, C2 => 
                           n61768, A => n5927, ZN => n5924);
   U7705 : AOI22_X1 port map( A1 => n51669, A2 => n61767, B1 => n51677, B2 => 
                           n61764, ZN => n5927);
   U7706 : OAI221_X1 port map( B1 => n61773, B2 => n1070, C1 => n52500, C2 => 
                           n61768, A => n5852, ZN => n5849);
   U7707 : AOI22_X1 port map( A1 => n51668, A2 => n61767, B1 => n51676, B2 => 
                           n61764, ZN => n5852);
   U7708 : OAI221_X1 port map( B1 => n52507, B2 => n61773, C1 => n52499, C2 => 
                           n61768, A => n5777, ZN => n5774);
   U7709 : AOI22_X1 port map( A1 => n51667, A2 => n61767, B1 => n51675, B2 => 
                           n61764, ZN => n5777);
   U7710 : OAI221_X1 port map( B1 => n52506, B2 => n61773, C1 => n52498, C2 => 
                           n61768, A => n5702, ZN => n5699);
   U7711 : AOI22_X1 port map( A1 => n51666, A2 => n61767, B1 => n51674, B2 => 
                           n61764, ZN => n5702);
   U7712 : OAI221_X1 port map( B1 => n52505, B2 => n61773, C1 => n52497, C2 => 
                           n61768, A => n5627, ZN => n5624);
   U7713 : AOI22_X1 port map( A1 => n51665, A2 => n61767, B1 => n51673, B2 => 
                           n61764, ZN => n5627);
   U7714 : OAI221_X1 port map( B1 => n52504, B2 => n61773, C1 => n52496, C2 => 
                           n61768, A => n5541, ZN => n5534);
   U7715 : AOI22_X1 port map( A1 => n51664, A2 => n61767, B1 => n51672, B2 => 
                           n61764, ZN => n5541);
   U7716 : OAI221_X1 port map( B1 => n61701, B2 => n2840, C1 => n61703, C2 => 
                           n2864, A => n7124, ZN => n7117);
   U7717 : AOI222_X1 port map( A1 => n16728, A2 => n62173, B1 => n653, B2 => 
                           n61867, C1 => n16752, C2 => n62171, ZN => n7124);
   U7718 : OAI221_X1 port map( B1 => n61681, B2 => n3908, C1 => n61683, C2 => 
                           n1800, A => n7144, ZN => n7137);
   U7719 : AOI222_X1 port map( A1 => n15525, A2 => n62141, B1 => n15717, B2 => 
                           n61819, C1 => n3112, C2 => n62143, ZN => n7144);
   U7720 : OAI221_X1 port map( B1 => n61701, B2 => n2839, C1 => n61703, C2 => 
                           n2863, A => n7049, ZN => n7042);
   U7721 : AOI222_X1 port map( A1 => n16729, A2 => n62173, B1 => n652, B2 => 
                           n61867, C1 => n16753, C2 => n62171, ZN => n7049);
   U7722 : OAI221_X1 port map( B1 => n61681, B2 => n3907, C1 => n61683, C2 => 
                           n1799, A => n7069, ZN => n7062);
   U7723 : AOI222_X1 port map( A1 => n15526, A2 => n62141, B1 => n15718, B2 => 
                           n61819, C1 => n3111, C2 => n62143, ZN => n7069);
   U7724 : OAI221_X1 port map( B1 => n61701, B2 => n2842, C1 => n61703, C2 => 
                           n2866, A => n7274, ZN => n7267);
   U7725 : AOI222_X1 port map( A1 => n16726, A2 => n62173, B1 => n655, B2 => 
                           n61867, C1 => n16750, C2 => n62171, ZN => n7274);
   U7726 : OAI221_X1 port map( B1 => n61681, B2 => n3910, C1 => n61683, C2 => 
                           n1802, A => n7294, ZN => n7287);
   U7727 : AOI222_X1 port map( A1 => n15523, A2 => n62141, B1 => n15715, B2 => 
                           n61819, C1 => n3114, C2 => n62143, ZN => n7294);
   U7728 : OAI221_X1 port map( B1 => n61701, B2 => n2850, C1 => n61703, C2 => 
                           n2874, A => n7899, ZN => n7891);
   U7729 : AOI222_X1 port map( A1 => n16718, A2 => n62173, B1 => n663, B2 => 
                           n61867, C1 => n16742, C2 => n62171, ZN => n7899);
   U7730 : OAI221_X1 port map( B1 => n61681, B2 => n3918, C1 => n61683, C2 => 
                           n4407, A => n7923, ZN => n7915);
   U7731 : AOI222_X1 port map( A1 => n62141, A2 => n59689, B1 => n15707, B2 => 
                           n61819, C1 => n3122, C2 => n62143, ZN => n7923);
   U7732 : OAI221_X1 port map( B1 => n61701, B2 => n2849, C1 => n61703, C2 => 
                           n2873, A => n7799, ZN => n7792);
   U7733 : AOI222_X1 port map( A1 => n16719, A2 => n62173, B1 => n662, B2 => 
                           n61867, C1 => n16743, C2 => n62171, ZN => n7799);
   U7734 : OAI221_X1 port map( B1 => n61681, B2 => n3917, C1 => n61683, C2 => 
                           n4406, A => n7819, ZN => n7812);
   U7735 : AOI222_X1 port map( A1 => n62141, A2 => n59690, B1 => n15708, B2 => 
                           n61820, C1 => n3121, C2 => n62143, ZN => n7819);
   U7736 : OAI221_X1 port map( B1 => n61701, B2 => n2848, C1 => n61703, C2 => 
                           n2872, A => n7724, ZN => n7717);
   U7737 : AOI222_X1 port map( A1 => n16720, A2 => n62173, B1 => n661, B2 => 
                           n61867, C1 => n16744, C2 => n62171, ZN => n7724);
   U7738 : OAI221_X1 port map( B1 => n61681, B2 => n3916, C1 => n61683, C2 => 
                           n4405, A => n7744, ZN => n7737);
   U7739 : AOI222_X1 port map( A1 => n62141, A2 => n59691, B1 => n15709, B2 => 
                           n61820, C1 => n3120, C2 => n62143, ZN => n7744);
   U7740 : OAI221_X1 port map( B1 => n61701, B2 => n2847, C1 => n61703, C2 => 
                           n2871, A => n7649, ZN => n7642);
   U7741 : AOI222_X1 port map( A1 => n16721, A2 => n62173, B1 => n660, B2 => 
                           n61867, C1 => n16745, C2 => n62171, ZN => n7649);
   U7742 : OAI221_X1 port map( B1 => n61681, B2 => n3915, C1 => n61683, C2 => 
                           n4404, A => n7669, ZN => n7662);
   U7743 : AOI222_X1 port map( A1 => n62141, A2 => n59692, B1 => n15710, B2 => 
                           n61820, C1 => n3119, C2 => n62143, ZN => n7669);
   U7744 : OAI221_X1 port map( B1 => n61701, B2 => n2846, C1 => n61703, C2 => 
                           n2870, A => n7574, ZN => n7567);
   U7745 : AOI222_X1 port map( A1 => n16722, A2 => n62173, B1 => n659, B2 => 
                           n61867, C1 => n16746, C2 => n62171, ZN => n7574);
   U7746 : OAI221_X1 port map( B1 => n61681, B2 => n3914, C1 => n61683, C2 => 
                           n4403, A => n7594, ZN => n7587);
   U7747 : AOI222_X1 port map( A1 => n62141, A2 => n59693, B1 => n15711, B2 => 
                           n61820, C1 => n3118, C2 => n62143, ZN => n7594);
   U7748 : OAI221_X1 port map( B1 => n61701, B2 => n2845, C1 => n61703, C2 => 
                           n2869, A => n7499, ZN => n7492);
   U7749 : AOI222_X1 port map( A1 => n16723, A2 => n62173, B1 => n658, B2 => 
                           n61867, C1 => n16747, C2 => n62171, ZN => n7499);
   U7750 : OAI221_X1 port map( B1 => n61681, B2 => n3913, C1 => n61683, C2 => 
                           n1805, A => n7519, ZN => n7512);
   U7751 : AOI222_X1 port map( A1 => n15520, A2 => n62141, B1 => n15712, B2 => 
                           n61820, C1 => n3117, C2 => n62143, ZN => n7519);
   U7752 : OAI221_X1 port map( B1 => n61701, B2 => n2844, C1 => n61703, C2 => 
                           n2868, A => n7424, ZN => n7417);
   U7753 : AOI222_X1 port map( A1 => n16724, A2 => n62173, B1 => n657, B2 => 
                           n61867, C1 => n16748, C2 => n62171, ZN => n7424);
   U7754 : OAI221_X1 port map( B1 => n61681, B2 => n3912, C1 => n61683, C2 => 
                           n1804, A => n7444, ZN => n7437);
   U7755 : AOI222_X1 port map( A1 => n15521, A2 => n62141, B1 => n15713, B2 => 
                           n61819, C1 => n3116, C2 => n62143, ZN => n7444);
   U7756 : OAI221_X1 port map( B1 => n61701, B2 => n2843, C1 => n61703, C2 => 
                           n2867, A => n7349, ZN => n7342);
   U7757 : AOI222_X1 port map( A1 => n16725, A2 => n62173, B1 => n656, B2 => 
                           n61867, C1 => n16749, C2 => n62171, ZN => n7349);
   U7758 : OAI221_X1 port map( B1 => n61681, B2 => n3911, C1 => n61683, C2 => 
                           n1803, A => n7369, ZN => n7362);
   U7759 : AOI222_X1 port map( A1 => n15522, A2 => n62141, B1 => n15714, B2 => 
                           n61819, C1 => n3115, C2 => n62143, ZN => n7369);
   U7760 : OAI221_X1 port map( B1 => n61701, B2 => n2841, C1 => n61703, C2 => 
                           n2865, A => n7199, ZN => n7192);
   U7761 : AOI222_X1 port map( A1 => n16727, A2 => n62173, B1 => n654, B2 => 
                           n61867, C1 => n16751, C2 => n62171, ZN => n7199);
   U7762 : OAI221_X1 port map( B1 => n61681, B2 => n3909, C1 => n61683, C2 => 
                           n1801, A => n7219, ZN => n7212);
   U7763 : AOI222_X1 port map( A1 => n15524, A2 => n62141, B1 => n15716, B2 => 
                           n61819, C1 => n3113, C2 => n62143, ZN => n7219);
   U7764 : OAI221_X1 port map( B1 => n61788, B2 => n1130, C1 => n61785, C2 => 
                           n1122, A => n6100, ZN => n6093);
   U7765 : AOI222_X1 port map( A1 => n61782, A2 => n4324, B1 => n1518, B2 => 
                           n61779, C1 => n52527, C2 => n61776, ZN => n6100);
   U7766 : OAI221_X1 port map( B1 => n61788, B2 => n1129, C1 => n61785, C2 => 
                           n1121, A => n5996, ZN => n5989);
   U7767 : AOI222_X1 port map( A1 => n61782, A2 => n4323, B1 => n61779, B2 => 
                           n4331, C1 => n52526, C2 => n61776, ZN => n5996);
   U7768 : OAI221_X1 port map( B1 => n61788, B2 => n1128, C1 => n61785, C2 => 
                           n1120, A => n5921, ZN => n5914);
   U7769 : AOI222_X1 port map( A1 => n61782, A2 => n4322, B1 => n61779, B2 => 
                           n4330, C1 => n52525, C2 => n61776, ZN => n5921);
   U7770 : OAI221_X1 port map( B1 => n61788, B2 => n1127, C1 => n61785, C2 => 
                           n1119, A => n5846, ZN => n5839);
   U7771 : AOI222_X1 port map( A1 => n61782, A2 => n4321, B1 => n61779, B2 => 
                           n4329, C1 => n52524, C2 => n61776, ZN => n5846);
   U7772 : OAI221_X1 port map( B1 => n61788, B2 => n1126, C1 => n61785, C2 => 
                           n1118, A => n5771, ZN => n5764);
   U7773 : AOI222_X1 port map( A1 => n61782, A2 => n4320, B1 => n61779, B2 => 
                           n4328, C1 => n52523, C2 => n61776, ZN => n5771);
   U7774 : OAI221_X1 port map( B1 => n61788, B2 => n1125, C1 => n61785, C2 => 
                           n1117, A => n5696, ZN => n5689);
   U7775 : AOI222_X1 port map( A1 => n61782, A2 => n4319, B1 => n61779, B2 => 
                           n4327, C1 => n52522, C2 => n61776, ZN => n5696);
   U7776 : OAI221_X1 port map( B1 => n61788, B2 => n1124, C1 => n61785, C2 => 
                           n1116, A => n5621, ZN => n5614);
   U7777 : AOI222_X1 port map( A1 => n61782, A2 => n4318, B1 => n61779, B2 => 
                           n4326, C1 => n52521, C2 => n61776, ZN => n5621);
   U7778 : OAI221_X1 port map( B1 => n61788, B2 => n1123, C1 => n61785, C2 => 
                           n1115, A => n5528, ZN => n5507);
   U7779 : AOI222_X1 port map( A1 => n61782, A2 => n4317, B1 => n61779, B2 => 
                           n4325, C1 => n52520, C2 => n61776, ZN => n5528);
   U7780 : OAI221_X1 port map( B1 => n2495, B2 => n61799, C1 => n3975, C2 => 
                           n61796, A => n6776, ZN => n6771);
   U7781 : AOI22_X1 port map( A1 => n15435, A2 => n62146, B1 => n15397, B2 => 
                           n62144, ZN => n6776);
   U7782 : OAI221_X1 port map( B1 => n2494, B2 => n61799, C1 => n3974, C2 => 
                           n61796, A => n6701, ZN => n6696);
   U7783 : AOI22_X1 port map( A1 => n15436, A2 => n62146, B1 => n15398, B2 => 
                           n62144, ZN => n6701);
   U7784 : OAI221_X1 port map( B1 => n2493, B2 => n61799, C1 => n3973, C2 => 
                           n61796, A => n6626, ZN => n6621);
   U7785 : AOI22_X1 port map( A1 => n15437, A2 => n62146, B1 => n15399, B2 => 
                           n62144, ZN => n6626);
   U7786 : OAI221_X1 port map( B1 => n2492, B2 => n61799, C1 => n3972, C2 => 
                           n61796, A => n6551, ZN => n6546);
   U7787 : AOI22_X1 port map( A1 => n15438, A2 => n62146, B1 => n15400, B2 => 
                           n62144, ZN => n6551);
   U7788 : OAI221_X1 port map( B1 => n2491, B2 => n61799, C1 => n3971, C2 => 
                           n61796, A => n6476, ZN => n6471);
   U7789 : AOI22_X1 port map( A1 => n15439, A2 => n62146, B1 => n15401, B2 => 
                           n62144, ZN => n6476);
   U7790 : OAI221_X1 port map( B1 => n2490, B2 => n61798, C1 => n3970, C2 => 
                           n61796, A => n6401, ZN => n6396);
   U7791 : AOI22_X1 port map( A1 => n16560, A2 => n62146, B1 => n15697, B2 => 
                           n62144, ZN => n6401);
   U7792 : OAI221_X1 port map( B1 => n2489, B2 => n61798, C1 => n3969, C2 => 
                           n61796, A => n6326, ZN => n6321);
   U7793 : AOI22_X1 port map( A1 => n16561, A2 => n62146, B1 => n15700, B2 => 
                           n62144, ZN => n6326);
   U7794 : OAI221_X1 port map( B1 => n2488, B2 => n61798, C1 => n3968, C2 => 
                           n61796, A => n6251, ZN => n6246);
   U7795 : AOI22_X1 port map( A1 => n16562, A2 => n62146, B1 => n15703, B2 => 
                           n62144, ZN => n6251);
   U7796 : OAI221_X1 port map( B1 => n2487, B2 => n61798, C1 => n3967, C2 => 
                           n61796, A => n6176, ZN => n6171);
   U7797 : AOI22_X1 port map( A1 => n16563, A2 => n62146, B1 => n15706, B2 => 
                           n62144, ZN => n6176);
   U7798 : OAI221_X1 port map( B1 => n2500, B2 => n61799, C1 => n3980, C2 => 
                           n61795, A => n7151, ZN => n7146);
   U7799 : AOI22_X1 port map( A1 => n16558, A2 => n62147, B1 => n15691, B2 => 
                           n62145, ZN => n7151);
   U7800 : OAI221_X1 port map( B1 => n2499, B2 => n61799, C1 => n3979, C2 => 
                           n61795, A => n7076, ZN => n7071);
   U7801 : AOI22_X1 port map( A1 => n16559, A2 => n62147, B1 => n15694, B2 => 
                           n62145, ZN => n7076);
   U7802 : OAI221_X1 port map( B1 => n2497, B2 => n61799, C1 => n3977, C2 => 
                           n61796, A => n6926, ZN => n6921);
   U7803 : AOI22_X1 port map( A1 => n15433, A2 => n62146, B1 => n15395, B2 => 
                           n62144, ZN => n6926);
   U7804 : OAI221_X1 port map( B1 => n2496, B2 => n61799, C1 => n3976, C2 => 
                           n61796, A => n6851, ZN => n6846);
   U7805 : AOI22_X1 port map( A1 => n15434, A2 => n62146, B1 => n15396, B2 => 
                           n62144, ZN => n6851);
   U7806 : OAI221_X1 port map( B1 => n2502, B2 => n61799, C1 => n3982, C2 => 
                           n61795, A => n7301, ZN => n7296);
   U7807 : AOI22_X1 port map( A1 => n16556, A2 => n62147, B1 => n15685, B2 => 
                           n62145, ZN => n7301);
   U7808 : OAI221_X1 port map( B1 => n2510, B2 => n61800, C1 => n3990, C2 => 
                           n61795, A => n7932, ZN => n7926);
   U7809 : AOI22_X1 port map( A1 => n15402, A2 => n62147, B1 => n15380, B2 => 
                           n62145, ZN => n7932);
   U7810 : OAI221_X1 port map( B1 => n2509, B2 => n61800, C1 => n3989, C2 => 
                           n61795, A => n7826, ZN => n7821);
   U7811 : AOI22_X1 port map( A1 => n15427, A2 => n62147, B1 => n15381, B2 => 
                           n62145, ZN => n7826);
   U7812 : OAI221_X1 port map( B1 => n2508, B2 => n61800, C1 => n3988, C2 => 
                           n61795, A => n7751, ZN => n7746);
   U7813 : AOI22_X1 port map( A1 => n15428, A2 => n62147, B1 => n15382, B2 => 
                           n62145, ZN => n7751);
   U7814 : OAI221_X1 port map( B1 => n2507, B2 => n61800, C1 => n3987, C2 => 
                           n61795, A => n7676, ZN => n7671);
   U7815 : AOI22_X1 port map( A1 => n15429, A2 => n62147, B1 => n15383, B2 => 
                           n62145, ZN => n7676);
   U7816 : OAI221_X1 port map( B1 => n2506, B2 => n61800, C1 => n3986, C2 => 
                           n61795, A => n7601, ZN => n7596);
   U7817 : AOI22_X1 port map( A1 => n15430, A2 => n62147, B1 => n15384, B2 => 
                           n62145, ZN => n7601);
   U7818 : OAI221_X1 port map( B1 => n2505, B2 => n61800, C1 => n3985, C2 => 
                           n61795, A => n7526, ZN => n7521);
   U7819 : AOI22_X1 port map( A1 => n15431, A2 => n62147, B1 => n15385, B2 => 
                           n62145, ZN => n7526);
   U7820 : OAI221_X1 port map( B1 => n2504, B2 => n61800, C1 => n3984, C2 => 
                           n61795, A => n7451, ZN => n7446);
   U7821 : AOI22_X1 port map( A1 => n16554, A2 => n62147, B1 => n15726, B2 => 
                           n62145, ZN => n7451);
   U7822 : OAI221_X1 port map( B1 => n2503, B2 => n61799, C1 => n3983, C2 => 
                           n61795, A => n7376, ZN => n7371);
   U7823 : AOI22_X1 port map( A1 => n16555, A2 => n62147, B1 => n15729, B2 => 
                           n62145, ZN => n7376);
   U7824 : OAI221_X1 port map( B1 => n2501, B2 => n61799, C1 => n3981, C2 => 
                           n61795, A => n7226, ZN => n7221);
   U7825 : AOI22_X1 port map( A1 => n16557, A2 => n62147, B1 => n15688, B2 => 
                           n62145, ZN => n7226);
   U7826 : OAI221_X1 port map( B1 => n2498, B2 => n61799, C1 => n3978, C2 => 
                           n61796, A => n7001, ZN => n6996);
   U7827 : AOI22_X1 port map( A1 => n15432, A2 => n62146, B1 => n15386, B2 => 
                           n62144, ZN => n7001);
   U7828 : OAI221_X1 port map( B1 => n9618, B2 => n61911, C1 => n831, C2 => 
                           n59740, A => n6035, ZN => n6026);
   U7829 : AOI222_X1 port map( A1 => n59635, A2 => n111, B1 => n61907, B2 => 
                           n3995, C1 => n52382, C2 => n61903, ZN => n6035);
   U7830 : OAI221_X1 port map( B1 => n9617, B2 => n61911, C1 => n830, C2 => 
                           n59741, A => n5952, ZN => n5945);
   U7831 : AOI222_X1 port map( A1 => n59635, A2 => n110, B1 => n61907, B2 => 
                           n3994, C1 => n52381, C2 => n61903, ZN => n5952);
   U7832 : OAI221_X1 port map( B1 => n9616, B2 => n61911, C1 => n829, C2 => 
                           n59742, A => n5877, ZN => n5870);
   U7833 : AOI222_X1 port map( A1 => n59635, A2 => n109, B1 => n61908, B2 => 
                           n3993, C1 => n52380, C2 => n61903, ZN => n5877);
   U7834 : OAI221_X1 port map( B1 => n9615, B2 => n61911, C1 => n828, C2 => 
                           n59743, A => n5802, ZN => n5795);
   U7835 : AOI222_X1 port map( A1 => n59635, A2 => n108, B1 => n61908, B2 => 
                           n3992, C1 => n52379, C2 => n61903, ZN => n5802);
   U7836 : OAI221_X1 port map( B1 => n9614, B2 => n61911, C1 => n827, C2 => 
                           n59742, A => n5727, ZN => n5720);
   U7837 : AOI222_X1 port map( A1 => n59635, A2 => n107, B1 => n61908, B2 => 
                           n3991, C1 => n52378, C2 => n61903, ZN => n5727);
   U7838 : OAI221_X1 port map( B1 => n9613, B2 => n61911, C1 => n826, C2 => 
                           n59743, A => n5652, ZN => n5645);
   U7839 : AOI222_X1 port map( A1 => n59635, A2 => n106, B1 => n61908, B2 => 
                           n3966, C1 => n52377, C2 => n61903, ZN => n5652);
   U7840 : OAI221_X1 port map( B1 => n9612, B2 => n61911, C1 => n825, C2 => 
                           n59740, A => n5577, ZN => n5570);
   U7841 : AOI222_X1 port map( A1 => n59635, A2 => n105, B1 => n61908, B2 => 
                           n3965, C1 => n52376, C2 => n61903, ZN => n5577);
   U7842 : OAI221_X1 port map( B1 => n9611, B2 => n61911, C1 => n824, C2 => 
                           n59741, A => n5420, ZN => n5401);
   U7843 : AOI222_X1 port map( A1 => n59635, A2 => n104, B1 => n61908, B2 => 
                           n3964, C1 => n52375, C2 => n61903, ZN => n5420);
   U7844 : OAI221_X1 port map( B1 => n15177, B2 => n61324, C1 => n15209, C2 => 
                           n61321, A => n8596, ZN => n8589);
   U7845 : AOI222_X1 port map( A1 => n61318, A2 => n52518, B1 => n61313, B2 => 
                           n52526, C1 => n61310, C2 => n52534, ZN => n8596);
   U7846 : OAI221_X1 port map( B1 => n15176, B2 => n61324, C1 => n15208, C2 => 
                           n61321, A => n8521, ZN => n8514);
   U7847 : AOI222_X1 port map( A1 => n61318, A2 => n52517, B1 => n61313, B2 => 
                           n52525, C1 => n61310, C2 => n52533, ZN => n8521);
   U7848 : OAI221_X1 port map( B1 => n15175, B2 => n61324, C1 => n15207, C2 => 
                           n61321, A => n8446, ZN => n8439);
   U7849 : AOI222_X1 port map( A1 => n61318, A2 => n52516, B1 => n61313, B2 => 
                           n52524, C1 => n61310, C2 => n52532, ZN => n8446);
   U7850 : OAI221_X1 port map( B1 => n15174, B2 => n61324, C1 => n15206, C2 => 
                           n61321, A => n8371, ZN => n8364);
   U7851 : AOI222_X1 port map( A1 => n61318, A2 => n52515, B1 => n61313, B2 => 
                           n52523, C1 => n61310, C2 => n52531, ZN => n8371);
   U7852 : OAI221_X1 port map( B1 => n15173, B2 => n61324, C1 => n15205, C2 => 
                           n61321, A => n8296, ZN => n8289);
   U7853 : AOI222_X1 port map( A1 => n61318, A2 => n52514, B1 => n61313, B2 => 
                           n52522, C1 => n61310, C2 => n52530, ZN => n8296);
   U7854 : OAI221_X1 port map( B1 => n15172, B2 => n61324, C1 => n15204, C2 => 
                           n61321, A => n8221, ZN => n8214);
   U7855 : AOI222_X1 port map( A1 => n61318, A2 => n52513, B1 => n61313, B2 => 
                           n52521, C1 => n61310, C2 => n52529, ZN => n8221);
   U7856 : OAI221_X1 port map( B1 => n15171, B2 => n61324, C1 => n15203, C2 => 
                           n61321, A => n8126, ZN => n8105);
   U7857 : AOI222_X1 port map( A1 => n61318, A2 => n52512, B1 => n61313, B2 => 
                           n52520, C1 => n61310, C2 => n52528, ZN => n8126);
   U7858 : OAI221_X1 port map( B1 => n51, B2 => n61579, C1 => n43, C2 => n61576
                           , A => n8627, ZN => n8620);
   U7859 : AOI222_X1 port map( A1 => n61573, A2 => n52382, B1 => n61568, B2 => 
                           n52390, C1 => n61565, C2 => n783, ZN => n8627);
   U7860 : OAI221_X1 port map( B1 => n4131, B2 => n61630, C1 => n4123, C2 => 
                           n61627, A => n8619, ZN => n8612);
   U7861 : AOI222_X1 port map( A1 => n61624, A2 => n51607, B1 => n61619, B2 => 
                           n855, C1 => n61616, C2 => n863, ZN => n8619);
   U7862 : OAI221_X1 port map( B1 => n1250, B2 => n61375, C1 => n1242, C2 => 
                           n61372, A => n8663, ZN => n8656);
   U7863 : AOI222_X1 port map( A1 => n61369, A2 => n52591, B1 => n61364, B2 => 
                           n52599, C1 => n61361, C2 => n52607, ZN => n8663);
   U7864 : OAI221_X1 port map( B1 => n284, B2 => n61426, C1 => n276, C2 => 
                           n61423, A => n8655, ZN => n8648);
   U7865 : AOI222_X1 port map( A1 => n61420, A2 => n52663, B1 => n61415, B2 => 
                           n4035, C1 => n61412, C2 => n4043, ZN => n8655);
   U7866 : OAI221_X1 port map( B1 => n283, B2 => n61426, C1 => n275, C2 => 
                           n61423, A => n8580, ZN => n8573);
   U7867 : AOI222_X1 port map( A1 => n61420, A2 => n52662, B1 => n61415, B2 => 
                           n4034, C1 => n61412, C2 => n4042, ZN => n8580);
   U7868 : OAI221_X1 port map( B1 => n282, B2 => n61426, C1 => n274, C2 => 
                           n61423, A => n8505, ZN => n8498);
   U7869 : AOI222_X1 port map( A1 => n61420, A2 => n52661, B1 => n61415, B2 => 
                           n4033, C1 => n61412, C2 => n4041, ZN => n8505);
   U7870 : OAI221_X1 port map( B1 => n281, B2 => n61426, C1 => n273, C2 => 
                           n61423, A => n8430, ZN => n8423);
   U7871 : AOI222_X1 port map( A1 => n61420, A2 => n52660, B1 => n61415, B2 => 
                           n4032, C1 => n61412, C2 => n4040, ZN => n8430);
   U7872 : OAI221_X1 port map( B1 => n280, B2 => n61426, C1 => n272, C2 => 
                           n61423, A => n8355, ZN => n8348);
   U7873 : AOI222_X1 port map( A1 => n61420, A2 => n52659, B1 => n61415, B2 => 
                           n4031, C1 => n61412, C2 => n4039, ZN => n8355);
   U7874 : OAI221_X1 port map( B1 => n279, B2 => n61426, C1 => n271, C2 => 
                           n61423, A => n8280, ZN => n8273);
   U7875 : AOI222_X1 port map( A1 => n61420, A2 => n52658, B1 => n61415, B2 => 
                           n4030, C1 => n61412, C2 => n4038, ZN => n8280);
   U7876 : OAI221_X1 port map( B1 => n278, B2 => n61426, C1 => n270, C2 => 
                           n61423, A => n8205, ZN => n8198);
   U7877 : AOI222_X1 port map( A1 => n61420, A2 => n52657, B1 => n61415, B2 => 
                           n4029, C1 => n61412, C2 => n4037, ZN => n8205);
   U7878 : OAI221_X1 port map( B1 => n277, B2 => n61426, C1 => n269, C2 => 
                           n61423, A => n8076, ZN => n8055);
   U7879 : AOI222_X1 port map( A1 => n61420, A2 => n52656, B1 => n61415, B2 => 
                           n4028, C1 => n61412, C2 => n4036, ZN => n8076);
   U7880 : OAI221_X1 port map( B1 => n4235, B2 => n61528, C1 => n4227, C2 => 
                           n61525, A => n8635, ZN => n8628);
   U7881 : AOI222_X1 port map( A1 => n61522, A2 => n52315, B1 => n61517, B2 => 
                           n52323, C1 => n61514, C2 => n52331, ZN => n8635);
   U7882 : OAI221_X1 port map( B1 => n1114, B2 => n61324, C1 => n15210, C2 => 
                           n61321, A => n8671, ZN => n8664);
   U7883 : AOI222_X1 port map( A1 => n61318, A2 => n52519, B1 => n61313, B2 => 
                           n52527, C1 => n61310, C2 => n52535, ZN => n8671);
   U7884 : OAI221_X1 port map( B1 => n4234, B2 => n61528, C1 => n4226, C2 => 
                           n61525, A => n8560, ZN => n8553);
   U7885 : AOI222_X1 port map( A1 => n61522, A2 => n52314, B1 => n61517, B2 => 
                           n52322, C1 => n61514, C2 => n52330, ZN => n8560);
   U7886 : OAI221_X1 port map( B1 => n50, B2 => n61579, C1 => n42, C2 => n61576
                           , A => n8552, ZN => n8545);
   U7887 : AOI222_X1 port map( A1 => n61573, A2 => n52381, B1 => n61568, B2 => 
                           n52389, C1 => n61565, C2 => n782, ZN => n8552);
   U7888 : OAI221_X1 port map( B1 => n4130, B2 => n61630, C1 => n4122, C2 => 
                           n61627, A => n8544, ZN => n8537);
   U7889 : AOI222_X1 port map( A1 => n61624, A2 => n51606, B1 => n61619, B2 => 
                           n854, C1 => n61616, C2 => n862, ZN => n8544);
   U7890 : OAI221_X1 port map( B1 => n1249, B2 => n61375, C1 => n1241, C2 => 
                           n61372, A => n8588, ZN => n8581);
   U7891 : AOI222_X1 port map( A1 => n61369, A2 => n52590, B1 => n61364, B2 => 
                           n52598, C1 => n61361, C2 => n52606, ZN => n8588);
   U7892 : OAI221_X1 port map( B1 => n4233, B2 => n61528, C1 => n4225, C2 => 
                           n61525, A => n8485, ZN => n8478);
   U7893 : AOI222_X1 port map( A1 => n61522, A2 => n52313, B1 => n61517, B2 => 
                           n52321, C1 => n61514, C2 => n52329, ZN => n8485);
   U7894 : OAI221_X1 port map( B1 => n49, B2 => n61579, C1 => n41, C2 => n61576
                           , A => n8477, ZN => n8470);
   U7895 : AOI222_X1 port map( A1 => n61573, A2 => n52380, B1 => n61568, B2 => 
                           n52388, C1 => n61565, C2 => n781, ZN => n8477);
   U7896 : OAI221_X1 port map( B1 => n4129, B2 => n61630, C1 => n4121, C2 => 
                           n61627, A => n8469, ZN => n8462);
   U7897 : AOI222_X1 port map( A1 => n61624, A2 => n51605, B1 => n61619, B2 => 
                           n853, C1 => n61616, C2 => n861, ZN => n8469);
   U7898 : OAI221_X1 port map( B1 => n1248, B2 => n61375, C1 => n1240, C2 => 
                           n61372, A => n8513, ZN => n8506);
   U7899 : AOI222_X1 port map( A1 => n61369, A2 => n52589, B1 => n61364, B2 => 
                           n52597, C1 => n61361, C2 => n52605, ZN => n8513);
   U7900 : OAI221_X1 port map( B1 => n4232, B2 => n61528, C1 => n4224, C2 => 
                           n61525, A => n8410, ZN => n8403);
   U7901 : AOI222_X1 port map( A1 => n61522, A2 => n52312, B1 => n61517, B2 => 
                           n52320, C1 => n61514, C2 => n52328, ZN => n8410);
   U7902 : OAI221_X1 port map( B1 => n48, B2 => n61579, C1 => n40, C2 => n61576
                           , A => n8402, ZN => n8395);
   U7903 : AOI222_X1 port map( A1 => n61573, A2 => n52379, B1 => n61568, B2 => 
                           n52387, C1 => n61565, C2 => n780, ZN => n8402);
   U7904 : OAI221_X1 port map( B1 => n4128, B2 => n61630, C1 => n4120, C2 => 
                           n61627, A => n8394, ZN => n8387);
   U7905 : AOI222_X1 port map( A1 => n61624, A2 => n51604, B1 => n61619, B2 => 
                           n852, C1 => n61616, C2 => n860, ZN => n8394);
   U7906 : OAI221_X1 port map( B1 => n1247, B2 => n61375, C1 => n1239, C2 => 
                           n61372, A => n8438, ZN => n8431);
   U7907 : AOI222_X1 port map( A1 => n61369, A2 => n52588, B1 => n61364, B2 => 
                           n52596, C1 => n61361, C2 => n52604, ZN => n8438);
   U7908 : OAI221_X1 port map( B1 => n4231, B2 => n61528, C1 => n4223, C2 => 
                           n61525, A => n8335, ZN => n8328);
   U7909 : AOI222_X1 port map( A1 => n61522, A2 => n52311, B1 => n61517, B2 => 
                           n52319, C1 => n61514, C2 => n52327, ZN => n8335);
   U7910 : OAI221_X1 port map( B1 => n47, B2 => n61579, C1 => n39, C2 => n61576
                           , A => n8327, ZN => n8320);
   U7911 : AOI222_X1 port map( A1 => n61573, A2 => n52378, B1 => n61568, B2 => 
                           n52386, C1 => n61565, C2 => n779, ZN => n8327);
   U7912 : OAI221_X1 port map( B1 => n4127, B2 => n61630, C1 => n4119, C2 => 
                           n61627, A => n8319, ZN => n8312);
   U7913 : AOI222_X1 port map( A1 => n61624, A2 => n51603, B1 => n61619, B2 => 
                           n851, C1 => n61616, C2 => n859, ZN => n8319);
   U7914 : OAI221_X1 port map( B1 => n1246, B2 => n61375, C1 => n1238, C2 => 
                           n61372, A => n8363, ZN => n8356);
   U7915 : AOI222_X1 port map( A1 => n61369, A2 => n52587, B1 => n61364, B2 => 
                           n52595, C1 => n61361, C2 => n52603, ZN => n8363);
   U7916 : OAI221_X1 port map( B1 => n4230, B2 => n61528, C1 => n4222, C2 => 
                           n61525, A => n8260, ZN => n8253);
   U7917 : AOI222_X1 port map( A1 => n61522, A2 => n52310, B1 => n61517, B2 => 
                           n52318, C1 => n61514, C2 => n52326, ZN => n8260);
   U7918 : OAI221_X1 port map( B1 => n46, B2 => n61579, C1 => n38, C2 => n61576
                           , A => n8252, ZN => n8245);
   U7919 : AOI222_X1 port map( A1 => n61573, A2 => n52377, B1 => n61568, B2 => 
                           n52385, C1 => n61565, C2 => n778, ZN => n8252);
   U7920 : OAI221_X1 port map( B1 => n4126, B2 => n61630, C1 => n4118, C2 => 
                           n61627, A => n8244, ZN => n8237);
   U7921 : AOI222_X1 port map( A1 => n61624, A2 => n51602, B1 => n61619, B2 => 
                           n850, C1 => n61616, C2 => n858, ZN => n8244);
   U7922 : OAI221_X1 port map( B1 => n1245, B2 => n61375, C1 => n1237, C2 => 
                           n61372, A => n8288, ZN => n8281);
   U7923 : AOI222_X1 port map( A1 => n61369, A2 => n52586, B1 => n61364, B2 => 
                           n52594, C1 => n61361, C2 => n52602, ZN => n8288);
   U7924 : OAI221_X1 port map( B1 => n4229, B2 => n61528, C1 => n4221, C2 => 
                           n61525, A => n8185, ZN => n8178);
   U7925 : AOI222_X1 port map( A1 => n61522, A2 => n52309, B1 => n61517, B2 => 
                           n52317, C1 => n61514, C2 => n52325, ZN => n8185);
   U7926 : OAI221_X1 port map( B1 => n45, B2 => n61579, C1 => n37, C2 => n61576
                           , A => n8177, ZN => n8170);
   U7927 : AOI222_X1 port map( A1 => n61573, A2 => n52376, B1 => n61568, B2 => 
                           n52384, C1 => n61565, C2 => n777, ZN => n8177);
   U7928 : OAI221_X1 port map( B1 => n4125, B2 => n61630, C1 => n4117, C2 => 
                           n61627, A => n8169, ZN => n8162);
   U7929 : AOI222_X1 port map( A1 => n61624, A2 => n51601, B1 => n61619, B2 => 
                           n849, C1 => n61616, C2 => n857, ZN => n8169);
   U7930 : OAI221_X1 port map( B1 => n1244, B2 => n61375, C1 => n1236, C2 => 
                           n61372, A => n8213, ZN => n8206);
   U7931 : AOI222_X1 port map( A1 => n61369, A2 => n52585, B1 => n61364, B2 => 
                           n52593, C1 => n61361, C2 => n52601, ZN => n8213);
   U7932 : OAI221_X1 port map( B1 => n4228, B2 => n61528, C1 => n4220, C2 => 
                           n61525, A => n8022, ZN => n8001);
   U7933 : AOI222_X1 port map( A1 => n61522, A2 => n52308, B1 => n61517, B2 => 
                           n52316, C1 => n61514, C2 => n52324, ZN => n8022);
   U7934 : OAI221_X1 port map( B1 => n44, B2 => n61579, C1 => n36, C2 => n61576
                           , A => n7997, ZN => n7976);
   U7935 : AOI222_X1 port map( A1 => n61573, A2 => n52375, B1 => n61568, B2 => 
                           n52383, C1 => n61565, C2 => n776, ZN => n7997);
   U7936 : OAI221_X1 port map( B1 => n4124, B2 => n61630, C1 => n4116, C2 => 
                           n61627, A => n7972, ZN => n7951);
   U7937 : AOI222_X1 port map( A1 => n61624, A2 => n51600, B1 => n61619, B2 => 
                           n848, C1 => n61616, C2 => n856, ZN => n7972);
   U7938 : OAI221_X1 port map( B1 => n1243, B2 => n61375, C1 => n1235, C2 => 
                           n61372, A => n8101, ZN => n8080);
   U7939 : AOI222_X1 port map( A1 => n61369, A2 => n52584, B1 => n61364, B2 => 
                           n52592, C1 => n61361, C2 => n52600, ZN => n8101);
   U7940 : OAI221_X1 port map( B1 => n61889, B2 => n3217, C1 => n61886, C2 => 
                           n3241, A => n6741, ZN => n6734);
   U7941 : AOI222_X1 port map( A1 => n16497, A2 => n62162, B1 => n62160, B2 => 
                           n4938, C1 => n16651, C2 => n62158, ZN => n6741);
   U7942 : OAI221_X1 port map( B1 => n6059, B2 => n2787, C1 => n61704, C2 => 
                           n2859, A => n6749, ZN => n6742);
   U7943 : AOI222_X1 port map( A1 => n16733, A2 => n62172, B1 => n648, B2 => 
                           n61868, C1 => n16757, C2 => n62170, ZN => n6749);
   U7944 : OAI221_X1 port map( B1 => n61955, B2 => n4656, C1 => n61952, C2 => 
                           n4680, A => n6725, ZN => n6718);
   U7945 : AOI222_X1 port map( A1 => n62180, A2 => n4632, B1 => n61937, B2 => 
                           n4440, C1 => n16802, C2 => n62176, ZN => n6725);
   U7946 : OAI221_X1 port map( B1 => n6089, B2 => n3903, C1 => n61684, C2 => 
                           n1795, A => n6769, ZN => n6762);
   U7947 : AOI222_X1 port map( A1 => n15530, A2 => n62140, B1 => n15722, B2 => 
                           n61819, C1 => n3107, C2 => n62142, ZN => n6769);
   U7948 : OAI221_X1 port map( B1 => n61889, B2 => n3216, C1 => n61886, C2 => 
                           n3240, A => n6666, ZN => n6659);
   U7949 : AOI222_X1 port map( A1 => n16498, A2 => n62162, B1 => n62160, B2 => 
                           n4937, C1 => n16652, C2 => n62158, ZN => n6666);
   U7950 : OAI221_X1 port map( B1 => n6059, B2 => n2786, C1 => n61704, C2 => 
                           n2858, A => n6674, ZN => n6667);
   U7951 : AOI222_X1 port map( A1 => n16734, A2 => n62172, B1 => n647, B2 => 
                           n61868, C1 => n16758, C2 => n62170, ZN => n6674);
   U7952 : OAI221_X1 port map( B1 => n61955, B2 => n4655, C1 => n61952, C2 => 
                           n4679, A => n6650, ZN => n6643);
   U7953 : AOI222_X1 port map( A1 => n62180, A2 => n4631, B1 => n61937, B2 => 
                           n4439, C1 => n16803, C2 => n62176, ZN => n6650);
   U7954 : OAI221_X1 port map( B1 => n6089, B2 => n3902, C1 => n61684, C2 => 
                           n1794, A => n6694, ZN => n6687);
   U7955 : AOI222_X1 port map( A1 => n15531, A2 => n62140, B1 => n15723, B2 => 
                           n61819, C1 => n3106, C2 => n62142, ZN => n6694);
   U7956 : OAI221_X1 port map( B1 => n61889, B2 => n3215, C1 => n61886, C2 => 
                           n3239, A => n6591, ZN => n6584);
   U7957 : AOI222_X1 port map( A1 => n16499, A2 => n62162, B1 => n62160, B2 => 
                           n4936, C1 => n16653, C2 => n62158, ZN => n6591);
   U7958 : OAI221_X1 port map( B1 => n6059, B2 => n2785, C1 => n61704, C2 => 
                           n2857, A => n6599, ZN => n6592);
   U7959 : AOI222_X1 port map( A1 => n16735, A2 => n62172, B1 => n646, B2 => 
                           n61868, C1 => n16759, C2 => n62170, ZN => n6599);
   U7960 : OAI221_X1 port map( B1 => n61955, B2 => n4654, C1 => n61952, C2 => 
                           n4678, A => n6575, ZN => n6568);
   U7961 : AOI222_X1 port map( A1 => n62180, A2 => n4630, B1 => n61937, B2 => 
                           n4438, C1 => n16804, C2 => n62176, ZN => n6575);
   U7962 : OAI221_X1 port map( B1 => n6089, B2 => n3901, C1 => n61684, C2 => 
                           n1793, A => n6619, ZN => n6612);
   U7963 : AOI222_X1 port map( A1 => n15532, A2 => n62140, B1 => n61821, B2 => 
                           n59730, C1 => n3105, C2 => n62142, ZN => n6619);
   U7964 : OAI221_X1 port map( B1 => n61889, B2 => n3214, C1 => n61886, C2 => 
                           n3238, A => n6516, ZN => n6509);
   U7965 : AOI222_X1 port map( A1 => n16500, A2 => n62162, B1 => n62160, B2 => 
                           n4935, C1 => n16654, C2 => n62158, ZN => n6516);
   U7966 : OAI221_X1 port map( B1 => n6059, B2 => n2784, C1 => n61704, C2 => 
                           n2856, A => n6524, ZN => n6517);
   U7967 : AOI222_X1 port map( A1 => n16736, A2 => n62172, B1 => n645, B2 => 
                           n61868, C1 => n16760, C2 => n62170, ZN => n6524);
   U7968 : OAI221_X1 port map( B1 => n61955, B2 => n4653, C1 => n61952, C2 => 
                           n4677, A => n6500, ZN => n6493);
   U7969 : AOI222_X1 port map( A1 => n62180, A2 => n4629, B1 => n61937, B2 => 
                           n4437, C1 => n16805, C2 => n62176, ZN => n6500);
   U7970 : OAI221_X1 port map( B1 => n6089, B2 => n3900, C1 => n61684, C2 => 
                           n1792, A => n6544, ZN => n6537);
   U7971 : AOI222_X1 port map( A1 => n15533, A2 => n62140, B1 => n61821, B2 => 
                           n59731, C1 => n3104, C2 => n62142, ZN => n6544);
   U7972 : OAI221_X1 port map( B1 => n61889, B2 => n3213, C1 => n61886, C2 => 
                           n3237, A => n6441, ZN => n6434);
   U7973 : AOI222_X1 port map( A1 => n16501, A2 => n62162, B1 => n62160, B2 => 
                           n4934, C1 => n16655, C2 => n62158, ZN => n6441);
   U7974 : OAI221_X1 port map( B1 => n6059, B2 => n2783, C1 => n61704, C2 => 
                           n2855, A => n6449, ZN => n6442);
   U7975 : AOI222_X1 port map( A1 => n16737, A2 => n62172, B1 => n644, B2 => 
                           n61868, C1 => n16761, C2 => n62170, ZN => n6449);
   U7976 : OAI221_X1 port map( B1 => n61955, B2 => n4652, C1 => n61952, C2 => 
                           n4676, A => n6425, ZN => n6418);
   U7977 : AOI222_X1 port map( A1 => n62180, A2 => n4628, B1 => n61937, B2 => 
                           n4436, C1 => n16806, C2 => n62176, ZN => n6425);
   U7978 : OAI221_X1 port map( B1 => n6089, B2 => n3899, C1 => n61684, C2 => 
                           n1791, A => n6469, ZN => n6462);
   U7979 : AOI222_X1 port map( A1 => n15534, A2 => n62140, B1 => n61821, B2 => 
                           n59732, C1 => n3103, C2 => n62142, ZN => n6469);
   U7980 : OAI221_X1 port map( B1 => n61889, B2 => n3212, C1 => n61886, C2 => 
                           n3236, A => n6366, ZN => n6359);
   U7981 : AOI222_X1 port map( A1 => n16502, A2 => n62162, B1 => n62160, B2 => 
                           n4933, C1 => n16656, C2 => n62158, ZN => n6366);
   U7982 : OAI221_X1 port map( B1 => n6059, B2 => n2782, C1 => n61704, C2 => 
                           n2854, A => n6374, ZN => n6367);
   U7983 : AOI222_X1 port map( A1 => n16738, A2 => n62172, B1 => n643, B2 => 
                           n61868, C1 => n16762, C2 => n62170, ZN => n6374);
   U7984 : OAI221_X1 port map( B1 => n61955, B2 => n4651, C1 => n61952, C2 => 
                           n4675, A => n6350, ZN => n6343);
   U7985 : AOI222_X1 port map( A1 => n62180, A2 => n4627, B1 => n61936, B2 => 
                           n4435, C1 => n16795, C2 => n62176, ZN => n6350);
   U7986 : OAI221_X1 port map( B1 => n6089, B2 => n3898, C1 => n61684, C2 => 
                           n1790, A => n6394, ZN => n6387);
   U7987 : AOI222_X1 port map( A1 => n15535, A2 => n62140, B1 => n61821, B2 => 
                           n59733, C1 => n3102, C2 => n62142, ZN => n6394);
   U7988 : OAI221_X1 port map( B1 => n61889, B2 => n3211, C1 => n61886, C2 => 
                           n3235, A => n6291, ZN => n6284);
   U7989 : AOI222_X1 port map( A1 => n16503, A2 => n62162, B1 => n62160, B2 => 
                           n4932, C1 => n16657, C2 => n62158, ZN => n6291);
   U7990 : OAI221_X1 port map( B1 => n6059, B2 => n2781, C1 => n61704, C2 => 
                           n2853, A => n6299, ZN => n6292);
   U7991 : AOI222_X1 port map( A1 => n16739, A2 => n62172, B1 => n642, B2 => 
                           n61868, C1 => n16763, C2 => n62170, ZN => n6299);
   U7992 : OAI221_X1 port map( B1 => n61955, B2 => n4650, C1 => n61952, C2 => 
                           n4674, A => n6275, ZN => n6268);
   U7993 : AOI222_X1 port map( A1 => n62180, A2 => n4626, B1 => n61936, B2 => 
                           n4434, C1 => n16796, C2 => n62176, ZN => n6275);
   U7994 : OAI221_X1 port map( B1 => n6089, B2 => n3897, C1 => n61684, C2 => 
                           n1789, A => n6319, ZN => n6312);
   U7995 : AOI222_X1 port map( A1 => n15536, A2 => n62140, B1 => n61821, B2 => 
                           n59734, C1 => n3101, C2 => n62142, ZN => n6319);
   U7996 : OAI221_X1 port map( B1 => n61889, B2 => n3210, C1 => n61886, C2 => 
                           n3234, A => n6216, ZN => n6209);
   U7997 : AOI222_X1 port map( A1 => n16504, A2 => n62162, B1 => n62160, B2 => 
                           n4931, C1 => n16658, C2 => n62158, ZN => n6216);
   U7998 : OAI221_X1 port map( B1 => n6059, B2 => n2780, C1 => n61704, C2 => 
                           n2852, A => n6224, ZN => n6217);
   U7999 : AOI222_X1 port map( A1 => n16740, A2 => n62172, B1 => n641, B2 => 
                           n61868, C1 => n16764, C2 => n62170, ZN => n6224);
   U8000 : OAI221_X1 port map( B1 => n61955, B2 => n4649, C1 => n61952, C2 => 
                           n4673, A => n6200, ZN => n6193);
   U8001 : AOI222_X1 port map( A1 => n62180, A2 => n4625, B1 => n61936, B2 => 
                           n4433, C1 => n16797, C2 => n62176, ZN => n6200);
   U8002 : OAI221_X1 port map( B1 => n6089, B2 => n3896, C1 => n61684, C2 => 
                           n1788, A => n6244, ZN => n6237);
   U8003 : AOI222_X1 port map( A1 => n15537, A2 => n62140, B1 => n61821, B2 => 
                           n59735, C1 => n3100, C2 => n62142, ZN => n6244);
   U8004 : OAI221_X1 port map( B1 => n61889, B2 => n3209, C1 => n61886, C2 => 
                           n3233, A => n6141, ZN => n6134);
   U8005 : AOI222_X1 port map( A1 => n16505, A2 => n62162, B1 => n62160, B2 => 
                           n4930, C1 => n16659, C2 => n62158, ZN => n6141);
   U8006 : OAI221_X1 port map( B1 => n6059, B2 => n2779, C1 => n61704, C2 => 
                           n2851, A => n6149, ZN => n6142);
   U8007 : AOI222_X1 port map( A1 => n16741, A2 => n62172, B1 => n640, B2 => 
                           n61868, C1 => n16765, C2 => n62170, ZN => n6149);
   U8008 : OAI221_X1 port map( B1 => n61955, B2 => n4648, C1 => n61952, C2 => 
                           n4672, A => n6125, ZN => n6118);
   U8009 : AOI222_X1 port map( A1 => n62180, A2 => n4624, B1 => n61936, B2 => 
                           n4432, C1 => n16798, C2 => n62176, ZN => n6125);
   U8010 : OAI221_X1 port map( B1 => n6089, B2 => n3895, C1 => n61684, C2 => 
                           n1787, A => n6169, ZN => n6162);
   U8011 : AOI222_X1 port map( A1 => n15538, A2 => n62140, B1 => n61821, B2 => 
                           n59736, C1 => n3099, C2 => n62142, ZN => n6169);
   U8012 : OAI221_X1 port map( B1 => n61888, B2 => n3222, C1 => n61885, C2 => 
                           n3246, A => n7116, ZN => n7109);
   U8013 : AOI222_X1 port map( A1 => n16492, A2 => n62163, B1 => n62161, B2 => 
                           n4943, C1 => n16646, C2 => n62159, ZN => n7116);
   U8014 : OAI221_X1 port map( B1 => n61954, B2 => n4661, C1 => n61951, C2 => 
                           n4685, A => n7100, ZN => n7093);
   U8015 : AOI222_X1 port map( A1 => n62181, A2 => n4637, B1 => n61937, B2 => 
                           n4445, C1 => n16807, C2 => n62177, ZN => n7100);
   U8016 : OAI221_X1 port map( B1 => n61888, B2 => n3221, C1 => n61885, C2 => 
                           n3245, A => n7041, ZN => n7034);
   U8017 : AOI222_X1 port map( A1 => n16493, A2 => n62163, B1 => n62161, B2 => 
                           n4942, C1 => n16647, C2 => n62159, ZN => n7041);
   U8018 : OAI221_X1 port map( B1 => n61954, B2 => n4660, C1 => n61951, C2 => 
                           n4684, A => n7025, ZN => n7018);
   U8019 : AOI222_X1 port map( A1 => n62181, A2 => n4636, B1 => n61937, B2 => 
                           n4444, C1 => n16808, C2 => n62177, ZN => n7025);
   U8020 : OAI221_X1 port map( B1 => n61889, B2 => n3219, C1 => n61886, C2 => 
                           n3243, A => n6891, ZN => n6884);
   U8021 : AOI222_X1 port map( A1 => n16495, A2 => n62162, B1 => n62160, B2 => 
                           n4940, C1 => n16649, C2 => n62158, ZN => n6891);
   U8022 : OAI221_X1 port map( B1 => n6059, B2 => n2789, C1 => n61704, C2 => 
                           n2861, A => n6899, ZN => n6892);
   U8023 : AOI222_X1 port map( A1 => n16731, A2 => n62172, B1 => n650, B2 => 
                           n61868, C1 => n16755, C2 => n62170, ZN => n6899);
   U8024 : OAI221_X1 port map( B1 => n61955, B2 => n4658, C1 => n61952, C2 => 
                           n4682, A => n6875, ZN => n6868);
   U8025 : AOI222_X1 port map( A1 => n62180, A2 => n4634, B1 => n61937, B2 => 
                           n4442, C1 => n16809, C2 => n62176, ZN => n6875);
   U8026 : OAI221_X1 port map( B1 => n6089, B2 => n3905, C1 => n61684, C2 => 
                           n1797, A => n6919, ZN => n6912);
   U8027 : AOI222_X1 port map( A1 => n15528, A2 => n62140, B1 => n15720, B2 => 
                           n61819, C1 => n3109, C2 => n62142, ZN => n6919);
   U8028 : OAI221_X1 port map( B1 => n61889, B2 => n3218, C1 => n61886, C2 => 
                           n3242, A => n6816, ZN => n6809);
   U8029 : AOI222_X1 port map( A1 => n16496, A2 => n62162, B1 => n62160, B2 => 
                           n4939, C1 => n16650, C2 => n62158, ZN => n6816);
   U8030 : OAI221_X1 port map( B1 => n6059, B2 => n2788, C1 => n61704, C2 => 
                           n2860, A => n6824, ZN => n6817);
   U8031 : AOI222_X1 port map( A1 => n16732, A2 => n62172, B1 => n649, B2 => 
                           n61868, C1 => n16756, C2 => n62170, ZN => n6824);
   U8032 : OAI221_X1 port map( B1 => n61955, B2 => n4657, C1 => n61952, C2 => 
                           n4681, A => n6800, ZN => n6793);
   U8033 : AOI222_X1 port map( A1 => n62180, A2 => n4633, B1 => n61937, B2 => 
                           n4441, C1 => n16810, C2 => n62176, ZN => n6800);
   U8034 : OAI221_X1 port map( B1 => n6089, B2 => n3904, C1 => n61684, C2 => 
                           n1796, A => n6844, ZN => n6837);
   U8035 : AOI222_X1 port map( A1 => n15529, A2 => n62140, B1 => n15721, B2 => 
                           n61819, C1 => n3108, C2 => n62142, ZN => n6844);
   U8036 : OAI221_X1 port map( B1 => n61888, B2 => n3224, C1 => n61885, C2 => 
                           n3248, A => n7266, ZN => n7259);
   U8037 : AOI222_X1 port map( A1 => n16490, A2 => n62163, B1 => n62161, B2 => 
                           n4945, C1 => n16644, C2 => n62159, ZN => n7266);
   U8038 : OAI221_X1 port map( B1 => n61954, B2 => n4663, C1 => n61951, C2 => 
                           n4687, A => n7250, ZN => n7243);
   U8039 : AOI222_X1 port map( A1 => n62181, A2 => n4639, B1 => n61937, B2 => 
                           n4447, C1 => n16794, C2 => n62177, ZN => n7250);
   U8040 : OAI221_X1 port map( B1 => n61888, B2 => n3232, C1 => n61885, C2 => 
                           n3256, A => n7888, ZN => n7878);
   U8041 : AOI222_X1 port map( A1 => n16482, A2 => n62163, B1 => n62161, B2 => 
                           n4953, C1 => n16636, C2 => n62159, ZN => n7888);
   U8042 : OAI221_X1 port map( B1 => n61954, B2 => n4671, C1 => n61951, C2 => 
                           n4695, A => n7863, ZN => n7843);
   U8043 : AOI222_X1 port map( A1 => n62181, A2 => n4647, B1 => n61938, B2 => 
                           n4455, C1 => n16811, C2 => n62177, ZN => n7863);
   U8044 : OAI221_X1 port map( B1 => n61888, B2 => n3231, C1 => n61885, C2 => 
                           n3255, A => n7791, ZN => n7784);
   U8045 : AOI222_X1 port map( A1 => n16483, A2 => n62163, B1 => n62161, B2 => 
                           n4952, C1 => n16637, C2 => n62159, ZN => n7791);
   U8046 : OAI221_X1 port map( B1 => n61954, B2 => n4670, C1 => n61951, C2 => 
                           n4694, A => n7775, ZN => n7768);
   U8047 : AOI222_X1 port map( A1 => n62181, A2 => n4646, B1 => n61938, B2 => 
                           n4454, C1 => n16812, C2 => n62177, ZN => n7775);
   U8048 : OAI221_X1 port map( B1 => n61888, B2 => n3230, C1 => n61885, C2 => 
                           n3254, A => n7716, ZN => n7709);
   U8049 : AOI222_X1 port map( A1 => n16484, A2 => n62163, B1 => n62161, B2 => 
                           n4951, C1 => n16638, C2 => n62159, ZN => n7716);
   U8050 : OAI221_X1 port map( B1 => n61954, B2 => n4669, C1 => n61951, C2 => 
                           n4693, A => n7700, ZN => n7693);
   U8051 : AOI222_X1 port map( A1 => n62181, A2 => n4645, B1 => n61938, B2 => 
                           n4453, C1 => n16813, C2 => n62177, ZN => n7700);
   U8052 : OAI221_X1 port map( B1 => n61888, B2 => n3229, C1 => n61885, C2 => 
                           n3253, A => n7641, ZN => n7634);
   U8053 : AOI222_X1 port map( A1 => n16485, A2 => n62163, B1 => n62161, B2 => 
                           n4950, C1 => n16639, C2 => n62159, ZN => n7641);
   U8054 : OAI221_X1 port map( B1 => n61954, B2 => n4668, C1 => n61951, C2 => 
                           n4692, A => n7625, ZN => n7618);
   U8055 : AOI222_X1 port map( A1 => n62181, A2 => n4644, B1 => n61938, B2 => 
                           n4452, C1 => n16790, C2 => n62177, ZN => n7625);
   U8056 : OAI221_X1 port map( B1 => n61888, B2 => n3228, C1 => n61885, C2 => 
                           n3252, A => n7566, ZN => n7559);
   U8057 : AOI222_X1 port map( A1 => n16486, A2 => n62163, B1 => n62161, B2 => 
                           n4949, C1 => n16640, C2 => n62159, ZN => n7566);
   U8058 : OAI221_X1 port map( B1 => n61954, B2 => n4667, C1 => n61951, C2 => 
                           n4691, A => n7550, ZN => n7543);
   U8059 : AOI222_X1 port map( A1 => n62181, A2 => n4643, B1 => n61938, B2 => 
                           n4451, C1 => n16791, C2 => n62177, ZN => n7550);
   U8060 : OAI221_X1 port map( B1 => n61888, B2 => n3227, C1 => n61885, C2 => 
                           n3251, A => n7491, ZN => n7484);
   U8061 : AOI222_X1 port map( A1 => n16487, A2 => n62163, B1 => n62161, B2 => 
                           n4948, C1 => n16641, C2 => n62159, ZN => n7491);
   U8062 : OAI221_X1 port map( B1 => n61954, B2 => n4666, C1 => n61951, C2 => 
                           n4690, A => n7475, ZN => n7468);
   U8063 : AOI222_X1 port map( A1 => n62181, A2 => n4642, B1 => n61938, B2 => 
                           n4450, C1 => n16792, C2 => n62177, ZN => n7475);
   U8064 : OAI221_X1 port map( B1 => n61888, B2 => n3226, C1 => n61885, C2 => 
                           n3250, A => n7416, ZN => n7409);
   U8065 : AOI222_X1 port map( A1 => n16488, A2 => n62163, B1 => n62161, B2 => 
                           n4947, C1 => n16642, C2 => n62159, ZN => n7416);
   U8066 : OAI221_X1 port map( B1 => n61954, B2 => n4665, C1 => n61951, C2 => 
                           n4689, A => n7400, ZN => n7393);
   U8067 : AOI222_X1 port map( A1 => n62181, A2 => n4641, B1 => n61938, B2 => 
                           n4449, C1 => n16793, C2 => n62177, ZN => n7400);
   U8068 : OAI221_X1 port map( B1 => n61888, B2 => n3225, C1 => n61885, C2 => 
                           n3249, A => n7341, ZN => n7334);
   U8069 : AOI222_X1 port map( A1 => n16489, A2 => n62163, B1 => n62161, B2 => 
                           n4946, C1 => n16643, C2 => n62159, ZN => n7341);
   U8070 : OAI221_X1 port map( B1 => n61954, B2 => n4664, C1 => n61951, C2 => 
                           n4688, A => n7325, ZN => n7318);
   U8071 : AOI222_X1 port map( A1 => n62181, A2 => n4640, B1 => n61937, B2 => 
                           n4448, C1 => n16799, C2 => n62177, ZN => n7325);
   U8072 : OAI221_X1 port map( B1 => n61888, B2 => n3223, C1 => n61885, C2 => 
                           n3247, A => n7191, ZN => n7184);
   U8073 : AOI222_X1 port map( A1 => n16491, A2 => n62163, B1 => n62161, B2 => 
                           n4944, C1 => n16645, C2 => n62159, ZN => n7191);
   U8074 : OAI221_X1 port map( B1 => n61954, B2 => n4662, C1 => n61951, C2 => 
                           n4686, A => n7175, ZN => n7168);
   U8075 : AOI222_X1 port map( A1 => n62181, A2 => n4638, B1 => n61937, B2 => 
                           n4446, C1 => n16800, C2 => n62177, ZN => n7175);
   U8076 : OAI221_X1 port map( B1 => n61889, B2 => n3220, C1 => n61886, C2 => 
                           n3244, A => n6966, ZN => n6959);
   U8077 : AOI222_X1 port map( A1 => n16494, A2 => n62162, B1 => n62160, B2 => 
                           n4941, C1 => n16648, C2 => n62158, ZN => n6966);
   U8078 : OAI221_X1 port map( B1 => n6059, B2 => n2790, C1 => n61704, C2 => 
                           n2862, A => n6974, ZN => n6967);
   U8079 : AOI222_X1 port map( A1 => n16730, A2 => n62172, B1 => n651, B2 => 
                           n61868, C1 => n16754, C2 => n62170, ZN => n6974);
   U8080 : OAI221_X1 port map( B1 => n61955, B2 => n4659, C1 => n61952, C2 => 
                           n4683, A => n6950, ZN => n6943);
   U8081 : AOI222_X1 port map( A1 => n62180, A2 => n4635, B1 => n61937, B2 => 
                           n4443, C1 => n16801, C2 => n62176, ZN => n6950);
   U8082 : OAI221_X1 port map( B1 => n6089, B2 => n3906, C1 => n61684, C2 => 
                           n1798, A => n6994, ZN => n6987);
   U8083 : AOI222_X1 port map( A1 => n15527, A2 => n62140, B1 => n15719, B2 => 
                           n61819, C1 => n3110, C2 => n62142, ZN => n6994);
   U8084 : OAI221_X1 port map( B1 => n4849, B2 => n61526, C1 => n3166, C2 => 
                           n61523, A => n14395, ZN => n14388);
   U8085 : AOI222_X1 port map( A1 => n61520, A2 => n53139, B1 => n61518, B2 => 
                           n4801, C1 => n61515, C2 => n53187, ZN => n14395);
   U8086 : OAI221_X1 port map( B1 => n1498, B2 => n61577, C1 => n1474, C2 => 
                           n61574, A => n14387, ZN => n14380);
   U8087 : AOI222_X1 port map( A1 => n61571, A2 => n5017, B1 => n61569, B2 => 
                           n5041, C1 => n61566, C2 => n52871, ZN => n14387);
   U8088 : OAI221_X1 port map( B1 => n4543, B2 => n61628, C1 => n4519, C2 => 
                           n61625, A => n14379, ZN => n14372);
   U8089 : AOI222_X1 port map( A1 => n61622, A2 => n4394, B1 => n61620, B2 => 
                           n4471, C1 => n61617, C2 => n4495, ZN => n14379);
   U8090 : OAI221_X1 port map( B1 => n3540, B2 => n61322, C1 => n3516, C2 => 
                           n61319, A => n14431, ZN => n14424);
   U8091 : AOI222_X1 port map( A1 => n61316, A2 => n53695, B1 => n61314, B2 => 
                           n53719, C1 => n61311, C2 => n53743, ZN => n14431);
   U8092 : OAI221_X1 port map( B1 => n3886, B2 => n61373, C1 => n3862, C2 => 
                           n61370, A => n14423, ZN => n14416);
   U8093 : AOI222_X1 port map( A1 => n61367, A2 => n53931, B1 => n61365, B2 => 
                           n53955, C1 => n61362, C2 => n53979, ZN => n14423);
   U8094 : OAI221_X1 port map( B1 => n2161, B2 => n61424, C1 => n2137, C2 => 
                           n61421, A => n14415, ZN => n14408);
   U8095 : AOI222_X1 port map( A1 => n61418, A2 => n54171, B1 => n61416, B2 => 
                           n54195, C1 => n61413, C2 => n54219, ZN => n14415);
   U8096 : OAI221_X1 port map( B1 => n4848, B2 => n61526, C1 => n3165, C2 => 
                           n61523, A => n9904, ZN => n9897);
   U8097 : AOI222_X1 port map( A1 => n61520, A2 => n53138, B1 => n61518, B2 => 
                           n4800, C1 => n61515, C2 => n53186, ZN => n9904);
   U8098 : OAI221_X1 port map( B1 => n1497, B2 => n61577, C1 => n1473, C2 => 
                           n61574, A => n9896, ZN => n9889);
   U8099 : AOI222_X1 port map( A1 => n61571, A2 => n5016, B1 => n61569, B2 => 
                           n5040, C1 => n61566, C2 => n52870, ZN => n9896);
   U8100 : OAI221_X1 port map( B1 => n4542, B2 => n61628, C1 => n4518, C2 => 
                           n61625, A => n9888, ZN => n9881);
   U8101 : AOI222_X1 port map( A1 => n61622, A2 => n4393, B1 => n61620, B2 => 
                           n4470, C1 => n61617, C2 => n4494, ZN => n9888);
   U8102 : OAI221_X1 port map( B1 => n3539, B2 => n61322, C1 => n3515, C2 => 
                           n61319, A => n14356, ZN => n14349);
   U8103 : AOI222_X1 port map( A1 => n61316, A2 => n53694, B1 => n61314, B2 => 
                           n53718, C1 => n61311, C2 => n53742, ZN => n14356);
   U8104 : OAI221_X1 port map( B1 => n3885, B2 => n61373, C1 => n3861, C2 => 
                           n61370, A => n14348, ZN => n14341);
   U8105 : AOI222_X1 port map( A1 => n61367, A2 => n53930, B1 => n61365, B2 => 
                           n53954, C1 => n61362, C2 => n53978, ZN => n14348);
   U8106 : OAI221_X1 port map( B1 => n2160, B2 => n61424, C1 => n2136, C2 => 
                           n61421, A => n9924, ZN => n9917);
   U8107 : AOI222_X1 port map( A1 => n61418, A2 => n54170, B1 => n61416, B2 => 
                           n54194, C1 => n61413, C2 => n54218, ZN => n9924);
   U8108 : OAI221_X1 port map( B1 => n4847, B2 => n61526, C1 => n3164, C2 => 
                           n61523, A => n9829, ZN => n9822);
   U8109 : AOI222_X1 port map( A1 => n61520, A2 => n53137, B1 => n61518, B2 => 
                           n4799, C1 => n61515, C2 => n4823, ZN => n9829);
   U8110 : OAI221_X1 port map( B1 => n1496, B2 => n61577, C1 => n1472, C2 => 
                           n61574, A => n9821, ZN => n9814);
   U8111 : AOI222_X1 port map( A1 => n61571, A2 => n5015, B1 => n61569, B2 => 
                           n5039, C1 => n61566, C2 => n52869, ZN => n9821);
   U8112 : OAI221_X1 port map( B1 => n4541, B2 => n61628, C1 => n4517, C2 => 
                           n61625, A => n9813, ZN => n9742);
   U8113 : AOI222_X1 port map( A1 => n61622, A2 => n4392, B1 => n61620, B2 => 
                           n4469, C1 => n61617, C2 => n4493, ZN => n9813);
   U8114 : OAI221_X1 port map( B1 => n3538, B2 => n61322, C1 => n3514, C2 => 
                           n61319, A => n9865, ZN => n9858);
   U8115 : AOI222_X1 port map( A1 => n61316, A2 => n53693, B1 => n61314, B2 => 
                           n53717, C1 => n61311, C2 => n53741, ZN => n9865);
   U8116 : OAI221_X1 port map( B1 => n3884, B2 => n61373, C1 => n3860, C2 => 
                           n61370, A => n9857, ZN => n9850);
   U8117 : AOI222_X1 port map( A1 => n61367, A2 => n53929, B1 => n61365, B2 => 
                           n53953, C1 => n61362, C2 => n53977, ZN => n9857);
   U8118 : OAI221_X1 port map( B1 => n2159, B2 => n61424, C1 => n2135, C2 => 
                           n61421, A => n9849, ZN => n9842);
   U8119 : AOI222_X1 port map( A1 => n61418, A2 => n54169, B1 => n61416, B2 => 
                           n54193, C1 => n61413, C2 => n54217, ZN => n9849);
   U8120 : OAI221_X1 port map( B1 => n4846, B2 => n61526, C1 => n3163, C2 => 
                           n61523, A => n9690, ZN => n9683);
   U8121 : AOI222_X1 port map( A1 => n61520, A2 => n53136, B1 => n61518, B2 => 
                           n4798, C1 => n61515, C2 => n4822, ZN => n9690);
   U8122 : OAI221_X1 port map( B1 => n1495, B2 => n61577, C1 => n1471, C2 => 
                           n61574, A => n9682, ZN => n9675);
   U8123 : AOI222_X1 port map( A1 => n61571, A2 => n5014, B1 => n61569, B2 => 
                           n5038, C1 => n61566, C2 => n52868, ZN => n9682);
   U8124 : OAI221_X1 port map( B1 => n4540, B2 => n61628, C1 => n4516, C2 => 
                           n61625, A => n9674, ZN => n9667);
   U8125 : AOI222_X1 port map( A1 => n61622, A2 => n4391, B1 => n61620, B2 => 
                           n4468, C1 => n61617, C2 => n4492, ZN => n9674);
   U8126 : OAI221_X1 port map( B1 => n3537, B2 => n61322, C1 => n3513, C2 => 
                           n61319, A => n9726, ZN => n9719);
   U8127 : AOI222_X1 port map( A1 => n61316, A2 => n53692, B1 => n61314, B2 => 
                           n53716, C1 => n61311, C2 => n53740, ZN => n9726);
   U8128 : OAI221_X1 port map( B1 => n3883, B2 => n61373, C1 => n3859, C2 => 
                           n61370, A => n9718, ZN => n9711);
   U8129 : AOI222_X1 port map( A1 => n61367, A2 => n53928, B1 => n61365, B2 => 
                           n53952, C1 => n61362, C2 => n53976, ZN => n9718);
   U8130 : OAI221_X1 port map( B1 => n2158, B2 => n61424, C1 => n2134, C2 => 
                           n61421, A => n9710, ZN => n9703);
   U8131 : AOI222_X1 port map( A1 => n61418, A2 => n54168, B1 => n61416, B2 => 
                           n54192, C1 => n61413, C2 => n54216, ZN => n9710);
   U8132 : OAI221_X1 port map( B1 => n4845, B2 => n61527, C1 => n3162, C2 => 
                           n61524, A => n9599, ZN => n9592);
   U8133 : AOI222_X1 port map( A1 => n61521, A2 => n53135, B1 => n61518, B2 => 
                           n4797, C1 => n61515, C2 => n4821, ZN => n9599);
   U8134 : OAI221_X1 port map( B1 => n1494, B2 => n61578, C1 => n1470, C2 => 
                           n61575, A => n9591, ZN => n9584);
   U8135 : AOI222_X1 port map( A1 => n61572, A2 => n5013, B1 => n61569, B2 => 
                           n5037, C1 => n61566, C2 => n52867, ZN => n9591);
   U8136 : OAI221_X1 port map( B1 => n4539, B2 => n61629, C1 => n4515, C2 => 
                           n61626, A => n9583, ZN => n9576);
   U8137 : AOI222_X1 port map( A1 => n61623, A2 => n4390, B1 => n61620, B2 => 
                           n4467, C1 => n61617, C2 => n4491, ZN => n9583);
   U8138 : OAI221_X1 port map( B1 => n3536, B2 => n61323, C1 => n3512, C2 => 
                           n61320, A => n9651, ZN => n9644);
   U8139 : AOI222_X1 port map( A1 => n61317, A2 => n53691, B1 => n61314, B2 => 
                           n53715, C1 => n61311, C2 => n53739, ZN => n9651);
   U8140 : OAI221_X1 port map( B1 => n3882, B2 => n61374, C1 => n3858, C2 => 
                           n61371, A => n9643, ZN => n9636);
   U8141 : AOI222_X1 port map( A1 => n61368, A2 => n53927, B1 => n61365, B2 => 
                           n53951, C1 => n61362, C2 => n53975, ZN => n9643);
   U8142 : OAI221_X1 port map( B1 => n2157, B2 => n61425, C1 => n2133, C2 => 
                           n61422, A => n9635, ZN => n9628);
   U8143 : AOI222_X1 port map( A1 => n61419, A2 => n54167, B1 => n61416, B2 => 
                           n54191, C1 => n61413, C2 => n54215, ZN => n9635);
   U8144 : OAI221_X1 port map( B1 => n4844, B2 => n61527, C1 => n3161, C2 => 
                           n61524, A => n9524, ZN => n9517);
   U8145 : AOI222_X1 port map( A1 => n61521, A2 => n53134, B1 => n61518, B2 => 
                           n4796, C1 => n61515, C2 => n4820, ZN => n9524);
   U8146 : OAI221_X1 port map( B1 => n1493, B2 => n61578, C1 => n1469, C2 => 
                           n61575, A => n9516, ZN => n9509);
   U8147 : AOI222_X1 port map( A1 => n61572, A2 => n5012, B1 => n61569, B2 => 
                           n5036, C1 => n61566, C2 => n52866, ZN => n9516);
   U8148 : OAI221_X1 port map( B1 => n4538, B2 => n61629, C1 => n4514, C2 => 
                           n61626, A => n9508, ZN => n9501);
   U8149 : AOI222_X1 port map( A1 => n61623, A2 => n4389, B1 => n61620, B2 => 
                           n4466, C1 => n61617, C2 => n4490, ZN => n9508);
   U8150 : OAI221_X1 port map( B1 => n3535, B2 => n61323, C1 => n3511, C2 => 
                           n61320, A => n9560, ZN => n9553);
   U8151 : AOI222_X1 port map( A1 => n61317, A2 => n53690, B1 => n61314, B2 => 
                           n53714, C1 => n61311, C2 => n53738, ZN => n9560);
   U8152 : OAI221_X1 port map( B1 => n3881, B2 => n61374, C1 => n3857, C2 => 
                           n61371, A => n9552, ZN => n9545);
   U8153 : AOI222_X1 port map( A1 => n61368, A2 => n53926, B1 => n61365, B2 => 
                           n53950, C1 => n61362, C2 => n53974, ZN => n9552);
   U8154 : OAI221_X1 port map( B1 => n2156, B2 => n61425, C1 => n2132, C2 => 
                           n61422, A => n9544, ZN => n9537);
   U8155 : AOI222_X1 port map( A1 => n61419, A2 => n54166, B1 => n61416, B2 => 
                           n54190, C1 => n61413, C2 => n54214, ZN => n9544);
   U8156 : OAI221_X1 port map( B1 => n4843, B2 => n61527, C1 => n4833, C2 => 
                           n61524, A => n9449, ZN => n9442);
   U8157 : AOI222_X1 port map( A1 => n61521, A2 => n53133, B1 => n61518, B2 => 
                           n4795, C1 => n61515, C2 => n4819, ZN => n9449);
   U8158 : OAI221_X1 port map( B1 => n1492, B2 => n61578, C1 => n1468, C2 => 
                           n61575, A => n9441, ZN => n9434);
   U8159 : AOI222_X1 port map( A1 => n61572, A2 => n5011, B1 => n61569, B2 => 
                           n5035, C1 => n61566, C2 => n52865, ZN => n9441);
   U8160 : OAI221_X1 port map( B1 => n4537, B2 => n61629, C1 => n4513, C2 => 
                           n61626, A => n9433, ZN => n9426);
   U8161 : AOI222_X1 port map( A1 => n61623, A2 => n4388, B1 => n61620, B2 => 
                           n4465, C1 => n61617, C2 => n4489, ZN => n9433);
   U8162 : OAI221_X1 port map( B1 => n3534, B2 => n61323, C1 => n3510, C2 => 
                           n61320, A => n9485, ZN => n9478);
   U8163 : AOI222_X1 port map( A1 => n61317, A2 => n53689, B1 => n61314, B2 => 
                           n53713, C1 => n61311, C2 => n53737, ZN => n9485);
   U8164 : OAI221_X1 port map( B1 => n3880, B2 => n61374, C1 => n3856, C2 => 
                           n61371, A => n9477, ZN => n9470);
   U8165 : AOI222_X1 port map( A1 => n61368, A2 => n53925, B1 => n61365, B2 => 
                           n53949, C1 => n61362, C2 => n53973, ZN => n9477);
   U8166 : OAI221_X1 port map( B1 => n2155, B2 => n61425, C1 => n2131, C2 => 
                           n61422, A => n9469, ZN => n9462);
   U8167 : AOI222_X1 port map( A1 => n61419, A2 => n54165, B1 => n61416, B2 => 
                           n54189, C1 => n61413, C2 => n54213, ZN => n9469);
   U8168 : OAI221_X1 port map( B1 => n4842, B2 => n61527, C1 => n4832, C2 => 
                           n61524, A => n9374, ZN => n9367);
   U8169 : AOI222_X1 port map( A1 => n61521, A2 => n53132, B1 => n61518, B2 => 
                           n4794, C1 => n61515, C2 => n4818, ZN => n9374);
   U8170 : OAI221_X1 port map( B1 => n1491, B2 => n61578, C1 => n1467, C2 => 
                           n61575, A => n9366, ZN => n9359);
   U8171 : AOI222_X1 port map( A1 => n61572, A2 => n5010, B1 => n61569, B2 => 
                           n5034, C1 => n61566, C2 => n52864, ZN => n9366);
   U8172 : OAI221_X1 port map( B1 => n4536, B2 => n61629, C1 => n4512, C2 => 
                           n61626, A => n9358, ZN => n9351);
   U8173 : AOI222_X1 port map( A1 => n61623, A2 => n4387, B1 => n61620, B2 => 
                           n4464, C1 => n61617, C2 => n4488, ZN => n9358);
   U8174 : OAI221_X1 port map( B1 => n3533, B2 => n61323, C1 => n3509, C2 => 
                           n61320, A => n9410, ZN => n9403);
   U8175 : AOI222_X1 port map( A1 => n61317, A2 => n53688, B1 => n61314, B2 => 
                           n53712, C1 => n61311, C2 => n53736, ZN => n9410);
   U8176 : OAI221_X1 port map( B1 => n3879, B2 => n61374, C1 => n3855, C2 => 
                           n61371, A => n9402, ZN => n9395);
   U8177 : AOI222_X1 port map( A1 => n61368, A2 => n53924, B1 => n61365, B2 => 
                           n53948, C1 => n61362, C2 => n53972, ZN => n9402);
   U8178 : OAI221_X1 port map( B1 => n2154, B2 => n61425, C1 => n2130, C2 => 
                           n61422, A => n9394, ZN => n9387);
   U8179 : AOI222_X1 port map( A1 => n61419, A2 => n54164, B1 => n61416, B2 => 
                           n54188, C1 => n61413, C2 => n54212, ZN => n9394);
   U8180 : OAI221_X1 port map( B1 => n4841, B2 => n61527, C1 => n4831, C2 => 
                           n61524, A => n9235, ZN => n9228);
   U8181 : AOI222_X1 port map( A1 => n61521, A2 => n53131, B1 => n61518, B2 => 
                           n4793, C1 => n61515, C2 => n4817, ZN => n9235);
   U8182 : OAI221_X1 port map( B1 => n1490, B2 => n61578, C1 => n1466, C2 => 
                           n61575, A => n9227, ZN => n9220);
   U8183 : AOI222_X1 port map( A1 => n61572, A2 => n5009, B1 => n61569, B2 => 
                           n5033, C1 => n61566, C2 => n52863, ZN => n9227);
   U8184 : OAI221_X1 port map( B1 => n4535, B2 => n61629, C1 => n4511, C2 => 
                           n61626, A => n9219, ZN => n9212);
   U8185 : AOI222_X1 port map( A1 => n61623, A2 => n4386, B1 => n61620, B2 => 
                           n4463, C1 => n61617, C2 => n4487, ZN => n9219);
   U8186 : OAI221_X1 port map( B1 => n3532, B2 => n61323, C1 => n3508, C2 => 
                           n61320, A => n9271, ZN => n9264);
   U8187 : AOI222_X1 port map( A1 => n61317, A2 => n53687, B1 => n61314, B2 => 
                           n53711, C1 => n61311, C2 => n53735, ZN => n9271);
   U8188 : OAI221_X1 port map( B1 => n3878, B2 => n61374, C1 => n3854, C2 => 
                           n61371, A => n9263, ZN => n9256);
   U8189 : AOI222_X1 port map( A1 => n61368, A2 => n53923, B1 => n61365, B2 => 
                           n53947, C1 => n61362, C2 => n53971, ZN => n9263);
   U8190 : OAI221_X1 port map( B1 => n2153, B2 => n61425, C1 => n2129, C2 => 
                           n61422, A => n9255, ZN => n9248);
   U8191 : AOI222_X1 port map( A1 => n61419, A2 => n54163, B1 => n61416, B2 => 
                           n54187, C1 => n61413, C2 => n54211, ZN => n9255);
   U8192 : OAI221_X1 port map( B1 => n4840, B2 => n61527, C1 => n4830, C2 => 
                           n61524, A => n9160, ZN => n9153);
   U8193 : AOI222_X1 port map( A1 => n61521, A2 => n53130, B1 => n61518, B2 => 
                           n4792, C1 => n61515, C2 => n4816, ZN => n9160);
   U8194 : OAI221_X1 port map( B1 => n1489, B2 => n61578, C1 => n1465, C2 => 
                           n61575, A => n9152, ZN => n9145);
   U8195 : AOI222_X1 port map( A1 => n61572, A2 => n5008, B1 => n61569, B2 => 
                           n5032, C1 => n61566, C2 => n52862, ZN => n9152);
   U8196 : OAI221_X1 port map( B1 => n4534, B2 => n61629, C1 => n4510, C2 => 
                           n61626, A => n9144, ZN => n9137);
   U8197 : AOI222_X1 port map( A1 => n61623, A2 => n4385, B1 => n61620, B2 => 
                           n4462, C1 => n61617, C2 => n4486, ZN => n9144);
   U8198 : OAI221_X1 port map( B1 => n3531, B2 => n61323, C1 => n3507, C2 => 
                           n61320, A => n9196, ZN => n9189);
   U8199 : AOI222_X1 port map( A1 => n61317, A2 => n53686, B1 => n61314, B2 => 
                           n53710, C1 => n61311, C2 => n53734, ZN => n9196);
   U8200 : OAI221_X1 port map( B1 => n3877, B2 => n61374, C1 => n3853, C2 => 
                           n61371, A => n9188, ZN => n9181);
   U8201 : AOI222_X1 port map( A1 => n61368, A2 => n53922, B1 => n61365, B2 => 
                           n53946, C1 => n61362, C2 => n53970, ZN => n9188);
   U8202 : OAI221_X1 port map( B1 => n2152, B2 => n61425, C1 => n2128, C2 => 
                           n61422, A => n9180, ZN => n9173);
   U8203 : AOI222_X1 port map( A1 => n61419, A2 => n54162, B1 => n61416, B2 => 
                           n54186, C1 => n61413, C2 => n54210, ZN => n9180);
   U8204 : OAI221_X1 port map( B1 => n4839, B2 => n61527, C1 => n4829, C2 => 
                           n61524, A => n9085, ZN => n9078);
   U8205 : AOI222_X1 port map( A1 => n61521, A2 => n53129, B1 => n61518, B2 => 
                           n4791, C1 => n61515, C2 => n4815, ZN => n9085);
   U8206 : OAI221_X1 port map( B1 => n1488, B2 => n61578, C1 => n1464, C2 => 
                           n61575, A => n9077, ZN => n9070);
   U8207 : AOI222_X1 port map( A1 => n61572, A2 => n5007, B1 => n61569, B2 => 
                           n5031, C1 => n61566, C2 => n52861, ZN => n9077);
   U8208 : OAI221_X1 port map( B1 => n4533, B2 => n61629, C1 => n4509, C2 => 
                           n61626, A => n9069, ZN => n9062);
   U8209 : AOI222_X1 port map( A1 => n61623, A2 => n4384, B1 => n61620, B2 => 
                           n4461, C1 => n61617, C2 => n4485, ZN => n9069);
   U8210 : OAI221_X1 port map( B1 => n3530, B2 => n61323, C1 => n3506, C2 => 
                           n61320, A => n9121, ZN => n9114);
   U8211 : AOI222_X1 port map( A1 => n61317, A2 => n53685, B1 => n61314, B2 => 
                           n53709, C1 => n61311, C2 => n53733, ZN => n9121);
   U8212 : OAI221_X1 port map( B1 => n3876, B2 => n61374, C1 => n3852, C2 => 
                           n61371, A => n9113, ZN => n9106);
   U8213 : AOI222_X1 port map( A1 => n61368, A2 => n53921, B1 => n61365, B2 => 
                           n53945, C1 => n61362, C2 => n53969, ZN => n9113);
   U8214 : OAI221_X1 port map( B1 => n2151, B2 => n61425, C1 => n2127, C2 => 
                           n61422, A => n9105, ZN => n9098);
   U8215 : AOI222_X1 port map( A1 => n61419, A2 => n54161, B1 => n61416, B2 => 
                           n54185, C1 => n61413, C2 => n54209, ZN => n9105);
   U8216 : OAI221_X1 port map( B1 => n4838, B2 => n61527, C1 => n4828, C2 => 
                           n61524, A => n9010, ZN => n9003);
   U8217 : AOI222_X1 port map( A1 => n61521, A2 => n53128, B1 => n61518, B2 => 
                           n4790, C1 => n61515, C2 => n4814, ZN => n9010);
   U8218 : OAI221_X1 port map( B1 => n1487, B2 => n61578, C1 => n1463, C2 => 
                           n61575, A => n9002, ZN => n8995);
   U8219 : AOI222_X1 port map( A1 => n61572, A2 => n5006, B1 => n61569, B2 => 
                           n5030, C1 => n61566, C2 => n52860, ZN => n9002);
   U8220 : OAI221_X1 port map( B1 => n4532, B2 => n61629, C1 => n4508, C2 => 
                           n61626, A => n8994, ZN => n8987);
   U8221 : AOI222_X1 port map( A1 => n61623, A2 => n4383, B1 => n61620, B2 => 
                           n4460, C1 => n61617, C2 => n4484, ZN => n8994);
   U8222 : OAI221_X1 port map( B1 => n3529, B2 => n61323, C1 => n3505, C2 => 
                           n61320, A => n9046, ZN => n9039);
   U8223 : AOI222_X1 port map( A1 => n61317, A2 => n53684, B1 => n61314, B2 => 
                           n53708, C1 => n61311, C2 => n53732, ZN => n9046);
   U8224 : OAI221_X1 port map( B1 => n3875, B2 => n61374, C1 => n3851, C2 => 
                           n61371, A => n9038, ZN => n9031);
   U8225 : AOI222_X1 port map( A1 => n61368, A2 => n53920, B1 => n61365, B2 => 
                           n53944, C1 => n61362, C2 => n53968, ZN => n9038);
   U8226 : OAI221_X1 port map( B1 => n2150, B2 => n61425, C1 => n2126, C2 => 
                           n61422, A => n9030, ZN => n9023);
   U8227 : AOI222_X1 port map( A1 => n61419, A2 => n54160, B1 => n61416, B2 => 
                           n54184, C1 => n61413, C2 => n54208, ZN => n9030);
   U8228 : OAI221_X1 port map( B1 => n4837, B2 => n61527, C1 => n4827, C2 => 
                           n61524, A => n8935, ZN => n8928);
   U8229 : AOI222_X1 port map( A1 => n61521, A2 => n53127, B1 => n61517, B2 => 
                           n4789, C1 => n61514, C2 => n4813, ZN => n8935);
   U8230 : OAI221_X1 port map( B1 => n1486, B2 => n61578, C1 => n1462, C2 => 
                           n61575, A => n8927, ZN => n8920);
   U8231 : AOI222_X1 port map( A1 => n61572, A2 => n5005, B1 => n61568, B2 => 
                           n5029, C1 => n61565, C2 => n52859, ZN => n8927);
   U8232 : OAI221_X1 port map( B1 => n4531, B2 => n61629, C1 => n4507, C2 => 
                           n61626, A => n8919, ZN => n8912);
   U8233 : AOI222_X1 port map( A1 => n61623, A2 => n4382, B1 => n61619, B2 => 
                           n4459, C1 => n61616, C2 => n4483, ZN => n8919);
   U8234 : OAI221_X1 port map( B1 => n3528, B2 => n61323, C1 => n3504, C2 => 
                           n61320, A => n8971, ZN => n8964);
   U8235 : AOI222_X1 port map( A1 => n61317, A2 => n53683, B1 => n61313, B2 => 
                           n53707, C1 => n61310, C2 => n53731, ZN => n8971);
   U8236 : OAI221_X1 port map( B1 => n3874, B2 => n61374, C1 => n3850, C2 => 
                           n61371, A => n8963, ZN => n8956);
   U8237 : AOI222_X1 port map( A1 => n61368, A2 => n53919, B1 => n61364, B2 => 
                           n53943, C1 => n61361, C2 => n53967, ZN => n8963);
   U8238 : OAI221_X1 port map( B1 => n2149, B2 => n61425, C1 => n2125, C2 => 
                           n61422, A => n8955, ZN => n8948);
   U8239 : AOI222_X1 port map( A1 => n61419, A2 => n54159, B1 => n61415, B2 => 
                           n54183, C1 => n61412, C2 => n54207, ZN => n8955);
   U8240 : OAI221_X1 port map( B1 => n4836, B2 => n61527, C1 => n4826, C2 => 
                           n61524, A => n8860, ZN => n8853);
   U8241 : AOI222_X1 port map( A1 => n61521, A2 => n53126, B1 => n61517, B2 => 
                           n4788, C1 => n61514, C2 => n4812, ZN => n8860);
   U8242 : OAI221_X1 port map( B1 => n1485, B2 => n61578, C1 => n1461, C2 => 
                           n61575, A => n8852, ZN => n8845);
   U8243 : AOI222_X1 port map( A1 => n61572, A2 => n5004, B1 => n61568, B2 => 
                           n5028, C1 => n61565, C2 => n52858, ZN => n8852);
   U8244 : OAI221_X1 port map( B1 => n4530, B2 => n61629, C1 => n4506, C2 => 
                           n61626, A => n8844, ZN => n8837);
   U8245 : AOI222_X1 port map( A1 => n61623, A2 => n4381, B1 => n61619, B2 => 
                           n4458, C1 => n61616, C2 => n4482, ZN => n8844);
   U8246 : OAI221_X1 port map( B1 => n3527, B2 => n61323, C1 => n3503, C2 => 
                           n61320, A => n8896, ZN => n8889);
   U8247 : AOI222_X1 port map( A1 => n61317, A2 => n53682, B1 => n61313, B2 => 
                           n53706, C1 => n61310, C2 => n53730, ZN => n8896);
   U8248 : OAI221_X1 port map( B1 => n3873, B2 => n61374, C1 => n3849, C2 => 
                           n61371, A => n8888, ZN => n8881);
   U8249 : AOI222_X1 port map( A1 => n61368, A2 => n53918, B1 => n61364, B2 => 
                           n53942, C1 => n61361, C2 => n53966, ZN => n8888);
   U8250 : OAI221_X1 port map( B1 => n2148, B2 => n61425, C1 => n2124, C2 => 
                           n61422, A => n8880, ZN => n8873);
   U8251 : AOI222_X1 port map( A1 => n61419, A2 => n54158, B1 => n61415, B2 => 
                           n54182, C1 => n61412, C2 => n54206, ZN => n8880);
   U8252 : OAI221_X1 port map( B1 => n4835, B2 => n61527, C1 => n4825, C2 => 
                           n61524, A => n8785, ZN => n8778);
   U8253 : AOI222_X1 port map( A1 => n61521, A2 => n53125, B1 => n61517, B2 => 
                           n4787, C1 => n61514, C2 => n4811, ZN => n8785);
   U8254 : OAI221_X1 port map( B1 => n1484, B2 => n61578, C1 => n1460, C2 => 
                           n61575, A => n8777, ZN => n8770);
   U8255 : AOI222_X1 port map( A1 => n61572, A2 => n5003, B1 => n61568, B2 => 
                           n5027, C1 => n61565, C2 => n52857, ZN => n8777);
   U8256 : OAI221_X1 port map( B1 => n4529, B2 => n61629, C1 => n4505, C2 => 
                           n61626, A => n8769, ZN => n8762);
   U8257 : AOI222_X1 port map( A1 => n61623, A2 => n4380, B1 => n61619, B2 => 
                           n4457, C1 => n61616, C2 => n4481, ZN => n8769);
   U8258 : OAI221_X1 port map( B1 => n3526, B2 => n61323, C1 => n3502, C2 => 
                           n61320, A => n8821, ZN => n8814);
   U8259 : AOI222_X1 port map( A1 => n61317, A2 => n53681, B1 => n61313, B2 => 
                           n53705, C1 => n61310, C2 => n53729, ZN => n8821);
   U8260 : OAI221_X1 port map( B1 => n3872, B2 => n61374, C1 => n3848, C2 => 
                           n61371, A => n8813, ZN => n8806);
   U8261 : AOI222_X1 port map( A1 => n61368, A2 => n53917, B1 => n61364, B2 => 
                           n53941, C1 => n61361, C2 => n53965, ZN => n8813);
   U8262 : OAI221_X1 port map( B1 => n2147, B2 => n61425, C1 => n2123, C2 => 
                           n61422, A => n8805, ZN => n8798);
   U8263 : AOI222_X1 port map( A1 => n61419, A2 => n54157, B1 => n61415, B2 => 
                           n54181, C1 => n61412, C2 => n54205, ZN => n8805);
   U8264 : OAI221_X1 port map( B1 => n4834, B2 => n61527, C1 => n4824, C2 => 
                           n61524, A => n8710, ZN => n8703);
   U8265 : AOI222_X1 port map( A1 => n61521, A2 => n53124, B1 => n61517, B2 => 
                           n4786, C1 => n61514, C2 => n4810, ZN => n8710);
   U8266 : OAI221_X1 port map( B1 => n1483, B2 => n61578, C1 => n1459, C2 => 
                           n61575, A => n8702, ZN => n8695);
   U8267 : AOI222_X1 port map( A1 => n61572, A2 => n5002, B1 => n61568, B2 => 
                           n5026, C1 => n61565, C2 => n52856, ZN => n8702);
   U8268 : OAI221_X1 port map( B1 => n4528, B2 => n61629, C1 => n4504, C2 => 
                           n61626, A => n8694, ZN => n8687);
   U8269 : AOI222_X1 port map( A1 => n61623, A2 => n4379, B1 => n61619, B2 => 
                           n4456, C1 => n61616, C2 => n4480, ZN => n8694);
   U8270 : OAI221_X1 port map( B1 => n3525, B2 => n61323, C1 => n3501, C2 => 
                           n61320, A => n8746, ZN => n8739);
   U8271 : AOI222_X1 port map( A1 => n61317, A2 => n53680, B1 => n61313, B2 => 
                           n53704, C1 => n61310, C2 => n53728, ZN => n8746);
   U8272 : OAI221_X1 port map( B1 => n3871, B2 => n61374, C1 => n3847, C2 => 
                           n61371, A => n8738, ZN => n8731);
   U8273 : AOI222_X1 port map( A1 => n61368, A2 => n53916, B1 => n61364, B2 => 
                           n53940, C1 => n61361, C2 => n53964, ZN => n8738);
   U8274 : OAI221_X1 port map( B1 => n2146, B2 => n61425, C1 => n2122, C2 => 
                           n61422, A => n8730, ZN => n8723);
   U8275 : AOI222_X1 port map( A1 => n61419, A2 => n54156, B1 => n61415, B2 => 
                           n54180, C1 => n61412, C2 => n54204, ZN => n8730);
   U8276 : OAI221_X1 port map( B1 => n4857, B2 => n61526, C1 => n3174, C2 => 
                           n61523, A => n15015, ZN => n15006);
   U8277 : AOI222_X1 port map( A1 => n61520, A2 => n53147, B1 => n61519, B2 => 
                           n4809, C1 => n61516, C2 => n53195, ZN => n15015);
   U8278 : OAI221_X1 port map( B1 => n1506, B2 => n61577, C1 => n1482, C2 => 
                           n61574, A => n15003, ZN => n14994);
   U8279 : AOI222_X1 port map( A1 => n61571, A2 => n5025, B1 => n61570, B2 => 
                           n5049, C1 => n61567, C2 => n52879, ZN => n15003);
   U8280 : OAI221_X1 port map( B1 => n4551, B2 => n61628, C1 => n4527, C2 => 
                           n61625, A => n14991, ZN => n14972);
   U8281 : AOI222_X1 port map( A1 => n61622, A2 => n4402, B1 => n61621, B2 => 
                           n4479, C1 => n61618, C2 => n4503, ZN => n14991);
   U8282 : OAI221_X1 port map( B1 => n3548, B2 => n61322, C1 => n3524, C2 => 
                           n61319, A => n15062, ZN => n15052);
   U8283 : AOI222_X1 port map( A1 => n61316, A2 => n53703, B1 => n61315, B2 => 
                           n53727, C1 => n61312, C2 => n53751, ZN => n15062);
   U8284 : OAI221_X1 port map( B1 => n3894, B2 => n61373, C1 => n3870, C2 => 
                           n61370, A => n15051, ZN => n15042);
   U8285 : AOI222_X1 port map( A1 => n61367, A2 => n53939, B1 => n61366, B2 => 
                           n53963, C1 => n61363, C2 => n53987, ZN => n15051);
   U8286 : OAI221_X1 port map( B1 => n2169, B2 => n61424, C1 => n2145, C2 => 
                           n61421, A => n15040, ZN => n15031);
   U8287 : AOI222_X1 port map( A1 => n61418, A2 => n54179, B1 => n61417, B2 => 
                           n54203, C1 => n61414, C2 => n54227, ZN => n15040);
   U8288 : OAI221_X1 port map( B1 => n4856, B2 => n61526, C1 => n3173, C2 => 
                           n61523, A => n14920, ZN => n14913);
   U8289 : AOI222_X1 port map( A1 => n61520, A2 => n53146, B1 => n61519, B2 => 
                           n4808, C1 => n61516, C2 => n53194, ZN => n14920);
   U8290 : OAI221_X1 port map( B1 => n1505, B2 => n61577, C1 => n1481, C2 => 
                           n61574, A => n14912, ZN => n14905);
   U8291 : AOI222_X1 port map( A1 => n61571, A2 => n5024, B1 => n61570, B2 => 
                           n5048, C1 => n61567, C2 => n52878, ZN => n14912);
   U8292 : OAI221_X1 port map( B1 => n4550, B2 => n61628, C1 => n4526, C2 => 
                           n61625, A => n14904, ZN => n14897);
   U8293 : AOI222_X1 port map( A1 => n61622, A2 => n4401, B1 => n61621, B2 => 
                           n4478, C1 => n61618, C2 => n4502, ZN => n14904);
   U8294 : OAI221_X1 port map( B1 => n3547, B2 => n61322, C1 => n3523, C2 => 
                           n61319, A => n14956, ZN => n14949);
   U8295 : AOI222_X1 port map( A1 => n61316, A2 => n53702, B1 => n61315, B2 => 
                           n53726, C1 => n61312, C2 => n53750, ZN => n14956);
   U8296 : OAI221_X1 port map( B1 => n3893, B2 => n61373, C1 => n3869, C2 => 
                           n61370, A => n14948, ZN => n14941);
   U8297 : AOI222_X1 port map( A1 => n61367, A2 => n53938, B1 => n61366, B2 => 
                           n53962, C1 => n61363, C2 => n53986, ZN => n14948);
   U8298 : OAI221_X1 port map( B1 => n2168, B2 => n61424, C1 => n2144, C2 => 
                           n61421, A => n14940, ZN => n14933);
   U8299 : AOI222_X1 port map( A1 => n61418, A2 => n54178, B1 => n61417, B2 => 
                           n54202, C1 => n61414, C2 => n54226, ZN => n14940);
   U8300 : OAI221_X1 port map( B1 => n4855, B2 => n61526, C1 => n3172, C2 => 
                           n61523, A => n14845, ZN => n14838);
   U8301 : AOI222_X1 port map( A1 => n61520, A2 => n53145, B1 => n61519, B2 => 
                           n4807, C1 => n61516, C2 => n53193, ZN => n14845);
   U8302 : OAI221_X1 port map( B1 => n1504, B2 => n61577, C1 => n1480, C2 => 
                           n61574, A => n14837, ZN => n14830);
   U8303 : AOI222_X1 port map( A1 => n61571, A2 => n5023, B1 => n61570, B2 => 
                           n5047, C1 => n61567, C2 => n52877, ZN => n14837);
   U8304 : OAI221_X1 port map( B1 => n4549, B2 => n61628, C1 => n4525, C2 => 
                           n61625, A => n14829, ZN => n14822);
   U8305 : AOI222_X1 port map( A1 => n61622, A2 => n4400, B1 => n61621, B2 => 
                           n4477, C1 => n61618, C2 => n4501, ZN => n14829);
   U8306 : OAI221_X1 port map( B1 => n3546, B2 => n61322, C1 => n3522, C2 => 
                           n61319, A => n14881, ZN => n14874);
   U8307 : AOI222_X1 port map( A1 => n61316, A2 => n53701, B1 => n61315, B2 => 
                           n53725, C1 => n61312, C2 => n53749, ZN => n14881);
   U8308 : OAI221_X1 port map( B1 => n3892, B2 => n61373, C1 => n3868, C2 => 
                           n61370, A => n14873, ZN => n14866);
   U8309 : AOI222_X1 port map( A1 => n61367, A2 => n53937, B1 => n61366, B2 => 
                           n53961, C1 => n61363, C2 => n53985, ZN => n14873);
   U8310 : OAI221_X1 port map( B1 => n2167, B2 => n61424, C1 => n2143, C2 => 
                           n61421, A => n14865, ZN => n14858);
   U8311 : AOI222_X1 port map( A1 => n61418, A2 => n54177, B1 => n61417, B2 => 
                           n54201, C1 => n61414, C2 => n54225, ZN => n14865);
   U8312 : OAI221_X1 port map( B1 => n4854, B2 => n61526, C1 => n3171, C2 => 
                           n61523, A => n14770, ZN => n14763);
   U8313 : AOI222_X1 port map( A1 => n61520, A2 => n53144, B1 => n61519, B2 => 
                           n4806, C1 => n61516, C2 => n53192, ZN => n14770);
   U8314 : OAI221_X1 port map( B1 => n1503, B2 => n61577, C1 => n1479, C2 => 
                           n61574, A => n14762, ZN => n14755);
   U8315 : AOI222_X1 port map( A1 => n61571, A2 => n5022, B1 => n61570, B2 => 
                           n5046, C1 => n61567, C2 => n52876, ZN => n14762);
   U8316 : OAI221_X1 port map( B1 => n4548, B2 => n61628, C1 => n4524, C2 => 
                           n61625, A => n14754, ZN => n14747);
   U8317 : AOI222_X1 port map( A1 => n61622, A2 => n4399, B1 => n61621, B2 => 
                           n4476, C1 => n61618, C2 => n4500, ZN => n14754);
   U8318 : OAI221_X1 port map( B1 => n3545, B2 => n61322, C1 => n3521, C2 => 
                           n61319, A => n14806, ZN => n14799);
   U8319 : AOI222_X1 port map( A1 => n61316, A2 => n53700, B1 => n61315, B2 => 
                           n53724, C1 => n61312, C2 => n53748, ZN => n14806);
   U8320 : OAI221_X1 port map( B1 => n3891, B2 => n61373, C1 => n3867, C2 => 
                           n61370, A => n14798, ZN => n14791);
   U8321 : AOI222_X1 port map( A1 => n61367, A2 => n53936, B1 => n61366, B2 => 
                           n53960, C1 => n61363, C2 => n53984, ZN => n14798);
   U8322 : OAI221_X1 port map( B1 => n2166, B2 => n61424, C1 => n2142, C2 => 
                           n61421, A => n14790, ZN => n14783);
   U8323 : AOI222_X1 port map( A1 => n61418, A2 => n54176, B1 => n61417, B2 => 
                           n54200, C1 => n61414, C2 => n54224, ZN => n14790);
   U8324 : OAI221_X1 port map( B1 => n4853, B2 => n61526, C1 => n3170, C2 => 
                           n61523, A => n14695, ZN => n14688);
   U8325 : AOI222_X1 port map( A1 => n61520, A2 => n53143, B1 => n61519, B2 => 
                           n4805, C1 => n61516, C2 => n53191, ZN => n14695);
   U8326 : OAI221_X1 port map( B1 => n1502, B2 => n61577, C1 => n1478, C2 => 
                           n61574, A => n14687, ZN => n14680);
   U8327 : AOI222_X1 port map( A1 => n61571, A2 => n5021, B1 => n61570, B2 => 
                           n5045, C1 => n61567, C2 => n52875, ZN => n14687);
   U8328 : OAI221_X1 port map( B1 => n4547, B2 => n61628, C1 => n4523, C2 => 
                           n61625, A => n14679, ZN => n14672);
   U8329 : AOI222_X1 port map( A1 => n61622, A2 => n4398, B1 => n61621, B2 => 
                           n4475, C1 => n61618, C2 => n4499, ZN => n14679);
   U8330 : OAI221_X1 port map( B1 => n3544, B2 => n61322, C1 => n3520, C2 => 
                           n61319, A => n14731, ZN => n14724);
   U8331 : AOI222_X1 port map( A1 => n61316, A2 => n53699, B1 => n61315, B2 => 
                           n53723, C1 => n61312, C2 => n53747, ZN => n14731);
   U8332 : OAI221_X1 port map( B1 => n3890, B2 => n61373, C1 => n3866, C2 => 
                           n61370, A => n14723, ZN => n14716);
   U8333 : AOI222_X1 port map( A1 => n61367, A2 => n53935, B1 => n61366, B2 => 
                           n53959, C1 => n61363, C2 => n53983, ZN => n14723);
   U8334 : OAI221_X1 port map( B1 => n2165, B2 => n61424, C1 => n2141, C2 => 
                           n61421, A => n14715, ZN => n14708);
   U8335 : AOI222_X1 port map( A1 => n61418, A2 => n54175, B1 => n61417, B2 => 
                           n54199, C1 => n61414, C2 => n54223, ZN => n14715);
   U8336 : OAI221_X1 port map( B1 => n4852, B2 => n61526, C1 => n3169, C2 => 
                           n61523, A => n14620, ZN => n14613);
   U8337 : AOI222_X1 port map( A1 => n61520, A2 => n53142, B1 => n61519, B2 => 
                           n4804, C1 => n61516, C2 => n53190, ZN => n14620);
   U8338 : OAI221_X1 port map( B1 => n1501, B2 => n61577, C1 => n1477, C2 => 
                           n61574, A => n14612, ZN => n14605);
   U8339 : AOI222_X1 port map( A1 => n61571, A2 => n5020, B1 => n61570, B2 => 
                           n5044, C1 => n61567, C2 => n52874, ZN => n14612);
   U8340 : OAI221_X1 port map( B1 => n4546, B2 => n61628, C1 => n4522, C2 => 
                           n61625, A => n14604, ZN => n14597);
   U8341 : AOI222_X1 port map( A1 => n61622, A2 => n4397, B1 => n61621, B2 => 
                           n4474, C1 => n61618, C2 => n4498, ZN => n14604);
   U8342 : OAI221_X1 port map( B1 => n3543, B2 => n61322, C1 => n3519, C2 => 
                           n61319, A => n14656, ZN => n14649);
   U8343 : AOI222_X1 port map( A1 => n61316, A2 => n53698, B1 => n61315, B2 => 
                           n53722, C1 => n61312, C2 => n53746, ZN => n14656);
   U8344 : OAI221_X1 port map( B1 => n3889, B2 => n61373, C1 => n3865, C2 => 
                           n61370, A => n14648, ZN => n14641);
   U8345 : AOI222_X1 port map( A1 => n61367, A2 => n53934, B1 => n61366, B2 => 
                           n53958, C1 => n61363, C2 => n53982, ZN => n14648);
   U8346 : OAI221_X1 port map( B1 => n2164, B2 => n61424, C1 => n2140, C2 => 
                           n61421, A => n14640, ZN => n14633);
   U8347 : AOI222_X1 port map( A1 => n61418, A2 => n54174, B1 => n61417, B2 => 
                           n54198, C1 => n61414, C2 => n54222, ZN => n14640);
   U8348 : OAI221_X1 port map( B1 => n4851, B2 => n61526, C1 => n3168, C2 => 
                           n61523, A => n14545, ZN => n14538);
   U8349 : AOI222_X1 port map( A1 => n61520, A2 => n53141, B1 => n61519, B2 => 
                           n4803, C1 => n61516, C2 => n53189, ZN => n14545);
   U8350 : OAI221_X1 port map( B1 => n1500, B2 => n61577, C1 => n1476, C2 => 
                           n61574, A => n14537, ZN => n14530);
   U8351 : AOI222_X1 port map( A1 => n61571, A2 => n5019, B1 => n61570, B2 => 
                           n5043, C1 => n61567, C2 => n52873, ZN => n14537);
   U8352 : OAI221_X1 port map( B1 => n4545, B2 => n61628, C1 => n4521, C2 => 
                           n61625, A => n14529, ZN => n14522);
   U8353 : AOI222_X1 port map( A1 => n61622, A2 => n4396, B1 => n61621, B2 => 
                           n4473, C1 => n61618, C2 => n4497, ZN => n14529);
   U8354 : OAI221_X1 port map( B1 => n3542, B2 => n61322, C1 => n3518, C2 => 
                           n61319, A => n14581, ZN => n14574);
   U8355 : AOI222_X1 port map( A1 => n61316, A2 => n53697, B1 => n61315, B2 => 
                           n53721, C1 => n61312, C2 => n53745, ZN => n14581);
   U8356 : OAI221_X1 port map( B1 => n3888, B2 => n61373, C1 => n3864, C2 => 
                           n61370, A => n14573, ZN => n14566);
   U8357 : AOI222_X1 port map( A1 => n61367, A2 => n53933, B1 => n61366, B2 => 
                           n53957, C1 => n61363, C2 => n53981, ZN => n14573);
   U8358 : OAI221_X1 port map( B1 => n2163, B2 => n61424, C1 => n2139, C2 => 
                           n61421, A => n14565, ZN => n14558);
   U8359 : AOI222_X1 port map( A1 => n61418, A2 => n54173, B1 => n61417, B2 => 
                           n54197, C1 => n61414, C2 => n54221, ZN => n14565);
   U8360 : OAI221_X1 port map( B1 => n4850, B2 => n61526, C1 => n3167, C2 => 
                           n61523, A => n14470, ZN => n14463);
   U8361 : AOI222_X1 port map( A1 => n61520, A2 => n53140, B1 => n61519, B2 => 
                           n4802, C1 => n61516, C2 => n53188, ZN => n14470);
   U8362 : OAI221_X1 port map( B1 => n1499, B2 => n61577, C1 => n1475, C2 => 
                           n61574, A => n14462, ZN => n14455);
   U8363 : AOI222_X1 port map( A1 => n61571, A2 => n5018, B1 => n61570, B2 => 
                           n5042, C1 => n61567, C2 => n52872, ZN => n14462);
   U8364 : OAI221_X1 port map( B1 => n4544, B2 => n61628, C1 => n4520, C2 => 
                           n61625, A => n14454, ZN => n14447);
   U8365 : AOI222_X1 port map( A1 => n61622, A2 => n4395, B1 => n61621, B2 => 
                           n4472, C1 => n61618, C2 => n4496, ZN => n14454);
   U8366 : OAI221_X1 port map( B1 => n3541, B2 => n61322, C1 => n3517, C2 => 
                           n61319, A => n14506, ZN => n14499);
   U8367 : AOI222_X1 port map( A1 => n61316, A2 => n53696, B1 => n61315, B2 => 
                           n53720, C1 => n61312, C2 => n53744, ZN => n14506);
   U8368 : OAI221_X1 port map( B1 => n3887, B2 => n61373, C1 => n3863, C2 => 
                           n61370, A => n14498, ZN => n14491);
   U8369 : AOI222_X1 port map( A1 => n61367, A2 => n53932, B1 => n61366, B2 => 
                           n53956, C1 => n61363, C2 => n53980, ZN => n14498);
   U8370 : OAI221_X1 port map( B1 => n2162, B2 => n61424, C1 => n2138, C2 => 
                           n61421, A => n14490, ZN => n14483);
   U8371 : AOI222_X1 port map( A1 => n61418, A2 => n54172, B1 => n61417, B2 => 
                           n54196, C1 => n61414, C2 => n54220, ZN => n14490);
   U8372 : OAI22_X1 port map( A1 => n62125, A2 => n396, B1 => n62118, B2 => 
                           n60969, ZN => n10000);
   U8373 : OAI22_X1 port map( A1 => n62125, A2 => n395, B1 => n62117, B2 => 
                           n60983, ZN => n10001);
   U8374 : OAI22_X1 port map( A1 => n62124, A2 => n394, B1 => n62118, B2 => 
                           n60997, ZN => n10002);
   U8375 : OAI22_X1 port map( A1 => n62124, A2 => n393, B1 => n62117, B2 => 
                           n61011, ZN => n10003);
   U8376 : OAI22_X1 port map( A1 => n62124, A2 => n392, B1 => n62118, B2 => 
                           n61025, ZN => n10004);
   U8377 : OAI22_X1 port map( A1 => n62124, A2 => n391, B1 => n62117, B2 => 
                           n61039, ZN => n10005);
   U8378 : OAI22_X1 port map( A1 => n62124, A2 => n390, B1 => n62118, B2 => 
                           n61053, ZN => n10006);
   U8379 : OAI22_X1 port map( A1 => n62123, A2 => n389, B1 => n62117, B2 => 
                           n61067, ZN => n10007);
   U8380 : AOI22_X1 port map( A1 => n16429, A2 => n61929, B1 => n16421, B2 => 
                           n61926, ZN => n6030);
   U8381 : AOI22_X1 port map( A1 => n15918, A2 => n61917, B1 => n15919, B2 => 
                           n61914, ZN => n6031);
   U8382 : AOI22_X1 port map( A1 => n16144, A2 => n61896, B1 => n16143, B2 => 
                           n61893, ZN => n6041);
   U8383 : AOI22_X1 port map( A1 => n51623, A2 => n61944, B1 => n51615, B2 => 
                           n61939, ZN => n6022);
   U8384 : AOI22_X1 port map( A1 => n52591, A2 => n61812, B1 => n52607, B2 => 
                           n61809, ZN => n6097);
   U8385 : AOI22_X1 port map( A1 => n387, A2 => n61806, B1 => n379, B2 => 
                           n61803, ZN => n6098);
   U8386 : AOI22_X1 port map( A1 => n355, A2 => n61794, B1 => n347, B2 => 
                           n61791, ZN => n6099);
   U8387 : AOI22_X1 port map( A1 => n16469, A2 => n61755, B1 => n15675, B2 => 
                           n61752, ZN => n6109);
   U8388 : AOI22_X1 port map( A1 => n51727, A2 => n61833, B1 => n51719, B2 => 
                           n61830, ZN => n6083);
   U8389 : AOI22_X1 port map( A1 => n451, A2 => n61842, B1 => n443, B2 => 
                           n61839, ZN => n6075);
   U8390 : AOI22_X1 port map( A1 => n16430, A2 => n61929, B1 => n16422, B2 => 
                           n61926, ZN => n5949);
   U8391 : AOI22_X1 port map( A1 => n15922, A2 => n61917, B1 => n15947, B2 => 
                           n61914, ZN => n5950);
   U8392 : AOI22_X1 port map( A1 => n16146, A2 => n61896, B1 => n16145, B2 => 
                           n61893, ZN => n5957);
   U8393 : AOI22_X1 port map( A1 => n51622, A2 => n61944, B1 => n51614, B2 => 
                           n61939, ZN => n5943);
   U8394 : AOI22_X1 port map( A1 => n52590, A2 => n61812, B1 => n52606, B2 => 
                           n61809, ZN => n5993);
   U8395 : AOI22_X1 port map( A1 => n386, A2 => n61806, B1 => n378, B2 => 
                           n61803, ZN => n5994);
   U8396 : AOI22_X1 port map( A1 => n354, A2 => n61794, B1 => n346, B2 => 
                           n61791, ZN => n5995);
   U8397 : AOI22_X1 port map( A1 => n16470, A2 => n61755, B1 => n15678, B2 => 
                           n61752, ZN => n6003);
   U8398 : AOI22_X1 port map( A1 => n51726, A2 => n61833, B1 => n51718, B2 => 
                           n61830, ZN => n5985);
   U8399 : AOI22_X1 port map( A1 => n450, A2 => n61842, B1 => n442, B2 => 
                           n61839, ZN => n5979);
   U8400 : AOI22_X1 port map( A1 => n16431, A2 => n61929, B1 => n16423, B2 => 
                           n61926, ZN => n5874);
   U8401 : AOI22_X1 port map( A1 => n15950, A2 => n61917, B1 => n15951, B2 => 
                           n61914, ZN => n5875);
   U8402 : AOI22_X1 port map( A1 => n16148, A2 => n61896, B1 => n16147, B2 => 
                           n61893, ZN => n5882);
   U8403 : AOI22_X1 port map( A1 => n51621, A2 => n61944, B1 => n51613, B2 => 
                           n61939, ZN => n5868);
   U8404 : AOI22_X1 port map( A1 => n52589, A2 => n61812, B1 => n52605, B2 => 
                           n61809, ZN => n5918);
   U8405 : AOI22_X1 port map( A1 => n385, A2 => n61806, B1 => n377, B2 => 
                           n61803, ZN => n5919);
   U8406 : AOI22_X1 port map( A1 => n353, A2 => n61794, B1 => n345, B2 => 
                           n61791, ZN => n5920);
   U8407 : AOI22_X1 port map( A1 => n16471, A2 => n61755, B1 => n15681, B2 => 
                           n61752, ZN => n5928);
   U8408 : AOI22_X1 port map( A1 => n51725, A2 => n61833, B1 => n51717, B2 => 
                           n61830, ZN => n5910);
   U8409 : AOI22_X1 port map( A1 => n449, A2 => n61842, B1 => n441, B2 => 
                           n61839, ZN => n5904);
   U8410 : AOI22_X1 port map( A1 => n16432, A2 => n61929, B1 => n16424, B2 => 
                           n61926, ZN => n5799);
   U8411 : AOI22_X1 port map( A1 => n15954, A2 => n61917, B1 => n15955, B2 => 
                           n61914, ZN => n5800);
   U8412 : AOI22_X1 port map( A1 => n16150, A2 => n61896, B1 => n16149, B2 => 
                           n61893, ZN => n5807);
   U8413 : AOI22_X1 port map( A1 => n51620, A2 => n61944, B1 => n51612, B2 => 
                           n61939, ZN => n5793);
   U8414 : AOI22_X1 port map( A1 => n52588, A2 => n61812, B1 => n52604, B2 => 
                           n61809, ZN => n5843);
   U8415 : AOI22_X1 port map( A1 => n384, A2 => n61806, B1 => n376, B2 => 
                           n61803, ZN => n5844);
   U8416 : AOI22_X1 port map( A1 => n352, A2 => n61794, B1 => n344, B2 => 
                           n61791, ZN => n5845);
   U8417 : AOI22_X1 port map( A1 => n16472, A2 => n61755, B1 => n15684, B2 => 
                           n61752, ZN => n5853);
   U8418 : AOI22_X1 port map( A1 => n51724, A2 => n61833, B1 => n51716, B2 => 
                           n61830, ZN => n5835);
   U8419 : AOI22_X1 port map( A1 => n448, A2 => n61842, B1 => n440, B2 => 
                           n61839, ZN => n5829);
   U8420 : AOI22_X1 port map( A1 => n16433, A2 => n61929, B1 => n16425, B2 => 
                           n61926, ZN => n5724);
   U8421 : AOI22_X1 port map( A1 => n15958, A2 => n61917, B1 => n15959, B2 => 
                           n61914, ZN => n5725);
   U8422 : AOI22_X1 port map( A1 => n16152, A2 => n61896, B1 => n16151, B2 => 
                           n61893, ZN => n5732);
   U8423 : AOI22_X1 port map( A1 => n51619, A2 => n61944, B1 => n51611, B2 => 
                           n61939, ZN => n5718);
   U8424 : AOI22_X1 port map( A1 => n52587, A2 => n61812, B1 => n52603, B2 => 
                           n61809, ZN => n5768);
   U8425 : AOI22_X1 port map( A1 => n383, A2 => n61806, B1 => n375, B2 => 
                           n61803, ZN => n5769);
   U8426 : AOI22_X1 port map( A1 => n351, A2 => n61794, B1 => n343, B2 => 
                           n61791, ZN => n5770);
   U8427 : AOI22_X1 port map( A1 => n16473, A2 => n61755, B1 => n15663, B2 => 
                           n61752, ZN => n5778);
   U8428 : AOI22_X1 port map( A1 => n51723, A2 => n61833, B1 => n51715, B2 => 
                           n61830, ZN => n5760);
   U8429 : AOI22_X1 port map( A1 => n447, A2 => n61842, B1 => n439, B2 => 
                           n61839, ZN => n5754);
   U8430 : AOI22_X1 port map( A1 => n16434, A2 => n61929, B1 => n16426, B2 => 
                           n61926, ZN => n5649);
   U8431 : AOI22_X1 port map( A1 => n15962, A2 => n61917, B1 => n15963, B2 => 
                           n61914, ZN => n5650);
   U8432 : AOI22_X1 port map( A1 => n16154, A2 => n61896, B1 => n16153, B2 => 
                           n61893, ZN => n5657);
   U8433 : AOI22_X1 port map( A1 => n51618, A2 => n61944, B1 => n51610, B2 => 
                           n61939, ZN => n5643);
   U8434 : AOI22_X1 port map( A1 => n52586, A2 => n61812, B1 => n52602, B2 => 
                           n61809, ZN => n5693);
   U8435 : AOI22_X1 port map( A1 => n382, A2 => n61806, B1 => n374, B2 => 
                           n61803, ZN => n5694);
   U8436 : AOI22_X1 port map( A1 => n350, A2 => n61794, B1 => n342, B2 => 
                           n61791, ZN => n5695);
   U8437 : AOI22_X1 port map( A1 => n16474, A2 => n61755, B1 => n15666, B2 => 
                           n61752, ZN => n5703);
   U8438 : AOI22_X1 port map( A1 => n51722, A2 => n61833, B1 => n51714, B2 => 
                           n61830, ZN => n5685);
   U8439 : AOI22_X1 port map( A1 => n446, A2 => n61842, B1 => n438, B2 => 
                           n61839, ZN => n5679);
   U8440 : AOI22_X1 port map( A1 => n16435, A2 => n61929, B1 => n16427, B2 => 
                           n61926, ZN => n5574);
   U8441 : AOI22_X1 port map( A1 => n15966, A2 => n61917, B1 => n15967, B2 => 
                           n61914, ZN => n5575);
   U8442 : AOI22_X1 port map( A1 => n16156, A2 => n61896, B1 => n16155, B2 => 
                           n61893, ZN => n5582);
   U8443 : AOI22_X1 port map( A1 => n51617, A2 => n61944, B1 => n51609, B2 => 
                           n61939, ZN => n5568);
   U8444 : AOI22_X1 port map( A1 => n52585, A2 => n61812, B1 => n52601, B2 => 
                           n61809, ZN => n5618);
   U8445 : AOI22_X1 port map( A1 => n381, A2 => n61806, B1 => n373, B2 => 
                           n61803, ZN => n5619);
   U8446 : AOI22_X1 port map( A1 => n349, A2 => n61794, B1 => n341, B2 => 
                           n61791, ZN => n5620);
   U8447 : AOI22_X1 port map( A1 => n16475, A2 => n61755, B1 => n15669, B2 => 
                           n61752, ZN => n5628);
   U8448 : AOI22_X1 port map( A1 => n51721, A2 => n61833, B1 => n51713, B2 => 
                           n61830, ZN => n5610);
   U8449 : AOI22_X1 port map( A1 => n445, A2 => n61842, B1 => n437, B2 => 
                           n61839, ZN => n5604);
   U8450 : AOI22_X1 port map( A1 => n16436, A2 => n61929, B1 => n16428, B2 => 
                           n61926, ZN => n5407);
   U8451 : AOI22_X1 port map( A1 => n15970, A2 => n61917, B1 => n15971, B2 => 
                           n61914, ZN => n5412);
   U8452 : AOI22_X1 port map( A1 => n16158, A2 => n61896, B1 => n16157, B2 => 
                           n61893, ZN => n5429);
   U8453 : AOI22_X1 port map( A1 => n51616, A2 => n61944, B1 => n51608, B2 => 
                           n61939, ZN => n5394);
   U8454 : AOI22_X1 port map( A1 => n52584, A2 => n61812, B1 => n52600, B2 => 
                           n61809, ZN => n5513);
   U8455 : AOI22_X1 port map( A1 => n380, A2 => n61806, B1 => n372, B2 => 
                           n61803, ZN => n5518);
   U8456 : AOI22_X1 port map( A1 => n348, A2 => n61794, B1 => n340, B2 => 
                           n61791, ZN => n5523);
   U8457 : AOI22_X1 port map( A1 => n16476, A2 => n61755, B1 => n15672, B2 => 
                           n61752, ZN => n5546);
   U8458 : AOI22_X1 port map( A1 => n51720, A2 => n61833, B1 => n51712, B2 => 
                           n61830, ZN => n5494);
   U8459 : AOI22_X1 port map( A1 => n444, A2 => n61842, B1 => n436, B2 => 
                           n61839, ZN => n5481);
   U8460 : OAI22_X1 port map( A1 => n62123, A2 => n1279, B1 => n62118, B2 => 
                           n61081, ZN => n10008);
   U8461 : OAI22_X1 port map( A1 => n62123, A2 => n1278, B1 => n62118, B2 => 
                           n61095, ZN => n10009);
   U8462 : OAI22_X1 port map( A1 => n62123, A2 => n1277, B1 => n62118, B2 => 
                           n61109, ZN => n10010);
   U8463 : OAI22_X1 port map( A1 => n62123, A2 => n1276, B1 => n62118, B2 => 
                           n61123, ZN => n10011);
   U8464 : OAI22_X1 port map( A1 => n62122, A2 => n1275, B1 => n62118, B2 => 
                           n61137, ZN => n10012);
   U8465 : OAI22_X1 port map( A1 => n62122, A2 => n1274, B1 => n62118, B2 => 
                           n61151, ZN => n10013);
   U8466 : OAI22_X1 port map( A1 => n62122, A2 => n1273, B1 => n62118, B2 => 
                           n61165, ZN => n10014);
   U8467 : OAI22_X1 port map( A1 => n62122, A2 => n1272, B1 => n62118, B2 => 
                           n61179, ZN => n10015);
   U8468 : OAI22_X1 port map( A1 => n62122, A2 => n1271, B1 => n62118, B2 => 
                           n61193, ZN => n10016);
   U8469 : OAI22_X1 port map( A1 => n62121, A2 => n1270, B1 => n62118, B2 => 
                           n61207, ZN => n10017);
   U8470 : OAI22_X1 port map( A1 => n62121, A2 => n1269, B1 => n62118, B2 => 
                           n61221, ZN => n10018);
   U8471 : OAI22_X1 port map( A1 => n62121, A2 => n1268, B1 => n62118, B2 => 
                           n61235, ZN => n10019);
   U8472 : OAI22_X1 port map( A1 => n62121, A2 => n1267, B1 => n62117, B2 => 
                           n61258, ZN => n10020);
   U8473 : OAI22_X1 port map( A1 => n3929, A2 => n15286, B1 => n59749, B2 => 
                           n61976, ZN => n10021);
   U8474 : OAI22_X1 port map( A1 => n3928, A2 => n15286, B1 => n59749, B2 => 
                           n61990, ZN => n10022);
   U8475 : OAI22_X1 port map( A1 => n3927, A2 => n15286, B1 => n59749, B2 => 
                           n62004, ZN => n10023);
   U8476 : OAI22_X1 port map( A1 => n99, A2 => n15286, B1 => n59749, B2 => 
                           n62018, ZN => n10024);
   U8477 : OAI22_X1 port map( A1 => n98, A2 => n15286, B1 => n59750, B2 => 
                           n62032, ZN => n10025);
   U8478 : OAI22_X1 port map( A1 => n97, A2 => n15286, B1 => n59750, B2 => 
                           n62046, ZN => n10026);
   U8479 : OAI22_X1 port map( A1 => n96, A2 => n59748, B1 => n59750, B2 => 
                           n62060, ZN => n10027);
   U8480 : OAI22_X1 port map( A1 => n95, A2 => n59748, B1 => n59750, B2 => 
                           n62074, ZN => n10028);
   U8481 : OAI22_X1 port map( A1 => n94, A2 => n59748, B1 => n59751, B2 => 
                           n62088, ZN => n10029);
   U8482 : OAI22_X1 port map( A1 => n93, A2 => n59748, B1 => n59751, B2 => 
                           n62102, ZN => n10030);
   U8483 : OAI22_X1 port map( A1 => n92, A2 => n59748, B1 => n59751, B2 => 
                           n62116, ZN => n10031);
   U8484 : OAI22_X1 port map( A1 => n62121, A2 => n1290, B1 => n62117, B2 => 
                           n61976, ZN => n9989);
   U8485 : OAI22_X1 port map( A1 => n62120, A2 => n1289, B1 => n62117, B2 => 
                           n61990, ZN => n9990);
   U8486 : OAI22_X1 port map( A1 => n62120, A2 => n1288, B1 => n62117, B2 => 
                           n62004, ZN => n9991);
   U8487 : OAI22_X1 port map( A1 => n62120, A2 => n1287, B1 => n62117, B2 => 
                           n62018, ZN => n9992);
   U8488 : OAI22_X1 port map( A1 => n62120, A2 => n1286, B1 => n62117, B2 => 
                           n62032, ZN => n9993);
   U8489 : OAI22_X1 port map( A1 => n62120, A2 => n1285, B1 => n62117, B2 => 
                           n62046, ZN => n9994);
   U8490 : OAI22_X1 port map( A1 => n62119, A2 => n1284, B1 => n62117, B2 => 
                           n62060, ZN => n9995);
   U8491 : OAI22_X1 port map( A1 => n62119, A2 => n1283, B1 => n62117, B2 => 
                           n62074, ZN => n9996);
   U8492 : OAI22_X1 port map( A1 => n62119, A2 => n1282, B1 => n62117, B2 => 
                           n62088, ZN => n9997);
   U8493 : OAI22_X1 port map( A1 => n62119, A2 => n1281, B1 => n62117, B2 => 
                           n62102, ZN => n9998);
   U8494 : OAI22_X1 port map( A1 => n62119, A2 => n1280, B1 => n62117, B2 => 
                           n62116, ZN => n9999);
   U8495 : OAI22_X1 port map( A1 => n59936, A2 => n61163, B1 => n15177, B2 => 
                           n59930, ZN => n10686);
   U8496 : OAI22_X1 port map( A1 => n59936, A2 => n61177, B1 => n15176, B2 => 
                           n59930, ZN => n10687);
   U8497 : OAI22_X1 port map( A1 => n59936, A2 => n61191, B1 => n15175, B2 => 
                           n59930, ZN => n10688);
   U8498 : OAI22_X1 port map( A1 => n59936, A2 => n61205, B1 => n15174, B2 => 
                           n15249, ZN => n10689);
   U8499 : OAI22_X1 port map( A1 => n59936, A2 => n61219, B1 => n15173, B2 => 
                           n15249, ZN => n10690);
   U8500 : OAI22_X1 port map( A1 => n59937, A2 => n61233, B1 => n15172, B2 => 
                           n15249, ZN => n10691);
   U8501 : OAI22_X1 port map( A1 => n59937, A2 => n61256, B1 => n15171, B2 => 
                           n15249, ZN => n10692);
   U8502 : OAI22_X1 port map( A1 => n59926, A2 => n61149, B1 => n15210, B2 => 
                           n59921, ZN => n10653);
   U8503 : OAI22_X1 port map( A1 => n59927, A2 => n61163, B1 => n15209, B2 => 
                           n59921, ZN => n10654);
   U8504 : OAI22_X1 port map( A1 => n59927, A2 => n61177, B1 => n15208, B2 => 
                           n59921, ZN => n10655);
   U8505 : OAI22_X1 port map( A1 => n59927, A2 => n61191, B1 => n15207, B2 => 
                           n59921, ZN => n10656);
   U8506 : OAI22_X1 port map( A1 => n59927, A2 => n61205, B1 => n15206, B2 => 
                           n15250, ZN => n10657);
   U8507 : OAI22_X1 port map( A1 => n59927, A2 => n61219, B1 => n15205, B2 => 
                           n15250, ZN => n10658);
   U8508 : OAI22_X1 port map( A1 => n59928, A2 => n61233, B1 => n15204, B2 => 
                           n15250, ZN => n10659);
   U8509 : OAI22_X1 port map( A1 => n59928, A2 => n61256, B1 => n15203, B2 => 
                           n15250, ZN => n10660);
   U8510 : OAI22_X1 port map( A1 => n59873, A2 => n61206, B1 => n52507, B2 => 
                           n15258, ZN => n10465);
   U8511 : OAI22_X1 port map( A1 => n59873, A2 => n61220, B1 => n52506, B2 => 
                           n15258, ZN => n10466);
   U8512 : OAI22_X1 port map( A1 => n59874, A2 => n61234, B1 => n52505, B2 => 
                           n15258, ZN => n10467);
   U8513 : OAI22_X1 port map( A1 => n59874, A2 => n61257, B1 => n52504, B2 => 
                           n15258, ZN => n10468);
   U8514 : OAI22_X1 port map( A1 => n59863, A2 => n61150, B1 => n52503, B2 => 
                           n59858, ZN => n10429);
   U8515 : OAI22_X1 port map( A1 => n59864, A2 => n61164, B1 => n52502, B2 => 
                           n59858, ZN => n10430);
   U8516 : OAI22_X1 port map( A1 => n59864, A2 => n61178, B1 => n52501, B2 => 
                           n59858, ZN => n10431);
   U8517 : OAI22_X1 port map( A1 => n59864, A2 => n61192, B1 => n52500, B2 => 
                           n59858, ZN => n10432);
   U8518 : OAI22_X1 port map( A1 => n59864, A2 => n61206, B1 => n52499, B2 => 
                           n15260, ZN => n10433);
   U8519 : OAI22_X1 port map( A1 => n59864, A2 => n61220, B1 => n52498, B2 => 
                           n15260, ZN => n10434);
   U8520 : OAI22_X1 port map( A1 => n59865, A2 => n61234, B1 => n52497, B2 => 
                           n15260, ZN => n10435);
   U8521 : OAI22_X1 port map( A1 => n59865, A2 => n61257, B1 => n52496, B2 => 
                           n15260, ZN => n10436);
   U8522 : OAI22_X1 port map( A1 => n59836, A2 => n61150, B1 => n15306, B2 => 
                           n59831, ZN => n10333);
   U8523 : OAI22_X1 port map( A1 => n59837, A2 => n61164, B1 => n15305, B2 => 
                           n59831, ZN => n10334);
   U8524 : OAI22_X1 port map( A1 => n59837, A2 => n61178, B1 => n15304, B2 => 
                           n59831, ZN => n10335);
   U8525 : OAI22_X1 port map( A1 => n59837, A2 => n61192, B1 => n15303, B2 => 
                           n59831, ZN => n10336);
   U8526 : OAI22_X1 port map( A1 => n59837, A2 => n61206, B1 => n15302, B2 => 
                           n15266, ZN => n10337);
   U8527 : OAI22_X1 port map( A1 => n59837, A2 => n61220, B1 => n15301, B2 => 
                           n15266, ZN => n10338);
   U8528 : OAI22_X1 port map( A1 => n59838, A2 => n61234, B1 => n15300, B2 => 
                           n15266, ZN => n10339);
   U8529 : OAI22_X1 port map( A1 => n59838, A2 => n61257, B1 => n15299, B2 => 
                           n15266, ZN => n10340);
   U8530 : OAI22_X1 port map( A1 => n59827, A2 => n61150, B1 => n15338, B2 => 
                           n59822, ZN => n10301);
   U8531 : OAI22_X1 port map( A1 => n59828, A2 => n61164, B1 => n15337, B2 => 
                           n59822, ZN => n10302);
   U8532 : OAI22_X1 port map( A1 => n59828, A2 => n61178, B1 => n15336, B2 => 
                           n59822, ZN => n10303);
   U8533 : OAI22_X1 port map( A1 => n59828, A2 => n61192, B1 => n15335, B2 => 
                           n59822, ZN => n10304);
   U8534 : OAI22_X1 port map( A1 => n59828, A2 => n61206, B1 => n15334, B2 => 
                           n15267, ZN => n10305);
   U8535 : OAI22_X1 port map( A1 => n59828, A2 => n61220, B1 => n15333, B2 => 
                           n15267, ZN => n10306);
   U8536 : OAI22_X1 port map( A1 => n59829, A2 => n61234, B1 => n15332, B2 => 
                           n15267, ZN => n10307);
   U8537 : OAI22_X1 port map( A1 => n59829, A2 => n61257, B1 => n15331, B2 => 
                           n15267, ZN => n10308);
   U8538 : OAI22_X1 port map( A1 => n60619, A2 => n61143, B1 => n9754, B2 => 
                           n60614, ZN => n13117);
   U8539 : OAI22_X1 port map( A1 => n60620, A2 => n61157, B1 => n9753, B2 => 
                           n60614, ZN => n13118);
   U8540 : OAI22_X1 port map( A1 => n60620, A2 => n61171, B1 => n9752, B2 => 
                           n60614, ZN => n13119);
   U8541 : OAI22_X1 port map( A1 => n60620, A2 => n61185, B1 => n9751, B2 => 
                           n60614, ZN => n13120);
   U8542 : OAI22_X1 port map( A1 => n60620, A2 => n61199, B1 => n9750, B2 => 
                           n15153, ZN => n13121);
   U8543 : OAI22_X1 port map( A1 => n60620, A2 => n61213, B1 => n9749, B2 => 
                           n15153, ZN => n13122);
   U8544 : OAI22_X1 port map( A1 => n60621, A2 => n61227, B1 => n9748, B2 => 
                           n15153, ZN => n13123);
   U8545 : OAI22_X1 port map( A1 => n60621, A2 => n61250, B1 => n9747, B2 => 
                           n15153, ZN => n13124);
   U8546 : OAI22_X1 port map( A1 => n60610, A2 => n61143, B1 => n9786, B2 => 
                           n60605, ZN => n13085);
   U8547 : OAI22_X1 port map( A1 => n60611, A2 => n61157, B1 => n9785, B2 => 
                           n60605, ZN => n13086);
   U8548 : OAI22_X1 port map( A1 => n60611, A2 => n61171, B1 => n9784, B2 => 
                           n60605, ZN => n13087);
   U8549 : OAI22_X1 port map( A1 => n60611, A2 => n61185, B1 => n9783, B2 => 
                           n60605, ZN => n13088);
   U8550 : OAI22_X1 port map( A1 => n60611, A2 => n61199, B1 => n9782, B2 => 
                           n15154, ZN => n13089);
   U8551 : OAI22_X1 port map( A1 => n60611, A2 => n61213, B1 => n9781, B2 => 
                           n15154, ZN => n13090);
   U8552 : OAI22_X1 port map( A1 => n60612, A2 => n61227, B1 => n9780, B2 => 
                           n15154, ZN => n13091);
   U8553 : OAI22_X1 port map( A1 => n60612, A2 => n61250, B1 => n9779, B2 => 
                           n15154, ZN => n13092);
   U8554 : OAI22_X1 port map( A1 => n60583, A2 => n61143, B1 => n4256, B2 => 
                           n60578, ZN => n12989);
   U8555 : OAI22_X1 port map( A1 => n60584, A2 => n61157, B1 => n4255, B2 => 
                           n60578, ZN => n12990);
   U8556 : OAI22_X1 port map( A1 => n60584, A2 => n61171, B1 => n4254, B2 => 
                           n60578, ZN => n12991);
   U8557 : OAI22_X1 port map( A1 => n60584, A2 => n61185, B1 => n4253, B2 => 
                           n60578, ZN => n12992);
   U8558 : OAI22_X1 port map( A1 => n60584, A2 => n61199, B1 => n4252, B2 => 
                           n15157, ZN => n12993);
   U8559 : OAI22_X1 port map( A1 => n60584, A2 => n61213, B1 => n4251, B2 => 
                           n15157, ZN => n12994);
   U8560 : OAI22_X1 port map( A1 => n60585, A2 => n61227, B1 => n4250, B2 => 
                           n15157, ZN => n12995);
   U8561 : OAI22_X1 port map( A1 => n60585, A2 => n61250, B1 => n4249, B2 => 
                           n15157, ZN => n12996);
   U8562 : OAI22_X1 port map( A1 => n60574, A2 => n61143, B1 => n4248, B2 => 
                           n60569, ZN => n12957);
   U8563 : OAI22_X1 port map( A1 => n60575, A2 => n61157, B1 => n4247, B2 => 
                           n60569, ZN => n12958);
   U8564 : OAI22_X1 port map( A1 => n60575, A2 => n61171, B1 => n4246, B2 => 
                           n60569, ZN => n12959);
   U8565 : OAI22_X1 port map( A1 => n60575, A2 => n61185, B1 => n4245, B2 => 
                           n60569, ZN => n12960);
   U8566 : OAI22_X1 port map( A1 => n60575, A2 => n61199, B1 => n4244, B2 => 
                           n15158, ZN => n12961);
   U8567 : OAI22_X1 port map( A1 => n60575, A2 => n61213, B1 => n4243, B2 => 
                           n15158, ZN => n12962);
   U8568 : OAI22_X1 port map( A1 => n60576, A2 => n61227, B1 => n4242, B2 => 
                           n15158, ZN => n12963);
   U8569 : OAI22_X1 port map( A1 => n60576, A2 => n61250, B1 => n4241, B2 => 
                           n15158, ZN => n12964);
   U8570 : OAI22_X1 port map( A1 => n60466, A2 => n61144, B1 => n4211, B2 => 
                           n60461, ZN => n12573);
   U8571 : OAI22_X1 port map( A1 => n60467, A2 => n61158, B1 => n4210, B2 => 
                           n60461, ZN => n12574);
   U8572 : OAI22_X1 port map( A1 => n60467, A2 => n61172, B1 => n4209, B2 => 
                           n60461, ZN => n12575);
   U8573 : OAI22_X1 port map( A1 => n60467, A2 => n61186, B1 => n4208, B2 => 
                           n60461, ZN => n12576);
   U8574 : OAI22_X1 port map( A1 => n60467, A2 => n61200, B1 => n4207, B2 => 
                           n15178, ZN => n12577);
   U8575 : OAI22_X1 port map( A1 => n60467, A2 => n61214, B1 => n4206, B2 => 
                           n15178, ZN => n12578);
   U8576 : OAI22_X1 port map( A1 => n60468, A2 => n61228, B1 => n4205, B2 => 
                           n15178, ZN => n12579);
   U8577 : OAI22_X1 port map( A1 => n60468, A2 => n61251, B1 => n4204, B2 => 
                           n15178, ZN => n12580);
   U8578 : OAI22_X1 port map( A1 => n60457, A2 => n61144, B1 => n4203, B2 => 
                           n60452, ZN => n12541);
   U8579 : OAI22_X1 port map( A1 => n60458, A2 => n61158, B1 => n4202, B2 => 
                           n60452, ZN => n12542);
   U8580 : OAI22_X1 port map( A1 => n60458, A2 => n61172, B1 => n4201, B2 => 
                           n60452, ZN => n12543);
   U8581 : OAI22_X1 port map( A1 => n60458, A2 => n61186, B1 => n4200, B2 => 
                           n60452, ZN => n12544);
   U8582 : OAI22_X1 port map( A1 => n60458, A2 => n61200, B1 => n4199, B2 => 
                           n15179, ZN => n12545);
   U8583 : OAI22_X1 port map( A1 => n60458, A2 => n61214, B1 => n4198, B2 => 
                           n15179, ZN => n12546);
   U8584 : OAI22_X1 port map( A1 => n60459, A2 => n61228, B1 => n4197, B2 => 
                           n15179, ZN => n12547);
   U8585 : OAI22_X1 port map( A1 => n60459, A2 => n61251, B1 => n4196, B2 => 
                           n15179, ZN => n12548);
   U8586 : OAI22_X1 port map( A1 => n60412, A2 => n61145, B1 => n4195, B2 => 
                           n60407, ZN => n12381);
   U8587 : OAI22_X1 port map( A1 => n60413, A2 => n61159, B1 => n4194, B2 => 
                           n60407, ZN => n12382);
   U8588 : OAI22_X1 port map( A1 => n60413, A2 => n61173, B1 => n4193, B2 => 
                           n60407, ZN => n12383);
   U8589 : OAI22_X1 port map( A1 => n60413, A2 => n61187, B1 => n4192, B2 => 
                           n60407, ZN => n12384);
   U8590 : OAI22_X1 port map( A1 => n60413, A2 => n61201, B1 => n4191, B2 => 
                           n15184, ZN => n12385);
   U8591 : OAI22_X1 port map( A1 => n60413, A2 => n61215, B1 => n4190, B2 => 
                           n15184, ZN => n12386);
   U8592 : OAI22_X1 port map( A1 => n60414, A2 => n61229, B1 => n4189, B2 => 
                           n15184, ZN => n12387);
   U8593 : OAI22_X1 port map( A1 => n60414, A2 => n61252, B1 => n4188, B2 => 
                           n15184, ZN => n12388);
   U8594 : OAI22_X1 port map( A1 => n60403, A2 => n61145, B1 => n4187, B2 => 
                           n60398, ZN => n12349);
   U8595 : OAI22_X1 port map( A1 => n60404, A2 => n61159, B1 => n4186, B2 => 
                           n60398, ZN => n12350);
   U8596 : OAI22_X1 port map( A1 => n60404, A2 => n61173, B1 => n4185, B2 => 
                           n60398, ZN => n12351);
   U8597 : OAI22_X1 port map( A1 => n60404, A2 => n61187, B1 => n4184, B2 => 
                           n60398, ZN => n12352);
   U8598 : OAI22_X1 port map( A1 => n60404, A2 => n61201, B1 => n4183, B2 => 
                           n15185, ZN => n12353);
   U8599 : OAI22_X1 port map( A1 => n60404, A2 => n61215, B1 => n4182, B2 => 
                           n15185, ZN => n12354);
   U8600 : OAI22_X1 port map( A1 => n60405, A2 => n61229, B1 => n4181, B2 => 
                           n15185, ZN => n12355);
   U8601 : OAI22_X1 port map( A1 => n60405, A2 => n61252, B1 => n4180, B2 => 
                           n15185, ZN => n12356);
   U8602 : OAI22_X1 port map( A1 => n60943, A2 => n61140, B1 => n51647, B2 => 
                           n60938, ZN => n14269);
   U8603 : OAI22_X1 port map( A1 => n60944, A2 => n61154, B1 => n51646, B2 => 
                           n60938, ZN => n14270);
   U8604 : OAI22_X1 port map( A1 => n60944, A2 => n61168, B1 => n51645, B2 => 
                           n60938, ZN => n14271);
   U8605 : OAI22_X1 port map( A1 => n60944, A2 => n61182, B1 => n51644, B2 => 
                           n60938, ZN => n14272);
   U8606 : OAI22_X1 port map( A1 => n60944, A2 => n61196, B1 => n51643, B2 => 
                           n15098, ZN => n14273);
   U8607 : OAI22_X1 port map( A1 => n60944, A2 => n61210, B1 => n51642, B2 => 
                           n15098, ZN => n14274);
   U8608 : OAI22_X1 port map( A1 => n60945, A2 => n61224, B1 => n51641, B2 => 
                           n15098, ZN => n14275);
   U8609 : OAI22_X1 port map( A1 => n60945, A2 => n61247, B1 => n51640, B2 => 
                           n15098, ZN => n14276);
   U8610 : OAI22_X1 port map( A1 => n60934, A2 => n61140, B1 => n51639, B2 => 
                           n60929, ZN => n14237);
   U8611 : OAI22_X1 port map( A1 => n60935, A2 => n61154, B1 => n51638, B2 => 
                           n60929, ZN => n14238);
   U8612 : OAI22_X1 port map( A1 => n60935, A2 => n61168, B1 => n51637, B2 => 
                           n60929, ZN => n14239);
   U8613 : OAI22_X1 port map( A1 => n60935, A2 => n61182, B1 => n51636, B2 => 
                           n60929, ZN => n14240);
   U8614 : OAI22_X1 port map( A1 => n60935, A2 => n61196, B1 => n51635, B2 => 
                           n15100, ZN => n14241);
   U8615 : OAI22_X1 port map( A1 => n60935, A2 => n61210, B1 => n51634, B2 => 
                           n15100, ZN => n14242);
   U8616 : OAI22_X1 port map( A1 => n60936, A2 => n61224, B1 => n51633, B2 => 
                           n15100, ZN => n14243);
   U8617 : OAI22_X1 port map( A1 => n60936, A2 => n61247, B1 => n51632, B2 => 
                           n15100, ZN => n14244);
   U8618 : OAI22_X1 port map( A1 => n60835, A2 => n61141, B1 => n4115, B2 => 
                           n60830, ZN => n13885);
   U8619 : OAI22_X1 port map( A1 => n60836, A2 => n61155, B1 => n4114, B2 => 
                           n60830, ZN => n13886);
   U8620 : OAI22_X1 port map( A1 => n60836, A2 => n61169, B1 => n4113, B2 => 
                           n60830, ZN => n13887);
   U8621 : OAI22_X1 port map( A1 => n60836, A2 => n61183, B1 => n4112, B2 => 
                           n60830, ZN => n13888);
   U8622 : OAI22_X1 port map( A1 => n60836, A2 => n61197, B1 => n4111, B2 => 
                           n15122, ZN => n13889);
   U8623 : OAI22_X1 port map( A1 => n60836, A2 => n61211, B1 => n4110, B2 => 
                           n15122, ZN => n13890);
   U8624 : OAI22_X1 port map( A1 => n60837, A2 => n61225, B1 => n4109, B2 => 
                           n15122, ZN => n13891);
   U8625 : OAI22_X1 port map( A1 => n60837, A2 => n61248, B1 => n4108, B2 => 
                           n15122, ZN => n13892);
   U8626 : OAI22_X1 port map( A1 => n60826, A2 => n61141, B1 => n4107, B2 => 
                           n60821, ZN => n13853);
   U8627 : OAI22_X1 port map( A1 => n60827, A2 => n61155, B1 => n4106, B2 => 
                           n60821, ZN => n13854);
   U8628 : OAI22_X1 port map( A1 => n60827, A2 => n61169, B1 => n4105, B2 => 
                           n60821, ZN => n13855);
   U8629 : OAI22_X1 port map( A1 => n60827, A2 => n61183, B1 => n4104, B2 => 
                           n60821, ZN => n13856);
   U8630 : OAI22_X1 port map( A1 => n60827, A2 => n61197, B1 => n4103, B2 => 
                           n15124, ZN => n13857);
   U8631 : OAI22_X1 port map( A1 => n60827, A2 => n61211, B1 => n4102, B2 => 
                           n15124, ZN => n13858);
   U8632 : OAI22_X1 port map( A1 => n60828, A2 => n61225, B1 => n4101, B2 => 
                           n15124, ZN => n13859);
   U8633 : OAI22_X1 port map( A1 => n60828, A2 => n61248, B1 => n4100, B2 => 
                           n15124, ZN => n13860);
   U8634 : OAI22_X1 port map( A1 => n60376, A2 => n61145, B1 => n52751, B2 => 
                           n60371, ZN => n12253);
   U8635 : OAI22_X1 port map( A1 => n60377, A2 => n61159, B1 => n52750, B2 => 
                           n60371, ZN => n12254);
   U8636 : OAI22_X1 port map( A1 => n60377, A2 => n61173, B1 => n52749, B2 => 
                           n60371, ZN => n12255);
   U8637 : OAI22_X1 port map( A1 => n60377, A2 => n61187, B1 => n52748, B2 => 
                           n60371, ZN => n12256);
   U8638 : OAI22_X1 port map( A1 => n60377, A2 => n61201, B1 => n52747, B2 => 
                           n15189, ZN => n12257);
   U8639 : OAI22_X1 port map( A1 => n60377, A2 => n61215, B1 => n52746, B2 => 
                           n15189, ZN => n12258);
   U8640 : OAI22_X1 port map( A1 => n60378, A2 => n61229, B1 => n52745, B2 => 
                           n15189, ZN => n12259);
   U8641 : OAI22_X1 port map( A1 => n60378, A2 => n61252, B1 => n52744, B2 => 
                           n15189, ZN => n12260);
   U8642 : OAI22_X1 port map( A1 => n60367, A2 => n61145, B1 => n52743, B2 => 
                           n60362, ZN => n12221);
   U8643 : OAI22_X1 port map( A1 => n60368, A2 => n61159, B1 => n52742, B2 => 
                           n60362, ZN => n12222);
   U8644 : OAI22_X1 port map( A1 => n60368, A2 => n61173, B1 => n52741, B2 => 
                           n60362, ZN => n12223);
   U8645 : OAI22_X1 port map( A1 => n60368, A2 => n61187, B1 => n52740, B2 => 
                           n60362, ZN => n12224);
   U8646 : OAI22_X1 port map( A1 => n60368, A2 => n61201, B1 => n52739, B2 => 
                           n15190, ZN => n12225);
   U8647 : OAI22_X1 port map( A1 => n60368, A2 => n61215, B1 => n52738, B2 => 
                           n15190, ZN => n12226);
   U8648 : OAI22_X1 port map( A1 => n60369, A2 => n61229, B1 => n52737, B2 => 
                           n15190, ZN => n12227);
   U8649 : OAI22_X1 port map( A1 => n60369, A2 => n61252, B1 => n52736, B2 => 
                           n15190, ZN => n12228);
   U8650 : OAI22_X1 port map( A1 => n60358, A2 => n61145, B1 => n52735, B2 => 
                           n60353, ZN => n12189);
   U8651 : OAI22_X1 port map( A1 => n60359, A2 => n61159, B1 => n52734, B2 => 
                           n60353, ZN => n12190);
   U8652 : OAI22_X1 port map( A1 => n60359, A2 => n61173, B1 => n52733, B2 => 
                           n60353, ZN => n12191);
   U8653 : OAI22_X1 port map( A1 => n60359, A2 => n61187, B1 => n52732, B2 => 
                           n60353, ZN => n12192);
   U8654 : OAI22_X1 port map( A1 => n60359, A2 => n61201, B1 => n52731, B2 => 
                           n15191, ZN => n12193);
   U8655 : OAI22_X1 port map( A1 => n60359, A2 => n61215, B1 => n52730, B2 => 
                           n15191, ZN => n12194);
   U8656 : OAI22_X1 port map( A1 => n60360, A2 => n61229, B1 => n52729, B2 => 
                           n15191, ZN => n12195);
   U8657 : OAI22_X1 port map( A1 => n60360, A2 => n61252, B1 => n52728, B2 => 
                           n15191, ZN => n12196);
   U8658 : OAI22_X1 port map( A1 => n60223, A2 => n61146, B1 => n52679, B2 => 
                           n60218, ZN => n11709);
   U8659 : OAI22_X1 port map( A1 => n60224, A2 => n61160, B1 => n52678, B2 => 
                           n60218, ZN => n11710);
   U8660 : OAI22_X1 port map( A1 => n60224, A2 => n61174, B1 => n52677, B2 => 
                           n60218, ZN => n11711);
   U8661 : OAI22_X1 port map( A1 => n60224, A2 => n61188, B1 => n52676, B2 => 
                           n60218, ZN => n11712);
   U8662 : OAI22_X1 port map( A1 => n60224, A2 => n61202, B1 => n52675, B2 => 
                           n15215, ZN => n11713);
   U8663 : OAI22_X1 port map( A1 => n60224, A2 => n61216, B1 => n52674, B2 => 
                           n15215, ZN => n11714);
   U8664 : OAI22_X1 port map( A1 => n60225, A2 => n61230, B1 => n52673, B2 => 
                           n15215, ZN => n11715);
   U8665 : OAI22_X1 port map( A1 => n60225, A2 => n61253, B1 => n52672, B2 => 
                           n15215, ZN => n11716);
   U8666 : OAI22_X1 port map( A1 => n60214, A2 => n61146, B1 => n52671, B2 => 
                           n60209, ZN => n11677);
   U8667 : OAI22_X1 port map( A1 => n60215, A2 => n61160, B1 => n52670, B2 => 
                           n60209, ZN => n11678);
   U8668 : OAI22_X1 port map( A1 => n60215, A2 => n61174, B1 => n52669, B2 => 
                           n60209, ZN => n11679);
   U8669 : OAI22_X1 port map( A1 => n60215, A2 => n61188, B1 => n52668, B2 => 
                           n60209, ZN => n11680);
   U8670 : OAI22_X1 port map( A1 => n60215, A2 => n61202, B1 => n52667, B2 => 
                           n15216, ZN => n11681);
   U8671 : OAI22_X1 port map( A1 => n60215, A2 => n61216, B1 => n52666, B2 => 
                           n15216, ZN => n11682);
   U8672 : OAI22_X1 port map( A1 => n60216, A2 => n61230, B1 => n52665, B2 => 
                           n15216, ZN => n11683);
   U8673 : OAI22_X1 port map( A1 => n60216, A2 => n61253, B1 => n52664, B2 => 
                           n15216, ZN => n11684);
   U8674 : OAI22_X1 port map( A1 => n60718, A2 => n61142, B1 => n9610, B2 => 
                           n60713, ZN => n13469);
   U8675 : OAI22_X1 port map( A1 => n60719, A2 => n61156, B1 => n9609, B2 => 
                           n60713, ZN => n13470);
   U8676 : OAI22_X1 port map( A1 => n60719, A2 => n61170, B1 => n9608, B2 => 
                           n60713, ZN => n13471);
   U8677 : OAI22_X1 port map( A1 => n60719, A2 => n61184, B1 => n9607, B2 => 
                           n60713, ZN => n13472);
   U8678 : OAI22_X1 port map( A1 => n60719, A2 => n61198, B1 => n9606, B2 => 
                           n15140, ZN => n13473);
   U8679 : OAI22_X1 port map( A1 => n60719, A2 => n61212, B1 => n9605, B2 => 
                           n15140, ZN => n13474);
   U8680 : OAI22_X1 port map( A1 => n60720, A2 => n61226, B1 => n9604, B2 => 
                           n15140, ZN => n13475);
   U8681 : OAI22_X1 port map( A1 => n60720, A2 => n61249, B1 => n9603, B2 => 
                           n15140, ZN => n13476);
   U8682 : OAI22_X1 port map( A1 => n60709, A2 => n61142, B1 => n9618, B2 => 
                           n60704, ZN => n13437);
   U8683 : OAI22_X1 port map( A1 => n60710, A2 => n61156, B1 => n9617, B2 => 
                           n60704, ZN => n13438);
   U8684 : OAI22_X1 port map( A1 => n60710, A2 => n61170, B1 => n9616, B2 => 
                           n60704, ZN => n13439);
   U8685 : OAI22_X1 port map( A1 => n60710, A2 => n61184, B1 => n9615, B2 => 
                           n60704, ZN => n13440);
   U8686 : OAI22_X1 port map( A1 => n60710, A2 => n61198, B1 => n9614, B2 => 
                           n15141, ZN => n13441);
   U8687 : OAI22_X1 port map( A1 => n60710, A2 => n61212, B1 => n9613, B2 => 
                           n15141, ZN => n13442);
   U8688 : OAI22_X1 port map( A1 => n60711, A2 => n61226, B1 => n9612, B2 => 
                           n15141, ZN => n13443);
   U8689 : OAI22_X1 port map( A1 => n60711, A2 => n61249, B1 => n9611, B2 => 
                           n15141, ZN => n13444);
   U8690 : OAI22_X1 port map( A1 => n59809, A2 => n61150, B1 => n3947, B2 => 
                           n59804, ZN => n10237);
   U8691 : OAI22_X1 port map( A1 => n59810, A2 => n61164, B1 => n3946, B2 => 
                           n59804, ZN => n10238);
   U8692 : OAI22_X1 port map( A1 => n59810, A2 => n61178, B1 => n3945, B2 => 
                           n59804, ZN => n10239);
   U8693 : OAI22_X1 port map( A1 => n59810, A2 => n61192, B1 => n3944, B2 => 
                           n59804, ZN => n10240);
   U8694 : OAI22_X1 port map( A1 => n59810, A2 => n61206, B1 => n3943, B2 => 
                           n15269, ZN => n10241);
   U8695 : OAI22_X1 port map( A1 => n59810, A2 => n61220, B1 => n3942, B2 => 
                           n15269, ZN => n10242);
   U8696 : OAI22_X1 port map( A1 => n59811, A2 => n61234, B1 => n3941, B2 => 
                           n15269, ZN => n10243);
   U8697 : OAI22_X1 port map( A1 => n59811, A2 => n61257, B1 => n3940, B2 => 
                           n15269, ZN => n10244);
   U8698 : OAI22_X1 port map( A1 => n59764, A2 => n61151, B1 => n52243, B2 => 
                           n59759, ZN => n10077);
   U8699 : OAI22_X1 port map( A1 => n59765, A2 => n61165, B1 => n52242, B2 => 
                           n59759, ZN => n10078);
   U8700 : OAI22_X1 port map( A1 => n59765, A2 => n61179, B1 => n52241, B2 => 
                           n59759, ZN => n10079);
   U8701 : OAI22_X1 port map( A1 => n59765, A2 => n61193, B1 => n52240, B2 => 
                           n59759, ZN => n10080);
   U8702 : OAI22_X1 port map( A1 => n59765, A2 => n61207, B1 => n52239, B2 => 
                           n15285, ZN => n10081);
   U8703 : OAI22_X1 port map( A1 => n59755, A2 => n61151, B1 => n1266, B2 => 
                           n59748, ZN => n10045);
   U8704 : OAI22_X1 port map( A1 => n59755, A2 => n61165, B1 => n1265, B2 => 
                           n59748, ZN => n10046);
   U8705 : OAI22_X1 port map( A1 => n59755, A2 => n61179, B1 => n1264, B2 => 
                           n59748, ZN => n10047);
   U8706 : OAI22_X1 port map( A1 => n59755, A2 => n61193, B1 => n1263, B2 => 
                           n59748, ZN => n10048);
   U8707 : OAI22_X1 port map( A1 => n59756, A2 => n61207, B1 => n1262, B2 => 
                           n15286, ZN => n10049);
   U8708 : OAI22_X1 port map( A1 => n59756, A2 => n61221, B1 => n1261, B2 => 
                           n15286, ZN => n10050);
   U8709 : OAI22_X1 port map( A1 => n59756, A2 => n61235, B1 => n1260, B2 => 
                           n15286, ZN => n10051);
   U8710 : OAI22_X1 port map( A1 => n59756, A2 => n61258, B1 => n1259, B2 => 
                           n15286, ZN => n10052);
   U8711 : OAI22_X1 port map( A1 => n60097, A2 => n61148, B1 => n1258, B2 => 
                           n60092, ZN => n11261);
   U8712 : OAI22_X1 port map( A1 => n60098, A2 => n61162, B1 => n1257, B2 => 
                           n60092, ZN => n11262);
   U8713 : OAI22_X1 port map( A1 => n60098, A2 => n61176, B1 => n1256, B2 => 
                           n60092, ZN => n11263);
   U8714 : OAI22_X1 port map( A1 => n60098, A2 => n61190, B1 => n1255, B2 => 
                           n60092, ZN => n11264);
   U8715 : OAI22_X1 port map( A1 => n60098, A2 => n61204, B1 => n1254, B2 => 
                           n15229, ZN => n11265);
   U8716 : OAI22_X1 port map( A1 => n60098, A2 => n61218, B1 => n1253, B2 => 
                           n15229, ZN => n11266);
   U8717 : OAI22_X1 port map( A1 => n60099, A2 => n61232, B1 => n1252, B2 => 
                           n15229, ZN => n11267);
   U8718 : OAI22_X1 port map( A1 => n60099, A2 => n61255, B1 => n1251, B2 => 
                           n15229, ZN => n11268);
   U8719 : OAI22_X1 port map( A1 => n60070, A2 => n61148, B1 => n1234, B2 => 
                           n60065, ZN => n11165);
   U8720 : OAI22_X1 port map( A1 => n60071, A2 => n61162, B1 => n1233, B2 => 
                           n60065, ZN => n11166);
   U8721 : OAI22_X1 port map( A1 => n60071, A2 => n61176, B1 => n1232, B2 => 
                           n60065, ZN => n11167);
   U8722 : OAI22_X1 port map( A1 => n60071, A2 => n61190, B1 => n1231, B2 => 
                           n60065, ZN => n11168);
   U8723 : OAI22_X1 port map( A1 => n60071, A2 => n61204, B1 => n1230, B2 => 
                           n15233, ZN => n11169);
   U8724 : OAI22_X1 port map( A1 => n60071, A2 => n61218, B1 => n1229, B2 => 
                           n15233, ZN => n11170);
   U8725 : OAI22_X1 port map( A1 => n60072, A2 => n61232, B1 => n1228, B2 => 
                           n15233, ZN => n11171);
   U8726 : OAI22_X1 port map( A1 => n60072, A2 => n61255, B1 => n1227, B2 => 
                           n15233, ZN => n11172);
   U8727 : OAI22_X1 port map( A1 => n60061, A2 => n61148, B1 => n1226, B2 => 
                           n60056, ZN => n11133);
   U8728 : OAI22_X1 port map( A1 => n60062, A2 => n61162, B1 => n1225, B2 => 
                           n60056, ZN => n11134);
   U8729 : OAI22_X1 port map( A1 => n60062, A2 => n61176, B1 => n1224, B2 => 
                           n60056, ZN => n11135);
   U8730 : OAI22_X1 port map( A1 => n60062, A2 => n61190, B1 => n1223, B2 => 
                           n60056, ZN => n11136);
   U8731 : OAI22_X1 port map( A1 => n60062, A2 => n61204, B1 => n1222, B2 => 
                           n15234, ZN => n11137);
   U8732 : OAI22_X1 port map( A1 => n60062, A2 => n61218, B1 => n1221, B2 => 
                           n15234, ZN => n11138);
   U8733 : OAI22_X1 port map( A1 => n60063, A2 => n61232, B1 => n1220, B2 => 
                           n15234, ZN => n11139);
   U8734 : OAI22_X1 port map( A1 => n60063, A2 => n61255, B1 => n1219, B2 => 
                           n15234, ZN => n11140);
   U8735 : OAI22_X1 port map( A1 => n60052, A2 => n61148, B1 => n1218, B2 => 
                           n60047, ZN => n11101);
   U8736 : OAI22_X1 port map( A1 => n60053, A2 => n61162, B1 => n1217, B2 => 
                           n60047, ZN => n11102);
   U8737 : OAI22_X1 port map( A1 => n60053, A2 => n61176, B1 => n1216, B2 => 
                           n60047, ZN => n11103);
   U8738 : OAI22_X1 port map( A1 => n60053, A2 => n61190, B1 => n1215, B2 => 
                           n60047, ZN => n11104);
   U8739 : OAI22_X1 port map( A1 => n60053, A2 => n61204, B1 => n1214, B2 => 
                           n15235, ZN => n11105);
   U8740 : OAI22_X1 port map( A1 => n60053, A2 => n61218, B1 => n1213, B2 => 
                           n15235, ZN => n11106);
   U8741 : OAI22_X1 port map( A1 => n60054, A2 => n61232, B1 => n1212, B2 => 
                           n15235, ZN => n11107);
   U8742 : OAI22_X1 port map( A1 => n60054, A2 => n61255, B1 => n1211, B2 => 
                           n15235, ZN => n11108);
   U8743 : OAI22_X1 port map( A1 => n60043, A2 => n61148, B1 => n1210, B2 => 
                           n60038, ZN => n11069);
   U8744 : OAI22_X1 port map( A1 => n60044, A2 => n61162, B1 => n1209, B2 => 
                           n60038, ZN => n11070);
   U8745 : OAI22_X1 port map( A1 => n60044, A2 => n61176, B1 => n1208, B2 => 
                           n60038, ZN => n11071);
   U8746 : OAI22_X1 port map( A1 => n60044, A2 => n61190, B1 => n1207, B2 => 
                           n60038, ZN => n11072);
   U8747 : OAI22_X1 port map( A1 => n60044, A2 => n61204, B1 => n1206, B2 => 
                           n15236, ZN => n11073);
   U8748 : OAI22_X1 port map( A1 => n60044, A2 => n61218, B1 => n1205, B2 => 
                           n15236, ZN => n11074);
   U8749 : OAI22_X1 port map( A1 => n60045, A2 => n61232, B1 => n1204, B2 => 
                           n15236, ZN => n11075);
   U8750 : OAI22_X1 port map( A1 => n60045, A2 => n61255, B1 => n1203, B2 => 
                           n15236, ZN => n11076);
   U8751 : OAI22_X1 port map( A1 => n60034, A2 => n61148, B1 => n1202, B2 => 
                           n60029, ZN => n11037);
   U8752 : OAI22_X1 port map( A1 => n60035, A2 => n61162, B1 => n1201, B2 => 
                           n60029, ZN => n11038);
   U8753 : OAI22_X1 port map( A1 => n60035, A2 => n61176, B1 => n1200, B2 => 
                           n60029, ZN => n11039);
   U8754 : OAI22_X1 port map( A1 => n60035, A2 => n61190, B1 => n1199, B2 => 
                           n60029, ZN => n11040);
   U8755 : OAI22_X1 port map( A1 => n60035, A2 => n61204, B1 => n1198, B2 => 
                           n15237, ZN => n11041);
   U8756 : OAI22_X1 port map( A1 => n60035, A2 => n61218, B1 => n1197, B2 => 
                           n15237, ZN => n11042);
   U8757 : OAI22_X1 port map( A1 => n60036, A2 => n61232, B1 => n1196, B2 => 
                           n15237, ZN => n11043);
   U8758 : OAI22_X1 port map( A1 => n60036, A2 => n61255, B1 => n1195, B2 => 
                           n15237, ZN => n11044);
   U8759 : OAI22_X1 port map( A1 => n59971, A2 => n61149, B1 => n1146, B2 => 
                           n59966, ZN => n10813);
   U8760 : OAI22_X1 port map( A1 => n59972, A2 => n61163, B1 => n1145, B2 => 
                           n59966, ZN => n10814);
   U8761 : OAI22_X1 port map( A1 => n59972, A2 => n61177, B1 => n1144, B2 => 
                           n59966, ZN => n10815);
   U8762 : OAI22_X1 port map( A1 => n59972, A2 => n61191, B1 => n1143, B2 => 
                           n59966, ZN => n10816);
   U8763 : OAI22_X1 port map( A1 => n59972, A2 => n61205, B1 => n1142, B2 => 
                           n15244, ZN => n10817);
   U8764 : OAI22_X1 port map( A1 => n59972, A2 => n61219, B1 => n1141, B2 => 
                           n15244, ZN => n10818);
   U8765 : OAI22_X1 port map( A1 => n59973, A2 => n61233, B1 => n1140, B2 => 
                           n15244, ZN => n10819);
   U8766 : OAI22_X1 port map( A1 => n59973, A2 => n61256, B1 => n1139, B2 => 
                           n15244, ZN => n10820);
   U8767 : OAI22_X1 port map( A1 => n59962, A2 => n61149, B1 => n1138, B2 => 
                           n59957, ZN => n10781);
   U8768 : OAI22_X1 port map( A1 => n59963, A2 => n61163, B1 => n1137, B2 => 
                           n59957, ZN => n10782);
   U8769 : OAI22_X1 port map( A1 => n59963, A2 => n61177, B1 => n1136, B2 => 
                           n59957, ZN => n10783);
   U8770 : OAI22_X1 port map( A1 => n59963, A2 => n61191, B1 => n1135, B2 => 
                           n59957, ZN => n10784);
   U8771 : OAI22_X1 port map( A1 => n59963, A2 => n61205, B1 => n1134, B2 => 
                           n15245, ZN => n10785);
   U8772 : OAI22_X1 port map( A1 => n59963, A2 => n61219, B1 => n1133, B2 => 
                           n15245, ZN => n10786);
   U8773 : OAI22_X1 port map( A1 => n59964, A2 => n61233, B1 => n1132, B2 => 
                           n15245, ZN => n10787);
   U8774 : OAI22_X1 port map( A1 => n59964, A2 => n61256, B1 => n1131, B2 => 
                           n15245, ZN => n10788);
   U8775 : OAI22_X1 port map( A1 => n59908, A2 => n61149, B1 => n1105, B2 => 
                           n59903, ZN => n10589);
   U8776 : OAI22_X1 port map( A1 => n59909, A2 => n61163, B1 => n1104, B2 => 
                           n59903, ZN => n10590);
   U8777 : OAI22_X1 port map( A1 => n59909, A2 => n61177, B1 => n1103, B2 => 
                           n59903, ZN => n10591);
   U8778 : OAI22_X1 port map( A1 => n59909, A2 => n61191, B1 => n1102, B2 => 
                           n59903, ZN => n10592);
   U8779 : OAI22_X1 port map( A1 => n59909, A2 => n61205, B1 => n1101, B2 => 
                           n15252, ZN => n10593);
   U8780 : OAI22_X1 port map( A1 => n59909, A2 => n61219, B1 => n1100, B2 => 
                           n15252, ZN => n10594);
   U8781 : OAI22_X1 port map( A1 => n59910, A2 => n61233, B1 => n1099, B2 => 
                           n15252, ZN => n10595);
   U8782 : OAI22_X1 port map( A1 => n59910, A2 => n61256, B1 => n1098, B2 => 
                           n15252, ZN => n10596);
   U8783 : OAI22_X1 port map( A1 => n59818, A2 => n61150, B1 => n1053, B2 => 
                           n59813, ZN => n10269);
   U8784 : OAI22_X1 port map( A1 => n59819, A2 => n61164, B1 => n1052, B2 => 
                           n59813, ZN => n10270);
   U8785 : OAI22_X1 port map( A1 => n59819, A2 => n61178, B1 => n1051, B2 => 
                           n59813, ZN => n10271);
   U8786 : OAI22_X1 port map( A1 => n59819, A2 => n61192, B1 => n1050, B2 => 
                           n59813, ZN => n10272);
   U8787 : OAI22_X1 port map( A1 => n59819, A2 => n61206, B1 => n1049, B2 => 
                           n15268, ZN => n10273);
   U8788 : OAI22_X1 port map( A1 => n59819, A2 => n61220, B1 => n1048, B2 => 
                           n15268, ZN => n10274);
   U8789 : OAI22_X1 port map( A1 => n59820, A2 => n61234, B1 => n1047, B2 => 
                           n15268, ZN => n10275);
   U8790 : OAI22_X1 port map( A1 => n59820, A2 => n61257, B1 => n1046, B2 => 
                           n15268, ZN => n10276);
   U8791 : OAI22_X1 port map( A1 => n60664, A2 => n61142, B1 => n1037, B2 => 
                           n60659, ZN => n13277);
   U8792 : OAI22_X1 port map( A1 => n60665, A2 => n61156, B1 => n1036, B2 => 
                           n60659, ZN => n13278);
   U8793 : OAI22_X1 port map( A1 => n60665, A2 => n61170, B1 => n1035, B2 => 
                           n60659, ZN => n13279);
   U8794 : OAI22_X1 port map( A1 => n60665, A2 => n61184, B1 => n1034, B2 => 
                           n60659, ZN => n13280);
   U8795 : OAI22_X1 port map( A1 => n60665, A2 => n61198, B1 => n1033, B2 => 
                           n15148, ZN => n13281);
   U8796 : OAI22_X1 port map( A1 => n60665, A2 => n61212, B1 => n1032, B2 => 
                           n15148, ZN => n13282);
   U8797 : OAI22_X1 port map( A1 => n60666, A2 => n61226, B1 => n1031, B2 => 
                           n15148, ZN => n13283);
   U8798 : OAI22_X1 port map( A1 => n60666, A2 => n61249, B1 => n1030, B2 => 
                           n15148, ZN => n13284);
   U8799 : OAI22_X1 port map( A1 => n60511, A2 => n61144, B1 => n810, B2 => 
                           n60506, ZN => n12733);
   U8800 : OAI22_X1 port map( A1 => n60512, A2 => n61158, B1 => n809, B2 => 
                           n60506, ZN => n12734);
   U8801 : OAI22_X1 port map( A1 => n60512, A2 => n61172, B1 => n808, B2 => 
                           n60506, ZN => n12735);
   U8802 : OAI22_X1 port map( A1 => n60512, A2 => n61186, B1 => n807, B2 => 
                           n60506, ZN => n12736);
   U8803 : OAI22_X1 port map( A1 => n60512, A2 => n61200, B1 => n806, B2 => 
                           n15166, ZN => n12737);
   U8804 : OAI22_X1 port map( A1 => n60512, A2 => n61214, B1 => n805, B2 => 
                           n15166, ZN => n12738);
   U8805 : OAI22_X1 port map( A1 => n60513, A2 => n61228, B1 => n804, B2 => 
                           n15166, ZN => n12739);
   U8806 : OAI22_X1 port map( A1 => n60513, A2 => n61251, B1 => n803, B2 => 
                           n15166, ZN => n12740);
   U8807 : OAI22_X1 port map( A1 => n60475, A2 => n61144, B1 => n546, B2 => 
                           n60470, ZN => n12605);
   U8808 : OAI22_X1 port map( A1 => n60476, A2 => n61158, B1 => n545, B2 => 
                           n60470, ZN => n12606);
   U8809 : OAI22_X1 port map( A1 => n60476, A2 => n61172, B1 => n544, B2 => 
                           n60470, ZN => n12607);
   U8810 : OAI22_X1 port map( A1 => n60476, A2 => n61186, B1 => n543, B2 => 
                           n60470, ZN => n12608);
   U8811 : OAI22_X1 port map( A1 => n60476, A2 => n61200, B1 => n542, B2 => 
                           n15170, ZN => n12609);
   U8812 : OAI22_X1 port map( A1 => n60476, A2 => n61214, B1 => n541, B2 => 
                           n15170, ZN => n12610);
   U8813 : OAI22_X1 port map( A1 => n60477, A2 => n61228, B1 => n540, B2 => 
                           n15170, ZN => n12611);
   U8814 : OAI22_X1 port map( A1 => n60477, A2 => n61251, B1 => n539, B2 => 
                           n15170, ZN => n12612);
   U8815 : OAI22_X1 port map( A1 => n60394, A2 => n61145, B1 => n505, B2 => 
                           n60389, ZN => n12317);
   U8816 : OAI22_X1 port map( A1 => n60395, A2 => n61159, B1 => n504, B2 => 
                           n60389, ZN => n12318);
   U8817 : OAI22_X1 port map( A1 => n60395, A2 => n61173, B1 => n503, B2 => 
                           n60389, ZN => n12319);
   U8818 : OAI22_X1 port map( A1 => n60395, A2 => n61187, B1 => n502, B2 => 
                           n60389, ZN => n12320);
   U8819 : OAI22_X1 port map( A1 => n60395, A2 => n61201, B1 => n501, B2 => 
                           n15186, ZN => n12321);
   U8820 : OAI22_X1 port map( A1 => n60395, A2 => n61215, B1 => n500, B2 => 
                           n15186, ZN => n12322);
   U8821 : OAI22_X1 port map( A1 => n60396, A2 => n61229, B1 => n475, B2 => 
                           n15186, ZN => n12323);
   U8822 : OAI22_X1 port map( A1 => n60396, A2 => n61252, B1 => n474, B2 => 
                           n15186, ZN => n12324);
   U8823 : OAI22_X1 port map( A1 => n60871, A2 => n61140, B1 => n460, B2 => 
                           n60866, ZN => n14013);
   U8824 : OAI22_X1 port map( A1 => n60872, A2 => n61154, B1 => n459, B2 => 
                           n60866, ZN => n14014);
   U8825 : OAI22_X1 port map( A1 => n60872, A2 => n61168, B1 => n458, B2 => 
                           n60866, ZN => n14015);
   U8826 : OAI22_X1 port map( A1 => n60872, A2 => n61182, B1 => n457, B2 => 
                           n60866, ZN => n14016);
   U8827 : OAI22_X1 port map( A1 => n60872, A2 => n61196, B1 => n456, B2 => 
                           n15114, ZN => n14017);
   U8828 : OAI22_X1 port map( A1 => n60872, A2 => n61210, B1 => n455, B2 => 
                           n15114, ZN => n14018);
   U8829 : OAI22_X1 port map( A1 => n60873, A2 => n61224, B1 => n454, B2 => 
                           n15114, ZN => n14019);
   U8830 : OAI22_X1 port map( A1 => n60873, A2 => n61247, B1 => n453, B2 => 
                           n15114, ZN => n14020);
   U8831 : OAI22_X1 port map( A1 => n60862, A2 => n61140, B1 => n412, B2 => 
                           n60857, ZN => n13981);
   U8832 : OAI22_X1 port map( A1 => n60863, A2 => n61154, B1 => n411, B2 => 
                           n60857, ZN => n13982);
   U8833 : OAI22_X1 port map( A1 => n60863, A2 => n61168, B1 => n410, B2 => 
                           n60857, ZN => n13983);
   U8834 : OAI22_X1 port map( A1 => n60863, A2 => n61182, B1 => n409, B2 => 
                           n60857, ZN => n13984);
   U8835 : OAI22_X1 port map( A1 => n60863, A2 => n61196, B1 => n408, B2 => 
                           n15116, ZN => n13985);
   U8836 : OAI22_X1 port map( A1 => n60863, A2 => n61210, B1 => n407, B2 => 
                           n15116, ZN => n13986);
   U8837 : OAI22_X1 port map( A1 => n60864, A2 => n61224, B1 => n406, B2 => 
                           n15116, ZN => n13987);
   U8838 : OAI22_X1 port map( A1 => n60864, A2 => n61247, B1 => n405, B2 => 
                           n15116, ZN => n13988);
   U8839 : OAI22_X1 port map( A1 => n60898, A2 => n61140, B1 => n404, B2 => 
                           n60893, ZN => n14109);
   U8840 : OAI22_X1 port map( A1 => n60899, A2 => n61154, B1 => n403, B2 => 
                           n60893, ZN => n14110);
   U8841 : OAI22_X1 port map( A1 => n60899, A2 => n61168, B1 => n402, B2 => 
                           n60893, ZN => n14111);
   U8842 : OAI22_X1 port map( A1 => n60899, A2 => n61182, B1 => n401, B2 => 
                           n60893, ZN => n14112);
   U8843 : OAI22_X1 port map( A1 => n60899, A2 => n61196, B1 => n400, B2 => 
                           n15108, ZN => n14113);
   U8844 : OAI22_X1 port map( A1 => n60899, A2 => n61210, B1 => n399, B2 => 
                           n15108, ZN => n14114);
   U8845 : OAI22_X1 port map( A1 => n60900, A2 => n61224, B1 => n398, B2 => 
                           n15108, ZN => n14115);
   U8846 : OAI22_X1 port map( A1 => n60900, A2 => n61247, B1 => n397, B2 => 
                           n15108, ZN => n14116);
   U8847 : OAI22_X1 port map( A1 => n60331, A2 => n61145, B1 => n364, B2 => 
                           n60326, ZN => n12093);
   U8848 : OAI22_X1 port map( A1 => n60332, A2 => n61159, B1 => n363, B2 => 
                           n60326, ZN => n12094);
   U8849 : OAI22_X1 port map( A1 => n60332, A2 => n61173, B1 => n362, B2 => 
                           n60326, ZN => n12095);
   U8850 : OAI22_X1 port map( A1 => n60332, A2 => n61187, B1 => n361, B2 => 
                           n60326, ZN => n12096);
   U8851 : OAI22_X1 port map( A1 => n60332, A2 => n61201, B1 => n360, B2 => 
                           n15194, ZN => n12097);
   U8852 : OAI22_X1 port map( A1 => n60332, A2 => n61215, B1 => n359, B2 => 
                           n15194, ZN => n12098);
   U8853 : OAI22_X1 port map( A1 => n60333, A2 => n61229, B1 => n358, B2 => 
                           n15194, ZN => n12099);
   U8854 : OAI22_X1 port map( A1 => n60333, A2 => n61252, B1 => n357, B2 => 
                           n15194, ZN => n12100);
   U8855 : OAI22_X1 port map( A1 => n60322, A2 => n61145, B1 => n356, B2 => 
                           n60317, ZN => n12061);
   U8856 : OAI22_X1 port map( A1 => n60323, A2 => n61159, B1 => n339, B2 => 
                           n60317, ZN => n12062);
   U8857 : OAI22_X1 port map( A1 => n60323, A2 => n61173, B1 => n338, B2 => 
                           n60317, ZN => n12063);
   U8858 : OAI22_X1 port map( A1 => n60323, A2 => n61187, B1 => n337, B2 => 
                           n60317, ZN => n12064);
   U8859 : OAI22_X1 port map( A1 => n60323, A2 => n61201, B1 => n336, B2 => 
                           n15195, ZN => n12065);
   U8860 : OAI22_X1 port map( A1 => n60323, A2 => n61215, B1 => n335, B2 => 
                           n15195, ZN => n12066);
   U8861 : OAI22_X1 port map( A1 => n60324, A2 => n61229, B1 => n334, B2 => 
                           n15195, ZN => n12067);
   U8862 : OAI22_X1 port map( A1 => n60324, A2 => n61252, B1 => n333, B2 => 
                           n15195, ZN => n12068);
   U8863 : OAI22_X1 port map( A1 => n60295, A2 => n61146, B1 => n316, B2 => 
                           n60290, ZN => n11965);
   U8864 : OAI22_X1 port map( A1 => n60296, A2 => n61160, B1 => n315, B2 => 
                           n60290, ZN => n11966);
   U8865 : OAI22_X1 port map( A1 => n60296, A2 => n61174, B1 => n314, B2 => 
                           n60290, ZN => n11967);
   U8866 : OAI22_X1 port map( A1 => n60296, A2 => n61188, B1 => n313, B2 => 
                           n60290, ZN => n11968);
   U8867 : OAI22_X1 port map( A1 => n60296, A2 => n61202, B1 => n312, B2 => 
                           n15198, ZN => n11969);
   U8868 : OAI22_X1 port map( A1 => n60296, A2 => n61216, B1 => n311, B2 => 
                           n15198, ZN => n11970);
   U8869 : OAI22_X1 port map( A1 => n60297, A2 => n61230, B1 => n310, B2 => 
                           n15198, ZN => n11971);
   U8870 : OAI22_X1 port map( A1 => n60297, A2 => n61253, B1 => n309, B2 => 
                           n15198, ZN => n11972);
   U8871 : OAI22_X1 port map( A1 => n60286, A2 => n61146, B1 => n308, B2 => 
                           n60281, ZN => n11933);
   U8872 : OAI22_X1 port map( A1 => n60287, A2 => n61160, B1 => n307, B2 => 
                           n60281, ZN => n11934);
   U8873 : OAI22_X1 port map( A1 => n60287, A2 => n61174, B1 => n306, B2 => 
                           n60281, ZN => n11935);
   U8874 : OAI22_X1 port map( A1 => n60287, A2 => n61188, B1 => n305, B2 => 
                           n60281, ZN => n11936);
   U8875 : OAI22_X1 port map( A1 => n60287, A2 => n61202, B1 => n304, B2 => 
                           n15199, ZN => n11937);
   U8876 : OAI22_X1 port map( A1 => n60287, A2 => n61216, B1 => n303, B2 => 
                           n15199, ZN => n11938);
   U8877 : OAI22_X1 port map( A1 => n60288, A2 => n61230, B1 => n302, B2 => 
                           n15199, ZN => n11939);
   U8878 : OAI22_X1 port map( A1 => n60288, A2 => n61253, B1 => n301, B2 => 
                           n15199, ZN => n11940);
   U8879 : OAI22_X1 port map( A1 => n60250, A2 => n61146, B1 => n292, B2 => 
                           n60245, ZN => n11805);
   U8880 : OAI22_X1 port map( A1 => n60251, A2 => n61160, B1 => n291, B2 => 
                           n60245, ZN => n11806);
   U8881 : OAI22_X1 port map( A1 => n60251, A2 => n61174, B1 => n290, B2 => 
                           n60245, ZN => n11807);
   U8882 : OAI22_X1 port map( A1 => n60251, A2 => n61188, B1 => n289, B2 => 
                           n60245, ZN => n11808);
   U8883 : OAI22_X1 port map( A1 => n60251, A2 => n61202, B1 => n288, B2 => 
                           n15211, ZN => n11809);
   U8884 : OAI22_X1 port map( A1 => n60251, A2 => n61216, B1 => n287, B2 => 
                           n15211, ZN => n11810);
   U8885 : OAI22_X1 port map( A1 => n60252, A2 => n61230, B1 => n286, B2 => 
                           n15211, ZN => n11811);
   U8886 : OAI22_X1 port map( A1 => n60252, A2 => n61253, B1 => n285, B2 => 
                           n15211, ZN => n11812);
   U8887 : OAI22_X1 port map( A1 => n60178, A2 => n61147, B1 => n244, B2 => 
                           n60173, ZN => n11549);
   U8888 : OAI22_X1 port map( A1 => n60179, A2 => n61161, B1 => n243, B2 => 
                           n60173, ZN => n11550);
   U8889 : OAI22_X1 port map( A1 => n60179, A2 => n61175, B1 => n242, B2 => 
                           n60173, ZN => n11551);
   U8890 : OAI22_X1 port map( A1 => n60179, A2 => n61189, B1 => n241, B2 => 
                           n60173, ZN => n11552);
   U8891 : OAI22_X1 port map( A1 => n60179, A2 => n61203, B1 => n240, B2 => 
                           n15220, ZN => n11553);
   U8892 : OAI22_X1 port map( A1 => n60179, A2 => n61217, B1 => n239, B2 => 
                           n15220, ZN => n11554);
   U8893 : OAI22_X1 port map( A1 => n60180, A2 => n61231, B1 => n238, B2 => 
                           n15220, ZN => n11555);
   U8894 : OAI22_X1 port map( A1 => n60180, A2 => n61254, B1 => n237, B2 => 
                           n15220, ZN => n11556);
   U8895 : OAI22_X1 port map( A1 => n60169, A2 => n61147, B1 => n236, B2 => 
                           n60164, ZN => n11517);
   U8896 : OAI22_X1 port map( A1 => n60170, A2 => n61161, B1 => n235, B2 => 
                           n60164, ZN => n11518);
   U8897 : OAI22_X1 port map( A1 => n60170, A2 => n61175, B1 => n234, B2 => 
                           n60164, ZN => n11519);
   U8898 : OAI22_X1 port map( A1 => n60170, A2 => n61189, B1 => n233, B2 => 
                           n60164, ZN => n11520);
   U8899 : OAI22_X1 port map( A1 => n60170, A2 => n61203, B1 => n232, B2 => 
                           n15221, ZN => n11521);
   U8900 : OAI22_X1 port map( A1 => n60170, A2 => n61217, B1 => n231, B2 => 
                           n15221, ZN => n11522);
   U8901 : OAI22_X1 port map( A1 => n60171, A2 => n61231, B1 => n230, B2 => 
                           n15221, ZN => n11523);
   U8902 : OAI22_X1 port map( A1 => n60171, A2 => n61254, B1 => n229, B2 => 
                           n15221, ZN => n11524);
   U8903 : OAI22_X1 port map( A1 => n60142, A2 => n61147, B1 => n228, B2 => 
                           n60137, ZN => n11421);
   U8904 : OAI22_X1 port map( A1 => n60143, A2 => n61161, B1 => n227, B2 => 
                           n60137, ZN => n11422);
   U8905 : OAI22_X1 port map( A1 => n60143, A2 => n61175, B1 => n226, B2 => 
                           n60137, ZN => n11423);
   U8906 : OAI22_X1 port map( A1 => n60143, A2 => n61189, B1 => n225, B2 => 
                           n60137, ZN => n11424);
   U8907 : OAI22_X1 port map( A1 => n60143, A2 => n61203, B1 => n224, B2 => 
                           n15224, ZN => n11425);
   U8908 : OAI22_X1 port map( A1 => n60143, A2 => n61217, B1 => n223, B2 => 
                           n15224, ZN => n11426);
   U8909 : OAI22_X1 port map( A1 => n60144, A2 => n61231, B1 => n222, B2 => 
                           n15224, ZN => n11427);
   U8910 : OAI22_X1 port map( A1 => n60144, A2 => n61254, B1 => n221, B2 => 
                           n15224, ZN => n11428);
   U8911 : OAI22_X1 port map( A1 => n60133, A2 => n61147, B1 => n220, B2 => 
                           n60128, ZN => n11389);
   U8912 : OAI22_X1 port map( A1 => n60134, A2 => n61161, B1 => n219, B2 => 
                           n60128, ZN => n11390);
   U8913 : OAI22_X1 port map( A1 => n60134, A2 => n61175, B1 => n218, B2 => 
                           n60128, ZN => n11391);
   U8914 : OAI22_X1 port map( A1 => n60134, A2 => n61189, B1 => n217, B2 => 
                           n60128, ZN => n11392);
   U8915 : OAI22_X1 port map( A1 => n60134, A2 => n61203, B1 => n216, B2 => 
                           n15225, ZN => n11393);
   U8916 : OAI22_X1 port map( A1 => n60134, A2 => n61217, B1 => n215, B2 => 
                           n15225, ZN => n11394);
   U8917 : OAI22_X1 port map( A1 => n60135, A2 => n61231, B1 => n214, B2 => 
                           n15225, ZN => n11395);
   U8918 : OAI22_X1 port map( A1 => n60135, A2 => n61254, B1 => n213, B2 => 
                           n15225, ZN => n11396);
   U8919 : OAI22_X1 port map( A1 => n60106, A2 => n61147, B1 => n143, B2 => 
                           n60101, ZN => n11293);
   U8920 : OAI22_X1 port map( A1 => n60107, A2 => n61161, B1 => n142, B2 => 
                           n60101, ZN => n11294);
   U8921 : OAI22_X1 port map( A1 => n60107, A2 => n61175, B1 => n141, B2 => 
                           n60101, ZN => n11295);
   U8922 : OAI22_X1 port map( A1 => n60107, A2 => n61189, B1 => n140, B2 => 
                           n60101, ZN => n11296);
   U8923 : OAI22_X1 port map( A1 => n60107, A2 => n61203, B1 => n139, B2 => 
                           n15228, ZN => n11297);
   U8924 : OAI22_X1 port map( A1 => n60107, A2 => n61217, B1 => n138, B2 => 
                           n15228, ZN => n11298);
   U8925 : OAI22_X1 port map( A1 => n60108, A2 => n61231, B1 => n137, B2 => 
                           n15228, ZN => n11299);
   U8926 : OAI22_X1 port map( A1 => n60108, A2 => n61254, B1 => n136, B2 => 
                           n15228, ZN => n11300);
   U8927 : OAI22_X1 port map( A1 => n60817, A2 => n61141, B1 => n135, B2 => 
                           n60812, ZN => n13821);
   U8928 : OAI22_X1 port map( A1 => n60818, A2 => n61155, B1 => n134, B2 => 
                           n60812, ZN => n13822);
   U8929 : OAI22_X1 port map( A1 => n60818, A2 => n61169, B1 => n133, B2 => 
                           n60812, ZN => n13823);
   U8930 : OAI22_X1 port map( A1 => n60818, A2 => n61183, B1 => n132, B2 => 
                           n60812, ZN => n13824);
   U8931 : OAI22_X1 port map( A1 => n60818, A2 => n61197, B1 => n131, B2 => 
                           n15128, ZN => n13825);
   U8932 : OAI22_X1 port map( A1 => n60818, A2 => n61211, B1 => n130, B2 => 
                           n15128, ZN => n13826);
   U8933 : OAI22_X1 port map( A1 => n60819, A2 => n61225, B1 => n129, B2 => 
                           n15128, ZN => n13827);
   U8934 : OAI22_X1 port map( A1 => n60819, A2 => n61248, B1 => n128, B2 => 
                           n15128, ZN => n13828);
   U8935 : OAI22_X1 port map( A1 => n60790, A2 => n61141, B1 => n2924, B2 => 
                           n60785, ZN => n13725);
   U8936 : OAI22_X1 port map( A1 => n60791, A2 => n61155, B1 => n2923, B2 => 
                           n60785, ZN => n13726);
   U8937 : OAI22_X1 port map( A1 => n60791, A2 => n61169, B1 => n2922, B2 => 
                           n60785, ZN => n13727);
   U8938 : OAI22_X1 port map( A1 => n60791, A2 => n61183, B1 => n2921, B2 => 
                           n60785, ZN => n13728);
   U8939 : OAI22_X1 port map( A1 => n60791, A2 => n61197, B1 => n2920, B2 => 
                           n15132, ZN => n13729);
   U8940 : OAI22_X1 port map( A1 => n60791, A2 => n61211, B1 => n2919, B2 => 
                           n15132, ZN => n13730);
   U8941 : OAI22_X1 port map( A1 => n60792, A2 => n61225, B1 => n2918, B2 => 
                           n15132, ZN => n13731);
   U8942 : OAI22_X1 port map( A1 => n60792, A2 => n61248, B1 => n2917, B2 => 
                           n15132, ZN => n13732);
   U8943 : OAI22_X1 port map( A1 => n60781, A2 => n61141, B1 => n2916, B2 => 
                           n60776, ZN => n13693);
   U8944 : OAI22_X1 port map( A1 => n60782, A2 => n61155, B1 => n2915, B2 => 
                           n60776, ZN => n13694);
   U8945 : OAI22_X1 port map( A1 => n60782, A2 => n61169, B1 => n2914, B2 => 
                           n60776, ZN => n13695);
   U8946 : OAI22_X1 port map( A1 => n60782, A2 => n61183, B1 => n2913, B2 => 
                           n60776, ZN => n13696);
   U8947 : OAI22_X1 port map( A1 => n60782, A2 => n61197, B1 => n2912, B2 => 
                           n15133, ZN => n13697);
   U8948 : OAI22_X1 port map( A1 => n60782, A2 => n61211, B1 => n2911, B2 => 
                           n15133, ZN => n13698);
   U8949 : OAI22_X1 port map( A1 => n60783, A2 => n61225, B1 => n2910, B2 => 
                           n15133, ZN => n13699);
   U8950 : OAI22_X1 port map( A1 => n60783, A2 => n61248, B1 => n2909, B2 => 
                           n15133, ZN => n13700);
   U8951 : OAI22_X1 port map( A1 => n60772, A2 => n61141, B1 => n831, B2 => 
                           n60767, ZN => n13661);
   U8952 : OAI22_X1 port map( A1 => n60773, A2 => n61155, B1 => n830, B2 => 
                           n60767, ZN => n13662);
   U8953 : OAI22_X1 port map( A1 => n60773, A2 => n61169, B1 => n829, B2 => 
                           n60767, ZN => n13663);
   U8954 : OAI22_X1 port map( A1 => n60773, A2 => n61183, B1 => n828, B2 => 
                           n60767, ZN => n13664);
   U8955 : OAI22_X1 port map( A1 => n60773, A2 => n61197, B1 => n827, B2 => 
                           n15134, ZN => n13665);
   U8956 : OAI22_X1 port map( A1 => n60773, A2 => n61211, B1 => n826, B2 => 
                           n15134, ZN => n13666);
   U8957 : OAI22_X1 port map( A1 => n60774, A2 => n61225, B1 => n825, B2 => 
                           n15134, ZN => n13667);
   U8958 : OAI22_X1 port map( A1 => n60774, A2 => n61248, B1 => n824, B2 => 
                           n15134, ZN => n13668);
   U8959 : OAI22_X1 port map( A1 => n60763, A2 => n61141, B1 => n823, B2 => 
                           n60758, ZN => n13629);
   U8960 : OAI22_X1 port map( A1 => n60764, A2 => n61155, B1 => n822, B2 => 
                           n60758, ZN => n13630);
   U8961 : OAI22_X1 port map( A1 => n60764, A2 => n61169, B1 => n821, B2 => 
                           n60758, ZN => n13631);
   U8962 : OAI22_X1 port map( A1 => n60764, A2 => n61183, B1 => n820, B2 => 
                           n60758, ZN => n13632);
   U8963 : OAI22_X1 port map( A1 => n60764, A2 => n61197, B1 => n819, B2 => 
                           n15135, ZN => n13633);
   U8964 : OAI22_X1 port map( A1 => n60764, A2 => n61211, B1 => n818, B2 => 
                           n15135, ZN => n13634);
   U8965 : OAI22_X1 port map( A1 => n60765, A2 => n61225, B1 => n817, B2 => 
                           n15135, ZN => n13635);
   U8966 : OAI22_X1 port map( A1 => n60765, A2 => n61248, B1 => n816, B2 => 
                           n15135, ZN => n13636);
   U8967 : OAI22_X1 port map( A1 => n60754, A2 => n61141, B1 => n103, B2 => 
                           n60749, ZN => n13597);
   U8968 : OAI22_X1 port map( A1 => n60755, A2 => n61155, B1 => n102, B2 => 
                           n60749, ZN => n13598);
   U8969 : OAI22_X1 port map( A1 => n60755, A2 => n61169, B1 => n101, B2 => 
                           n60749, ZN => n13599);
   U8970 : OAI22_X1 port map( A1 => n60755, A2 => n61183, B1 => n100, B2 => 
                           n60749, ZN => n13600);
   U8971 : OAI22_X1 port map( A1 => n60755, A2 => n61197, B1 => n79, B2 => 
                           n15136, ZN => n13601);
   U8972 : OAI22_X1 port map( A1 => n60755, A2 => n61211, B1 => n78, B2 => 
                           n15136, ZN => n13602);
   U8973 : OAI22_X1 port map( A1 => n60756, A2 => n61225, B1 => n77, B2 => 
                           n15136, ZN => n13603);
   U8974 : OAI22_X1 port map( A1 => n60756, A2 => n61248, B1 => n76, B2 => 
                           n15136, ZN => n13604);
   U8975 : OAI22_X1 port map( A1 => n60745, A2 => n61142, B1 => n75, B2 => 
                           n60740, ZN => n13565);
   U8976 : OAI22_X1 port map( A1 => n60746, A2 => n61156, B1 => n74, B2 => 
                           n60740, ZN => n13566);
   U8977 : OAI22_X1 port map( A1 => n60746, A2 => n61170, B1 => n73, B2 => 
                           n60740, ZN => n13567);
   U8978 : OAI22_X1 port map( A1 => n60746, A2 => n61184, B1 => n72, B2 => 
                           n60740, ZN => n13568);
   U8979 : OAI22_X1 port map( A1 => n60746, A2 => n61198, B1 => n71, B2 => 
                           n15137, ZN => n13569);
   U8980 : OAI22_X1 port map( A1 => n60746, A2 => n61212, B1 => n70, B2 => 
                           n15137, ZN => n13570);
   U8981 : OAI22_X1 port map( A1 => n60747, A2 => n61226, B1 => n69, B2 => 
                           n15137, ZN => n13571);
   U8982 : OAI22_X1 port map( A1 => n60747, A2 => n61249, B1 => n68, B2 => 
                           n15137, ZN => n13572);
   U8983 : OAI22_X1 port map( A1 => n59765, A2 => n61221, B1 => n3, B2 => 
                           n15285, ZN => n10082);
   U8984 : OAI22_X1 port map( A1 => n59766, A2 => n61235, B1 => n2, B2 => 
                           n15285, ZN => n10083);
   U8985 : OAI22_X1 port map( A1 => n59766, A2 => n61258, B1 => n1, B2 => 
                           n15285, ZN => n10084);
   U8986 : AOI22_X1 port map( A1 => n2327, A2 => n62154, B1 => n2303, B2 => 
                           n62152, ZN => n6746);
   U8987 : AOI22_X1 port map( A1 => n62156, A2 => n5034, B1 => n52864, B2 => 
                           n62178, ZN => n6723);
   U8988 : AOI22_X1 port map( A1 => n2326, A2 => n62154, B1 => n2302, B2 => 
                           n62152, ZN => n6671);
   U8989 : AOI22_X1 port map( A1 => n62156, A2 => n5033, B1 => n52863, B2 => 
                           n62178, ZN => n6648);
   U8990 : AOI22_X1 port map( A1 => n2325, A2 => n62154, B1 => n2301, B2 => 
                           n62152, ZN => n6596);
   U8991 : AOI22_X1 port map( A1 => n62156, A2 => n5032, B1 => n52862, B2 => 
                           n62178, ZN => n6573);
   U8992 : AOI22_X1 port map( A1 => n2324, A2 => n62154, B1 => n2300, B2 => 
                           n62152, ZN => n6521);
   U8993 : AOI22_X1 port map( A1 => n62156, A2 => n5031, B1 => n52861, B2 => 
                           n62178, ZN => n6498);
   U8994 : AOI22_X1 port map( A1 => n2323, A2 => n62154, B1 => n2299, B2 => 
                           n62152, ZN => n6446);
   U8995 : AOI22_X1 port map( A1 => n62156, A2 => n5030, B1 => n52860, B2 => 
                           n62178, ZN => n6423);
   U8996 : AOI22_X1 port map( A1 => n2322, A2 => n62154, B1 => n999, B2 => 
                           n62152, ZN => n6371);
   U8997 : AOI22_X1 port map( A1 => n62156, A2 => n5029, B1 => n52859, B2 => 
                           n62178, ZN => n6348);
   U8998 : AOI22_X1 port map( A1 => n2321, A2 => n62154, B1 => n998, B2 => 
                           n62152, ZN => n6296);
   U8999 : AOI22_X1 port map( A1 => n62156, A2 => n5028, B1 => n52858, B2 => 
                           n62178, ZN => n6273);
   U9000 : AOI22_X1 port map( A1 => n2320, A2 => n62154, B1 => n997, B2 => 
                           n62152, ZN => n6221);
   U9001 : AOI22_X1 port map( A1 => n62156, A2 => n5027, B1 => n52857, B2 => 
                           n62178, ZN => n6198);
   U9002 : AOI22_X1 port map( A1 => n2319, A2 => n62154, B1 => n996, B2 => 
                           n62152, ZN => n6146);
   U9003 : AOI22_X1 port map( A1 => n62156, A2 => n5026, B1 => n52856, B2 => 
                           n62178, ZN => n6123);
   U9004 : AOI22_X1 port map( A1 => n2332, A2 => n62155, B1 => n2308, B2 => 
                           n62153, ZN => n7121);
   U9005 : AOI22_X1 port map( A1 => n62157, A2 => n5039, B1 => n52869, B2 => 
                           n62179, ZN => n7098);
   U9006 : AOI22_X1 port map( A1 => n2331, A2 => n62155, B1 => n2307, B2 => 
                           n62153, ZN => n7046);
   U9007 : AOI22_X1 port map( A1 => n62157, A2 => n5038, B1 => n52868, B2 => 
                           n62179, ZN => n7023);
   U9008 : AOI22_X1 port map( A1 => n2329, A2 => n62154, B1 => n2305, B2 => 
                           n62152, ZN => n6896);
   U9009 : AOI22_X1 port map( A1 => n62156, A2 => n5036, B1 => n52866, B2 => 
                           n62178, ZN => n6873);
   U9010 : AOI22_X1 port map( A1 => n2328, A2 => n62154, B1 => n2304, B2 => 
                           n62152, ZN => n6821);
   U9011 : AOI22_X1 port map( A1 => n62156, A2 => n5035, B1 => n52865, B2 => 
                           n62178, ZN => n6798);
   U9012 : AOI22_X1 port map( A1 => n2334, A2 => n62155, B1 => n2310, B2 => 
                           n62153, ZN => n7271);
   U9013 : AOI22_X1 port map( A1 => n62157, A2 => n5041, B1 => n52871, B2 => 
                           n62179, ZN => n7248);
   U9014 : AOI22_X1 port map( A1 => n2342, A2 => n62155, B1 => n2318, B2 => 
                           n62153, ZN => n7895);
   U9015 : AOI22_X1 port map( A1 => n62157, A2 => n5049, B1 => n52879, B2 => 
                           n62179, ZN => n7854);
   U9016 : AOI22_X1 port map( A1 => n2341, A2 => n62155, B1 => n2317, B2 => 
                           n62153, ZN => n7796);
   U9017 : AOI22_X1 port map( A1 => n62157, A2 => n5048, B1 => n52878, B2 => 
                           n62179, ZN => n7773);
   U9018 : AOI22_X1 port map( A1 => n2340, A2 => n62155, B1 => n2316, B2 => 
                           n62153, ZN => n7721);
   U9019 : AOI22_X1 port map( A1 => n62157, A2 => n5047, B1 => n52877, B2 => 
                           n62179, ZN => n7698);
   U9020 : AOI22_X1 port map( A1 => n2339, A2 => n62155, B1 => n2315, B2 => 
                           n62153, ZN => n7646);
   U9021 : AOI22_X1 port map( A1 => n62157, A2 => n5046, B1 => n52876, B2 => 
                           n62179, ZN => n7623);
   U9022 : AOI22_X1 port map( A1 => n2338, A2 => n62155, B1 => n2314, B2 => 
                           n62153, ZN => n7571);
   U9023 : AOI22_X1 port map( A1 => n62157, A2 => n5045, B1 => n52875, B2 => 
                           n62179, ZN => n7548);
   U9024 : AOI22_X1 port map( A1 => n2337, A2 => n62155, B1 => n2313, B2 => 
                           n62153, ZN => n7496);
   U9025 : AOI22_X1 port map( A1 => n62157, A2 => n5044, B1 => n52874, B2 => 
                           n62179, ZN => n7473);
   U9026 : AOI22_X1 port map( A1 => n2336, A2 => n62155, B1 => n2312, B2 => 
                           n62153, ZN => n7421);
   U9027 : AOI22_X1 port map( A1 => n62157, A2 => n5043, B1 => n52873, B2 => 
                           n62179, ZN => n7398);
   U9028 : AOI22_X1 port map( A1 => n2335, A2 => n62155, B1 => n2311, B2 => 
                           n62153, ZN => n7346);
   U9029 : AOI22_X1 port map( A1 => n62157, A2 => n5042, B1 => n52872, B2 => 
                           n62179, ZN => n7323);
   U9030 : AOI22_X1 port map( A1 => n2333, A2 => n62155, B1 => n2309, B2 => 
                           n62153, ZN => n7196);
   U9031 : AOI22_X1 port map( A1 => n62157, A2 => n5040, B1 => n52870, B2 => 
                           n62179, ZN => n7173);
   U9032 : AOI22_X1 port map( A1 => n2330, A2 => n62154, B1 => n2306, B2 => 
                           n62152, ZN => n6971);
   U9033 : AOI22_X1 port map( A1 => n62156, A2 => n5037, B1 => n52867, B2 => 
                           n62178, ZN => n6948);
   U9034 : AOI22_X1 port map( A1 => n16675, A2 => n61883, B1 => n16521, B2 => 
                           n61880, ZN => n6740);
   U9035 : AOI22_X1 port map( A1 => n15842, A2 => n61895, B1 => n15818, B2 => 
                           n61892, ZN => n6739);
   U9036 : AOI22_X1 port map( A1 => n696, A2 => n62168, B1 => n720, B2 => 
                           n62166, ZN => n6748);
   U9037 : AOI22_X1 port map( A1 => n16709, A2 => n61874, B1 => n16699, B2 => 
                           n61871, ZN => n6747);
   U9038 : AOI22_X1 port map( A1 => n16627, A2 => n61928, B1 => n16603, B2 => 
                           n61925, ZN => n6731);
   U9039 : AOI22_X1 port map( A1 => n15786, A2 => n61916, B1 => n15787, B2 => 
                           n61913, ZN => n6732);
   U9040 : AOI22_X1 port map( A1 => n2895, A2 => n61793, B1 => n2447, B2 => 
                           n61790, ZN => n6722);
   U9041 : AOI22_X1 port map( A1 => n53484, A2 => n61943, B1 => n61940, B2 => 
                           n4560, ZN => n6724);
   U9042 : AOI22_X1 port map( A1 => n54212, A2 => n62134, B1 => n54164, B2 => 
                           n62132, ZN => n6767);
   U9043 : AOI22_X1 port map( A1 => n15784, A2 => n62138, B1 => n15783, B2 => 
                           n62136, ZN => n6768);
   U9044 : AOI22_X1 port map( A1 => n16545, A2 => n61832, B1 => n15785, B2 => 
                           n61829, ZN => n6766);
   U9045 : AOI22_X1 port map( A1 => n54356, A2 => n61853, B1 => n54332, B2 => 
                           n61850, ZN => n6759);
   U9046 : AOI22_X1 port map( A1 => n54486, A2 => n61841, B1 => n54630, B2 => 
                           n61838, ZN => n6760);
   U9047 : AOI22_X1 port map( A1 => n52168, A2 => n61766, B1 => n52192, B2 => 
                           n61763, ZN => n6783);
   U9048 : AOI22_X1 port map( A1 => n15511, A2 => n61754, B1 => n15455, B2 => 
                           n61751, ZN => n6784);
   U9049 : AOI22_X1 port map( A1 => n53924, A2 => n61811, B1 => n53972, B2 => 
                           n61808, ZN => n6774);
   U9050 : AOI22_X1 port map( A1 => n3011, A2 => n61805, B1 => n2987, B2 => 
                           n61802, ZN => n6775);
   U9051 : AOI22_X1 port map( A1 => n16676, A2 => n61883, B1 => n16522, B2 => 
                           n61880, ZN => n6665);
   U9052 : AOI22_X1 port map( A1 => n15843, A2 => n61895, B1 => n15819, B2 => 
                           n61892, ZN => n6664);
   U9053 : AOI22_X1 port map( A1 => n695, A2 => n62168, B1 => n719, B2 => 
                           n62166, ZN => n6673);
   U9054 : AOI22_X1 port map( A1 => n16710, A2 => n61874, B1 => n16700, B2 => 
                           n61871, ZN => n6672);
   U9055 : AOI22_X1 port map( A1 => n16628, A2 => n61928, B1 => n16604, B2 => 
                           n61925, ZN => n6656);
   U9056 : AOI22_X1 port map( A1 => n15791, A2 => n61916, B1 => n15792, B2 => 
                           n61913, ZN => n6657);
   U9057 : AOI22_X1 port map( A1 => n2894, A2 => n61793, B1 => n2446, B2 => 
                           n61790, ZN => n6647);
   U9058 : AOI22_X1 port map( A1 => n53483, A2 => n61943, B1 => n61940, B2 => 
                           n4559, ZN => n6649);
   U9059 : AOI22_X1 port map( A1 => n54211, A2 => n62134, B1 => n54163, B2 => 
                           n62132, ZN => n6692);
   U9060 : AOI22_X1 port map( A1 => n15789, A2 => n62138, B1 => n15788, B2 => 
                           n62136, ZN => n6693);
   U9061 : AOI22_X1 port map( A1 => n16546, A2 => n61832, B1 => n15790, B2 => 
                           n61829, ZN => n6691);
   U9062 : AOI22_X1 port map( A1 => n54355, A2 => n61853, B1 => n54331, B2 => 
                           n61850, ZN => n6684);
   U9063 : AOI22_X1 port map( A1 => n54487, A2 => n61841, B1 => n54631, B2 => 
                           n61838, ZN => n6685);
   U9064 : AOI22_X1 port map( A1 => n52167, A2 => n61766, B1 => n52191, B2 => 
                           n61763, ZN => n6708);
   U9065 : AOI22_X1 port map( A1 => n15512, A2 => n61754, B1 => n15456, B2 => 
                           n61751, ZN => n6709);
   U9066 : AOI22_X1 port map( A1 => n53923, A2 => n61811, B1 => n53971, B2 => 
                           n61808, ZN => n6699);
   U9067 : AOI22_X1 port map( A1 => n3010, A2 => n61805, B1 => n2986, B2 => 
                           n61802, ZN => n6700);
   U9068 : AOI22_X1 port map( A1 => n16677, A2 => n61883, B1 => n16523, B2 => 
                           n61880, ZN => n6590);
   U9069 : AOI22_X1 port map( A1 => n15844, A2 => n61895, B1 => n15820, B2 => 
                           n61892, ZN => n6589);
   U9070 : AOI22_X1 port map( A1 => n694, A2 => n62168, B1 => n718, B2 => 
                           n62166, ZN => n6598);
   U9071 : AOI22_X1 port map( A1 => n16711, A2 => n61874, B1 => n16701, B2 => 
                           n61871, ZN => n6597);
   U9072 : AOI22_X1 port map( A1 => n16629, A2 => n61928, B1 => n16605, B2 => 
                           n61925, ZN => n6581);
   U9073 : AOI22_X1 port map( A1 => n15796, A2 => n61916, B1 => n15797, B2 => 
                           n61913, ZN => n6582);
   U9074 : AOI22_X1 port map( A1 => n2893, A2 => n61793, B1 => n2445, B2 => 
                           n61790, ZN => n6572);
   U9075 : AOI22_X1 port map( A1 => n53482, A2 => n61943, B1 => n61940, B2 => 
                           n4558, ZN => n6574);
   U9076 : AOI22_X1 port map( A1 => n54210, A2 => n62134, B1 => n54162, B2 => 
                           n62132, ZN => n6617);
   U9077 : AOI22_X1 port map( A1 => n15794, A2 => n62138, B1 => n15793, B2 => 
                           n62136, ZN => n6618);
   U9078 : AOI22_X1 port map( A1 => n16547, A2 => n61832, B1 => n15795, B2 => 
                           n61829, ZN => n6616);
   U9079 : AOI22_X1 port map( A1 => n54354, A2 => n61853, B1 => n54330, B2 => 
                           n61850, ZN => n6609);
   U9080 : AOI22_X1 port map( A1 => n54488, A2 => n61841, B1 => n54632, B2 => 
                           n61838, ZN => n6610);
   U9081 : AOI22_X1 port map( A1 => n52166, A2 => n61766, B1 => n52190, B2 => 
                           n61763, ZN => n6633);
   U9082 : AOI22_X1 port map( A1 => n15513, A2 => n61754, B1 => n15457, B2 => 
                           n61751, ZN => n6634);
   U9083 : AOI22_X1 port map( A1 => n53922, A2 => n61811, B1 => n53970, B2 => 
                           n61808, ZN => n6624);
   U9084 : AOI22_X1 port map( A1 => n3009, A2 => n61805, B1 => n2985, B2 => 
                           n61802, ZN => n6625);
   U9085 : AOI22_X1 port map( A1 => n16678, A2 => n61883, B1 => n16524, B2 => 
                           n61880, ZN => n6515);
   U9086 : AOI22_X1 port map( A1 => n15845, A2 => n61895, B1 => n15821, B2 => 
                           n61892, ZN => n6514);
   U9087 : AOI22_X1 port map( A1 => n693, A2 => n62168, B1 => n717, B2 => 
                           n62166, ZN => n6523);
   U9088 : AOI22_X1 port map( A1 => n16712, A2 => n61874, B1 => n16702, B2 => 
                           n61871, ZN => n6522);
   U9089 : AOI22_X1 port map( A1 => n16630, A2 => n61928, B1 => n16606, B2 => 
                           n61925, ZN => n6506);
   U9090 : AOI22_X1 port map( A1 => n15801, A2 => n61916, B1 => n15802, B2 => 
                           n61913, ZN => n6507);
   U9091 : AOI22_X1 port map( A1 => n2892, A2 => n61793, B1 => n2444, B2 => 
                           n61790, ZN => n6497);
   U9092 : AOI22_X1 port map( A1 => n53481, A2 => n61943, B1 => n61940, B2 => 
                           n4557, ZN => n6499);
   U9093 : AOI22_X1 port map( A1 => n54209, A2 => n62134, B1 => n54161, B2 => 
                           n62132, ZN => n6542);
   U9094 : AOI22_X1 port map( A1 => n15799, A2 => n62138, B1 => n15798, B2 => 
                           n62136, ZN => n6543);
   U9095 : AOI22_X1 port map( A1 => n16548, A2 => n61832, B1 => n15800, B2 => 
                           n61829, ZN => n6541);
   U9096 : AOI22_X1 port map( A1 => n54353, A2 => n61853, B1 => n54329, B2 => 
                           n61850, ZN => n6534);
   U9097 : AOI22_X1 port map( A1 => n54489, A2 => n61841, B1 => n54633, B2 => 
                           n61838, ZN => n6535);
   U9098 : AOI22_X1 port map( A1 => n52165, A2 => n61766, B1 => n52189, B2 => 
                           n61763, ZN => n6558);
   U9099 : AOI22_X1 port map( A1 => n15514, A2 => n61754, B1 => n15458, B2 => 
                           n61751, ZN => n6559);
   U9100 : AOI22_X1 port map( A1 => n53921, A2 => n61811, B1 => n53969, B2 => 
                           n61808, ZN => n6549);
   U9101 : AOI22_X1 port map( A1 => n3008, A2 => n61805, B1 => n2984, B2 => 
                           n61802, ZN => n6550);
   U9102 : AOI22_X1 port map( A1 => n16679, A2 => n61883, B1 => n16525, B2 => 
                           n61880, ZN => n6440);
   U9103 : AOI22_X1 port map( A1 => n15846, A2 => n61895, B1 => n15822, B2 => 
                           n61892, ZN => n6439);
   U9104 : AOI22_X1 port map( A1 => n692, A2 => n62168, B1 => n716, B2 => 
                           n62166, ZN => n6448);
   U9105 : AOI22_X1 port map( A1 => n16713, A2 => n61874, B1 => n16703, B2 => 
                           n61871, ZN => n6447);
   U9106 : AOI22_X1 port map( A1 => n16631, A2 => n61928, B1 => n16607, B2 => 
                           n61925, ZN => n6431);
   U9107 : AOI22_X1 port map( A1 => n15854, A2 => n61916, B1 => n15855, B2 => 
                           n61913, ZN => n6432);
   U9108 : AOI22_X1 port map( A1 => n2891, A2 => n61793, B1 => n2443, B2 => 
                           n61790, ZN => n6422);
   U9109 : AOI22_X1 port map( A1 => n53480, A2 => n61943, B1 => n61940, B2 => 
                           n4556, ZN => n6424);
   U9110 : AOI22_X1 port map( A1 => n54208, A2 => n62134, B1 => n54160, B2 => 
                           n62132, ZN => n6467);
   U9111 : AOI22_X1 port map( A1 => n15852, A2 => n62138, B1 => n15851, B2 => 
                           n62136, ZN => n6468);
   U9112 : AOI22_X1 port map( A1 => n16549, A2 => n61832, B1 => n15853, B2 => 
                           n61829, ZN => n6466);
   U9113 : AOI22_X1 port map( A1 => n54352, A2 => n61853, B1 => n54328, B2 => 
                           n61850, ZN => n6459);
   U9114 : AOI22_X1 port map( A1 => n54490, A2 => n61841, B1 => n54634, B2 => 
                           n61838, ZN => n6460);
   U9115 : AOI22_X1 port map( A1 => n52164, A2 => n61766, B1 => n52188, B2 => 
                           n61763, ZN => n6483);
   U9116 : AOI22_X1 port map( A1 => n15515, A2 => n61754, B1 => n15459, B2 => 
                           n61751, ZN => n6484);
   U9117 : AOI22_X1 port map( A1 => n53920, A2 => n61811, B1 => n53968, B2 => 
                           n61808, ZN => n6474);
   U9118 : AOI22_X1 port map( A1 => n3007, A2 => n61805, B1 => n2983, B2 => 
                           n61802, ZN => n6475);
   U9119 : AOI22_X1 port map( A1 => n16680, A2 => n61883, B1 => n16526, B2 => 
                           n61880, ZN => n6365);
   U9120 : AOI22_X1 port map( A1 => n15847, A2 => n61895, B1 => n15823, B2 => 
                           n61892, ZN => n6364);
   U9121 : AOI22_X1 port map( A1 => n691, A2 => n62168, B1 => n715, B2 => 
                           n62166, ZN => n6373);
   U9122 : AOI22_X1 port map( A1 => n16714, A2 => n61874, B1 => n16704, B2 => 
                           n61871, ZN => n6372);
   U9123 : AOI22_X1 port map( A1 => n16632, A2 => n61928, B1 => n16608, B2 => 
                           n61925, ZN => n6356);
   U9124 : AOI22_X1 port map( A1 => n15859, A2 => n61916, B1 => n15860, B2 => 
                           n61913, ZN => n6357);
   U9125 : AOI22_X1 port map( A1 => n2890, A2 => n61793, B1 => n2442, B2 => 
                           n61790, ZN => n6347);
   U9126 : AOI22_X1 port map( A1 => n53479, A2 => n61943, B1 => n61939, B2 => 
                           n4555, ZN => n6349);
   U9127 : AOI22_X1 port map( A1 => n54207, A2 => n62134, B1 => n54159, B2 => 
                           n62132, ZN => n6392);
   U9128 : AOI22_X1 port map( A1 => n15857, A2 => n62138, B1 => n15856, B2 => 
                           n62136, ZN => n6393);
   U9129 : AOI22_X1 port map( A1 => n16550, A2 => n61832, B1 => n15858, B2 => 
                           n61829, ZN => n6391);
   U9130 : AOI22_X1 port map( A1 => n54351, A2 => n61853, B1 => n54327, B2 => 
                           n61850, ZN => n6384);
   U9131 : AOI22_X1 port map( A1 => n54491, A2 => n61841, B1 => n54635, B2 => 
                           n61838, ZN => n6385);
   U9132 : AOI22_X1 port map( A1 => n52163, A2 => n61766, B1 => n52187, B2 => 
                           n61763, ZN => n6408);
   U9133 : AOI22_X1 port map( A1 => n15516, A2 => n61754, B1 => n15460, B2 => 
                           n61751, ZN => n6409);
   U9134 : AOI22_X1 port map( A1 => n53919, A2 => n61811, B1 => n53967, B2 => 
                           n61808, ZN => n6399);
   U9135 : AOI22_X1 port map( A1 => n3006, A2 => n61805, B1 => n2982, B2 => 
                           n61802, ZN => n6400);
   U9136 : AOI22_X1 port map( A1 => n16681, A2 => n61883, B1 => n16527, B2 => 
                           n61880, ZN => n6290);
   U9137 : AOI22_X1 port map( A1 => n15848, A2 => n61895, B1 => n15824, B2 => 
                           n61892, ZN => n6289);
   U9138 : AOI22_X1 port map( A1 => n690, A2 => n62168, B1 => n714, B2 => 
                           n62166, ZN => n6298);
   U9139 : AOI22_X1 port map( A1 => n16715, A2 => n61874, B1 => n16705, B2 => 
                           n61871, ZN => n6297);
   U9140 : AOI22_X1 port map( A1 => n16633, A2 => n61928, B1 => n16609, B2 => 
                           n61925, ZN => n6281);
   U9141 : AOI22_X1 port map( A1 => n15864, A2 => n61916, B1 => n15865, B2 => 
                           n61913, ZN => n6282);
   U9142 : AOI22_X1 port map( A1 => n2889, A2 => n61793, B1 => n2441, B2 => 
                           n61790, ZN => n6272);
   U9143 : AOI22_X1 port map( A1 => n53478, A2 => n61943, B1 => n61939, B2 => 
                           n4554, ZN => n6274);
   U9144 : AOI22_X1 port map( A1 => n54206, A2 => n62134, B1 => n54158, B2 => 
                           n62132, ZN => n6317);
   U9145 : AOI22_X1 port map( A1 => n15862, A2 => n62138, B1 => n15861, B2 => 
                           n62136, ZN => n6318);
   U9146 : AOI22_X1 port map( A1 => n16551, A2 => n61832, B1 => n15863, B2 => 
                           n61829, ZN => n6316);
   U9147 : AOI22_X1 port map( A1 => n54350, A2 => n61853, B1 => n54326, B2 => 
                           n61850, ZN => n6309);
   U9148 : AOI22_X1 port map( A1 => n54492, A2 => n61841, B1 => n54636, B2 => 
                           n61838, ZN => n6310);
   U9149 : AOI22_X1 port map( A1 => n52162, A2 => n61766, B1 => n52186, B2 => 
                           n61763, ZN => n6333);
   U9150 : AOI22_X1 port map( A1 => n15517, A2 => n61754, B1 => n15461, B2 => 
                           n61751, ZN => n6334);
   U9151 : AOI22_X1 port map( A1 => n53918, A2 => n61811, B1 => n53966, B2 => 
                           n61808, ZN => n6324);
   U9152 : AOI22_X1 port map( A1 => n3005, A2 => n61805, B1 => n2981, B2 => 
                           n61802, ZN => n6325);
   U9153 : AOI22_X1 port map( A1 => n16682, A2 => n61883, B1 => n16528, B2 => 
                           n61880, ZN => n6215);
   U9154 : AOI22_X1 port map( A1 => n15849, A2 => n61895, B1 => n15825, B2 => 
                           n61892, ZN => n6214);
   U9155 : AOI22_X1 port map( A1 => n689, A2 => n62168, B1 => n713, B2 => 
                           n62166, ZN => n6223);
   U9156 : AOI22_X1 port map( A1 => n16716, A2 => n61874, B1 => n16706, B2 => 
                           n61871, ZN => n6222);
   U9157 : AOI22_X1 port map( A1 => n16634, A2 => n61928, B1 => n16610, B2 => 
                           n61925, ZN => n6206);
   U9158 : AOI22_X1 port map( A1 => n15869, A2 => n61916, B1 => n15870, B2 => 
                           n61913, ZN => n6207);
   U9159 : AOI22_X1 port map( A1 => n2888, A2 => n61793, B1 => n2440, B2 => 
                           n61790, ZN => n6197);
   U9160 : AOI22_X1 port map( A1 => n53477, A2 => n61943, B1 => n61939, B2 => 
                           n4553, ZN => n6199);
   U9161 : AOI22_X1 port map( A1 => n54205, A2 => n62134, B1 => n54157, B2 => 
                           n62132, ZN => n6242);
   U9162 : AOI22_X1 port map( A1 => n15867, A2 => n62138, B1 => n15866, B2 => 
                           n62136, ZN => n6243);
   U9163 : AOI22_X1 port map( A1 => n16552, A2 => n61832, B1 => n15868, B2 => 
                           n61829, ZN => n6241);
   U9164 : AOI22_X1 port map( A1 => n54349, A2 => n61853, B1 => n54325, B2 => 
                           n61850, ZN => n6234);
   U9165 : AOI22_X1 port map( A1 => n54493, A2 => n61841, B1 => n54637, B2 => 
                           n61838, ZN => n6235);
   U9166 : AOI22_X1 port map( A1 => n52161, A2 => n61766, B1 => n52185, B2 => 
                           n61763, ZN => n6258);
   U9167 : AOI22_X1 port map( A1 => n15518, A2 => n61754, B1 => n15462, B2 => 
                           n61751, ZN => n6259);
   U9168 : AOI22_X1 port map( A1 => n53917, A2 => n61811, B1 => n53965, B2 => 
                           n61808, ZN => n6249);
   U9169 : AOI22_X1 port map( A1 => n3004, A2 => n61805, B1 => n2980, B2 => 
                           n61802, ZN => n6250);
   U9170 : AOI22_X1 port map( A1 => n16683, A2 => n61883, B1 => n16529, B2 => 
                           n61880, ZN => n6140);
   U9171 : AOI22_X1 port map( A1 => n15850, A2 => n61895, B1 => n15826, B2 => 
                           n61892, ZN => n6139);
   U9172 : AOI22_X1 port map( A1 => n688, A2 => n62168, B1 => n712, B2 => 
                           n62166, ZN => n6148);
   U9173 : AOI22_X1 port map( A1 => n16717, A2 => n61874, B1 => n16707, B2 => 
                           n61871, ZN => n6147);
   U9174 : AOI22_X1 port map( A1 => n16635, A2 => n61928, B1 => n16611, B2 => 
                           n61925, ZN => n6131);
   U9175 : AOI22_X1 port map( A1 => n15874, A2 => n61916, B1 => n15875, B2 => 
                           n61913, ZN => n6132);
   U9176 : AOI22_X1 port map( A1 => n2887, A2 => n61793, B1 => n2439, B2 => 
                           n61790, ZN => n6122);
   U9177 : AOI22_X1 port map( A1 => n53476, A2 => n61943, B1 => n61939, B2 => 
                           n4552, ZN => n6124);
   U9178 : AOI22_X1 port map( A1 => n54204, A2 => n62134, B1 => n54156, B2 => 
                           n62132, ZN => n6167);
   U9179 : AOI22_X1 port map( A1 => n15872, A2 => n62138, B1 => n15871, B2 => 
                           n62136, ZN => n6168);
   U9180 : AOI22_X1 port map( A1 => n16553, A2 => n61832, B1 => n15873, B2 => 
                           n61829, ZN => n6166);
   U9181 : AOI22_X1 port map( A1 => n54348, A2 => n61853, B1 => n54324, B2 => 
                           n61850, ZN => n6159);
   U9182 : AOI22_X1 port map( A1 => n54494, A2 => n61841, B1 => n54638, B2 => 
                           n61838, ZN => n6160);
   U9183 : AOI22_X1 port map( A1 => n52160, A2 => n61766, B1 => n52184, B2 => 
                           n61763, ZN => n6183);
   U9184 : AOI22_X1 port map( A1 => n15519, A2 => n61754, B1 => n15463, B2 => 
                           n61751, ZN => n6184);
   U9185 : AOI22_X1 port map( A1 => n53916, A2 => n61811, B1 => n53964, B2 => 
                           n61808, ZN => n6174);
   U9186 : AOI22_X1 port map( A1 => n3003, A2 => n61805, B1 => n2979, B2 => 
                           n61802, ZN => n6175);
   U9187 : AOI22_X1 port map( A1 => n16670, A2 => n61882, B1 => n16516, B2 => 
                           n61879, ZN => n7115);
   U9188 : AOI22_X1 port map( A1 => n15837, A2 => n61894, B1 => n15813, B2 => 
                           n61891, ZN => n7114);
   U9189 : AOI22_X1 port map( A1 => n701, A2 => n62169, B1 => n725, B2 => 
                           n62167, ZN => n7123);
   U9190 : AOI22_X1 port map( A1 => n16302, A2 => n61873, B1 => n16694, B2 => 
                           n61870, ZN => n7122);
   U9191 : AOI22_X1 port map( A1 => n16622, A2 => n61927, B1 => n16598, B2 => 
                           n61924, ZN => n7106);
   U9192 : AOI22_X1 port map( A1 => n15761, A2 => n61915, B1 => n15762, B2 => 
                           n61912, ZN => n7107);
   U9193 : AOI22_X1 port map( A1 => n2900, A2 => n61792, B1 => n2452, B2 => 
                           n61789, ZN => n7097);
   U9194 : AOI22_X1 port map( A1 => n53489, A2 => n61942, B1 => n61940, B2 => 
                           n4565, ZN => n7099);
   U9195 : AOI22_X1 port map( A1 => n54217, A2 => n62135, B1 => n54169, B2 => 
                           n62133, ZN => n7142);
   U9196 : AOI22_X1 port map( A1 => n15759, A2 => n62139, B1 => n15758, B2 => 
                           n62137, ZN => n7143);
   U9197 : AOI22_X1 port map( A1 => n16540, A2 => n61831, B1 => n15760, B2 => 
                           n61828, ZN => n7141);
   U9198 : AOI22_X1 port map( A1 => n54361, A2 => n61852, B1 => n54337, B2 => 
                           n61849, ZN => n7134);
   U9199 : AOI22_X1 port map( A1 => n54481, A2 => n61840, B1 => n54625, B2 => 
                           n61837, ZN => n7135);
   U9200 : AOI22_X1 port map( A1 => n52173, A2 => n61765, B1 => n52197, B2 => 
                           n61762, ZN => n7158);
   U9201 : AOI22_X1 port map( A1 => n15506, A2 => n61753, B1 => n15450, B2 => 
                           n61750, ZN => n7159);
   U9202 : AOI22_X1 port map( A1 => n53929, A2 => n61810, B1 => n53977, B2 => 
                           n61807, ZN => n7149);
   U9203 : AOI22_X1 port map( A1 => n3016, A2 => n61804, B1 => n2992, B2 => 
                           n61801, ZN => n7150);
   U9204 : AOI22_X1 port map( A1 => n16671, A2 => n61882, B1 => n16517, B2 => 
                           n61879, ZN => n7040);
   U9205 : AOI22_X1 port map( A1 => n15838, A2 => n61894, B1 => n15814, B2 => 
                           n61891, ZN => n7039);
   U9206 : AOI22_X1 port map( A1 => n700, A2 => n62169, B1 => n724, B2 => 
                           n62167, ZN => n7048);
   U9207 : AOI22_X1 port map( A1 => n16304, A2 => n61873, B1 => n16695, B2 => 
                           n61870, ZN => n7047);
   U9208 : AOI22_X1 port map( A1 => n16623, A2 => n61927, B1 => n16599, B2 => 
                           n61924, ZN => n7031);
   U9209 : AOI22_X1 port map( A1 => n15766, A2 => n61915, B1 => n15767, B2 => 
                           n61912, ZN => n7032);
   U9210 : AOI22_X1 port map( A1 => n2899, A2 => n61792, B1 => n2451, B2 => 
                           n61789, ZN => n7022);
   U9211 : AOI22_X1 port map( A1 => n53488, A2 => n61942, B1 => n61940, B2 => 
                           n4564, ZN => n7024);
   U9212 : AOI22_X1 port map( A1 => n54216, A2 => n62135, B1 => n54168, B2 => 
                           n62133, ZN => n7067);
   U9213 : AOI22_X1 port map( A1 => n15764, A2 => n62139, B1 => n15763, B2 => 
                           n62137, ZN => n7068);
   U9214 : AOI22_X1 port map( A1 => n16541, A2 => n61831, B1 => n15765, B2 => 
                           n61828, ZN => n7066);
   U9215 : AOI22_X1 port map( A1 => n54360, A2 => n61852, B1 => n54336, B2 => 
                           n61849, ZN => n7059);
   U9216 : AOI22_X1 port map( A1 => n54482, A2 => n61840, B1 => n54626, B2 => 
                           n61837, ZN => n7060);
   U9217 : AOI22_X1 port map( A1 => n52172, A2 => n61765, B1 => n52196, B2 => 
                           n61762, ZN => n7083);
   U9218 : AOI22_X1 port map( A1 => n15507, A2 => n61753, B1 => n15451, B2 => 
                           n61750, ZN => n7084);
   U9219 : AOI22_X1 port map( A1 => n53928, A2 => n61810, B1 => n53976, B2 => 
                           n61807, ZN => n7074);
   U9220 : AOI22_X1 port map( A1 => n3015, A2 => n61804, B1 => n2991, B2 => 
                           n61801, ZN => n7075);
   U9221 : AOI22_X1 port map( A1 => n16673, A2 => n61883, B1 => n16519, B2 => 
                           n61880, ZN => n6890);
   U9222 : AOI22_X1 port map( A1 => n15840, A2 => n61895, B1 => n15816, B2 => 
                           n61892, ZN => n6889);
   U9223 : AOI22_X1 port map( A1 => n698, A2 => n62168, B1 => n722, B2 => 
                           n62166, ZN => n6898);
   U9224 : AOI22_X1 port map( A1 => n16308, A2 => n61874, B1 => n16697, B2 => 
                           n61871, ZN => n6897);
   U9225 : AOI22_X1 port map( A1 => n16625, A2 => n61928, B1 => n16601, B2 => 
                           n61925, ZN => n6881);
   U9226 : AOI22_X1 port map( A1 => n15776, A2 => n61916, B1 => n15777, B2 => 
                           n61913, ZN => n6882);
   U9227 : AOI22_X1 port map( A1 => n2897, A2 => n61793, B1 => n2449, B2 => 
                           n61790, ZN => n6872);
   U9228 : AOI22_X1 port map( A1 => n53486, A2 => n61943, B1 => n61940, B2 => 
                           n4562, ZN => n6874);
   U9229 : AOI22_X1 port map( A1 => n54214, A2 => n62134, B1 => n54166, B2 => 
                           n62132, ZN => n6917);
   U9230 : AOI22_X1 port map( A1 => n15774, A2 => n62138, B1 => n15773, B2 => 
                           n62136, ZN => n6918);
   U9231 : AOI22_X1 port map( A1 => n16543, A2 => n61832, B1 => n15775, B2 => 
                           n61829, ZN => n6916);
   U9232 : AOI22_X1 port map( A1 => n54358, A2 => n61853, B1 => n54334, B2 => 
                           n61850, ZN => n6909);
   U9233 : AOI22_X1 port map( A1 => n54484, A2 => n61841, B1 => n54628, B2 => 
                           n61838, ZN => n6910);
   U9234 : AOI22_X1 port map( A1 => n52170, A2 => n61766, B1 => n52194, B2 => 
                           n61763, ZN => n6933);
   U9235 : AOI22_X1 port map( A1 => n15509, A2 => n61754, B1 => n15453, B2 => 
                           n61751, ZN => n6934);
   U9236 : AOI22_X1 port map( A1 => n53926, A2 => n61811, B1 => n53974, B2 => 
                           n61808, ZN => n6924);
   U9237 : AOI22_X1 port map( A1 => n3013, A2 => n61805, B1 => n2989, B2 => 
                           n61802, ZN => n6925);
   U9238 : AOI22_X1 port map( A1 => n16674, A2 => n61883, B1 => n16520, B2 => 
                           n61880, ZN => n6815);
   U9239 : AOI22_X1 port map( A1 => n15841, A2 => n61895, B1 => n15817, B2 => 
                           n61892, ZN => n6814);
   U9240 : AOI22_X1 port map( A1 => n697, A2 => n62168, B1 => n721, B2 => 
                           n62166, ZN => n6823);
   U9241 : AOI22_X1 port map( A1 => n16708, A2 => n61874, B1 => n16698, B2 => 
                           n61871, ZN => n6822);
   U9242 : AOI22_X1 port map( A1 => n16626, A2 => n61928, B1 => n16602, B2 => 
                           n61925, ZN => n6806);
   U9243 : AOI22_X1 port map( A1 => n15781, A2 => n61916, B1 => n15782, B2 => 
                           n61913, ZN => n6807);
   U9244 : AOI22_X1 port map( A1 => n2896, A2 => n61793, B1 => n2448, B2 => 
                           n61790, ZN => n6797);
   U9245 : AOI22_X1 port map( A1 => n53485, A2 => n61943, B1 => n61940, B2 => 
                           n4561, ZN => n6799);
   U9246 : AOI22_X1 port map( A1 => n54213, A2 => n62134, B1 => n54165, B2 => 
                           n62132, ZN => n6842);
   U9247 : AOI22_X1 port map( A1 => n15779, A2 => n62138, B1 => n15778, B2 => 
                           n62136, ZN => n6843);
   U9248 : AOI22_X1 port map( A1 => n16544, A2 => n61832, B1 => n15780, B2 => 
                           n61829, ZN => n6841);
   U9249 : AOI22_X1 port map( A1 => n54357, A2 => n61853, B1 => n54333, B2 => 
                           n61850, ZN => n6834);
   U9250 : AOI22_X1 port map( A1 => n54485, A2 => n61841, B1 => n54629, B2 => 
                           n61838, ZN => n6835);
   U9251 : AOI22_X1 port map( A1 => n52169, A2 => n61766, B1 => n52193, B2 => 
                           n61763, ZN => n6858);
   U9252 : AOI22_X1 port map( A1 => n15510, A2 => n61754, B1 => n15454, B2 => 
                           n61751, ZN => n6859);
   U9253 : AOI22_X1 port map( A1 => n53925, A2 => n61811, B1 => n53973, B2 => 
                           n61808, ZN => n6849);
   U9254 : AOI22_X1 port map( A1 => n3012, A2 => n61805, B1 => n2988, B2 => 
                           n61802, ZN => n6850);
   U9255 : AOI22_X1 port map( A1 => n839, A2 => n61720, B1 => n847, B2 => 
                           n61722, ZN => n6032);
   U9256 : AOI22_X1 port map( A1 => n15587, A2 => n61706, B1 => n15588, B2 => 
                           n59636, ZN => n6054);
   U9257 : AOI22_X1 port map( A1 => n513, A2 => n61702, B1 => n522, B2 => 
                           n59637, ZN => n6057);
   U9258 : AOI22_X1 port map( A1 => n52374, A2 => n61714, B1 => n52366, B2 => 
                           n59638, ZN => n6042);
   U9259 : AOI22_X1 port map( A1 => n15419, A2 => n61728, B1 => n15411, B2 => 
                           n59639, ZN => n6019);
   U9260 : AOI22_X1 port map( A1 => n863, A2 => n61732, B1 => n855, B2 => 
                           n59640, ZN => n6016);
   U9261 : AOI22_X1 port map( A1 => n15491, A2 => n61674, B1 => n15483, B2 => 
                           n59641, ZN => n6105);
   U9262 : AOI22_X1 port map( A1 => n50971, A2 => n61682, B1 => n50939, B2 => 
                           n59642, ZN => n6087);
   U9263 : AOI22_X1 port map( A1 => n15475, A2 => n61686, B1 => n15467, B2 => 
                           n59643, ZN => n6084);
   U9264 : AOI22_X1 port map( A1 => n16349, A2 => n61694, B1 => n16341, B2 => 
                           n59644, ZN => n6071);
   U9265 : AOI22_X1 port map( A1 => n838, A2 => n61720, B1 => n846, B2 => 
                           n61722, ZN => n5951);
   U9266 : AOI22_X1 port map( A1 => n15589, A2 => n61706, B1 => n15590, B2 => 
                           n59636, ZN => n5966);
   U9267 : AOI22_X1 port map( A1 => n512, A2 => n61702, B1 => n521, B2 => 
                           n59637, ZN => n5967);
   U9268 : AOI22_X1 port map( A1 => n52373, A2 => n61714, B1 => n52365, B2 => 
                           n59638, ZN => n5958);
   U9269 : AOI22_X1 port map( A1 => n15420, A2 => n61728, B1 => n15412, B2 => 
                           n59639, ZN => n5942);
   U9270 : AOI22_X1 port map( A1 => n862, A2 => n61732, B1 => n854, B2 => 
                           n59640, ZN => n5941);
   U9271 : AOI22_X1 port map( A1 => n15492, A2 => n61674, B1 => n15484, B2 => 
                           n59641, ZN => n6001);
   U9272 : AOI22_X1 port map( A1 => n50970, A2 => n61682, B1 => n50938, B2 => 
                           n59642, ZN => n5987);
   U9273 : AOI22_X1 port map( A1 => n15476, A2 => n61686, B1 => n15468, B2 => 
                           n59643, ZN => n5986);
   U9274 : AOI22_X1 port map( A1 => n16350, A2 => n61694, B1 => n16342, B2 => 
                           n59644, ZN => n5977);
   U9275 : AOI22_X1 port map( A1 => n837, A2 => n61720, B1 => n845, B2 => 
                           n61722, ZN => n5876);
   U9276 : AOI22_X1 port map( A1 => n15591, A2 => n61706, B1 => n15592, B2 => 
                           n59636, ZN => n5891);
   U9277 : AOI22_X1 port map( A1 => n511, A2 => n61702, B1 => n520, B2 => 
                           n59637, ZN => n5892);
   U9278 : AOI22_X1 port map( A1 => n52372, A2 => n61714, B1 => n52364, B2 => 
                           n59638, ZN => n5883);
   U9279 : AOI22_X1 port map( A1 => n15421, A2 => n61728, B1 => n15413, B2 => 
                           n59639, ZN => n5867);
   U9280 : AOI22_X1 port map( A1 => n861, A2 => n61732, B1 => n853, B2 => 
                           n59640, ZN => n5866);
   U9281 : AOI22_X1 port map( A1 => n15493, A2 => n61674, B1 => n15485, B2 => 
                           n59641, ZN => n5926);
   U9282 : AOI22_X1 port map( A1 => n50969, A2 => n61682, B1 => n50937, B2 => 
                           n59642, ZN => n5912);
   U9283 : AOI22_X1 port map( A1 => n15477, A2 => n61686, B1 => n15469, B2 => 
                           n59643, ZN => n5911);
   U9284 : AOI22_X1 port map( A1 => n16351, A2 => n61694, B1 => n16343, B2 => 
                           n59644, ZN => n5902);
   U9285 : AOI22_X1 port map( A1 => n836, A2 => n61720, B1 => n844, B2 => 
                           n61722, ZN => n5801);
   U9286 : AOI22_X1 port map( A1 => n15593, A2 => n61706, B1 => n15594, B2 => 
                           n59636, ZN => n5816);
   U9287 : AOI22_X1 port map( A1 => n510, A2 => n61702, B1 => n518, B2 => 
                           n59637, ZN => n5817);
   U9288 : AOI22_X1 port map( A1 => n52371, A2 => n61714, B1 => n52363, B2 => 
                           n59638, ZN => n5808);
   U9289 : AOI22_X1 port map( A1 => n15422, A2 => n61728, B1 => n15414, B2 => 
                           n59639, ZN => n5792);
   U9290 : AOI22_X1 port map( A1 => n860, A2 => n61732, B1 => n852, B2 => 
                           n59640, ZN => n5791);
   U9291 : AOI22_X1 port map( A1 => n15494, A2 => n61674, B1 => n15486, B2 => 
                           n59641, ZN => n5851);
   U9292 : AOI22_X1 port map( A1 => n50968, A2 => n61682, B1 => n50936, B2 => 
                           n59642, ZN => n5837);
   U9293 : AOI22_X1 port map( A1 => n15478, A2 => n61686, B1 => n15470, B2 => 
                           n59643, ZN => n5836);
   U9294 : AOI22_X1 port map( A1 => n16352, A2 => n61694, B1 => n16344, B2 => 
                           n59644, ZN => n5827);
   U9295 : AOI22_X1 port map( A1 => n835, A2 => n61720, B1 => n843, B2 => 
                           n61722, ZN => n5726);
   U9296 : AOI22_X1 port map( A1 => n15595, A2 => n61706, B1 => n15596, B2 => 
                           n59636, ZN => n5741);
   U9297 : AOI22_X1 port map( A1 => n509, A2 => n61702, B1 => n517, B2 => 
                           n59637, ZN => n5742);
   U9298 : AOI22_X1 port map( A1 => n52370, A2 => n61714, B1 => n52362, B2 => 
                           n59638, ZN => n5733);
   U9299 : AOI22_X1 port map( A1 => n15423, A2 => n61728, B1 => n15415, B2 => 
                           n59639, ZN => n5717);
   U9300 : AOI22_X1 port map( A1 => n859, A2 => n61732, B1 => n851, B2 => 
                           n59640, ZN => n5716);
   U9301 : AOI22_X1 port map( A1 => n15495, A2 => n61674, B1 => n15487, B2 => 
                           n59641, ZN => n5776);
   U9302 : AOI22_X1 port map( A1 => n50967, A2 => n61682, B1 => n50935, B2 => 
                           n59642, ZN => n5762);
   U9303 : AOI22_X1 port map( A1 => n15479, A2 => n61686, B1 => n15471, B2 => 
                           n59643, ZN => n5761);
   U9304 : AOI22_X1 port map( A1 => n16353, A2 => n61694, B1 => n16345, B2 => 
                           n59644, ZN => n5752);
   U9305 : AOI22_X1 port map( A1 => n834, A2 => n61720, B1 => n842, B2 => 
                           n61722, ZN => n5651);
   U9306 : AOI22_X1 port map( A1 => n15597, A2 => n61706, B1 => n15598, B2 => 
                           n59636, ZN => n5666);
   U9307 : AOI22_X1 port map( A1 => n508, A2 => n61702, B1 => n516, B2 => 
                           n59637, ZN => n5667);
   U9308 : AOI22_X1 port map( A1 => n52369, A2 => n61714, B1 => n52361, B2 => 
                           n59638, ZN => n5658);
   U9309 : AOI22_X1 port map( A1 => n15424, A2 => n61728, B1 => n15416, B2 => 
                           n59639, ZN => n5642);
   U9310 : AOI22_X1 port map( A1 => n858, A2 => n61732, B1 => n850, B2 => 
                           n59640, ZN => n5641);
   U9311 : AOI22_X1 port map( A1 => n15496, A2 => n61674, B1 => n15488, B2 => 
                           n59641, ZN => n5701);
   U9312 : AOI22_X1 port map( A1 => n50966, A2 => n61682, B1 => n50934, B2 => 
                           n59642, ZN => n5687);
   U9313 : AOI22_X1 port map( A1 => n15480, A2 => n61686, B1 => n15472, B2 => 
                           n59643, ZN => n5686);
   U9314 : AOI22_X1 port map( A1 => n16354, A2 => n61694, B1 => n16346, B2 => 
                           n59644, ZN => n5677);
   U9315 : AOI22_X1 port map( A1 => n833, A2 => n61720, B1 => n841, B2 => 
                           n61722, ZN => n5576);
   U9316 : AOI22_X1 port map( A1 => n15599, A2 => n61706, B1 => n15600, B2 => 
                           n59636, ZN => n5591);
   U9317 : AOI22_X1 port map( A1 => n507, A2 => n61702, B1 => n515, B2 => 
                           n59637, ZN => n5592);
   U9318 : AOI22_X1 port map( A1 => n52368, A2 => n61714, B1 => n52360, B2 => 
                           n59638, ZN => n5583);
   U9319 : AOI22_X1 port map( A1 => n15425, A2 => n61728, B1 => n15417, B2 => 
                           n59639, ZN => n5567);
   U9320 : AOI22_X1 port map( A1 => n857, A2 => n61732, B1 => n849, B2 => 
                           n59640, ZN => n5566);
   U9321 : AOI22_X1 port map( A1 => n15497, A2 => n61674, B1 => n15489, B2 => 
                           n59641, ZN => n5626);
   U9322 : AOI22_X1 port map( A1 => n50965, A2 => n61682, B1 => n50933, B2 => 
                           n59642, ZN => n5612);
   U9323 : AOI22_X1 port map( A1 => n15481, A2 => n61686, B1 => n15473, B2 => 
                           n59643, ZN => n5611);
   U9324 : AOI22_X1 port map( A1 => n16355, A2 => n61694, B1 => n16347, B2 => 
                           n59644, ZN => n5602);
   U9325 : AOI22_X1 port map( A1 => n832, A2 => n61720, B1 => n840, B2 => 
                           n61722, ZN => n5417);
   U9326 : AOI22_X1 port map( A1 => n15611, A2 => n61706, B1 => n15612, B2 => 
                           n59636, ZN => n5455);
   U9327 : AOI22_X1 port map( A1 => n506, A2 => n61702, B1 => n514, B2 => 
                           n59637, ZN => n5458);
   U9328 : AOI22_X1 port map( A1 => n52367, A2 => n61714, B1 => n52359, B2 => 
                           n59638, ZN => n5434);
   U9329 : AOI22_X1 port map( A1 => n15426, A2 => n61728, B1 => n15418, B2 => 
                           n59639, ZN => n5391);
   U9330 : AOI22_X1 port map( A1 => n856, A2 => n61732, B1 => n848, B2 => 
                           n59640, ZN => n5388);
   U9331 : AOI22_X1 port map( A1 => n15498, A2 => n61674, B1 => n15490, B2 => 
                           n59641, ZN => n5538);
   U9332 : AOI22_X1 port map( A1 => n50964, A2 => n61682, B1 => n50932, B2 => 
                           n59642, ZN => n5502);
   U9333 : AOI22_X1 port map( A1 => n15482, A2 => n61686, B1 => n15474, B2 => 
                           n59643, ZN => n5499);
   U9334 : AOI22_X1 port map( A1 => n16356, A2 => n61694, B1 => n16348, B2 => 
                           n59644, ZN => n5473);
   U9335 : AOI22_X1 port map( A1 => n16668, A2 => n61882, B1 => n16514, B2 => 
                           n61879, ZN => n7265);
   U9336 : AOI22_X1 port map( A1 => n15835, A2 => n61894, B1 => n15811, B2 => 
                           n61891, ZN => n7264);
   U9337 : AOI22_X1 port map( A1 => n703, A2 => n62169, B1 => n727, B2 => 
                           n62167, ZN => n7273);
   U9338 : AOI22_X1 port map( A1 => n16298, A2 => n61873, B1 => n16692, B2 => 
                           n61870, ZN => n7272);
   U9339 : AOI22_X1 port map( A1 => n16620, A2 => n61927, B1 => n16596, B2 => 
                           n61924, ZN => n7256);
   U9340 : AOI22_X1 port map( A1 => n15751, A2 => n61915, B1 => n15752, B2 => 
                           n61912, ZN => n7257);
   U9341 : AOI22_X1 port map( A1 => n2902, A2 => n61792, B1 => n2454, B2 => 
                           n61789, ZN => n7247);
   U9342 : AOI22_X1 port map( A1 => n53491, A2 => n61942, B1 => n61940, B2 => 
                           n4567, ZN => n7249);
   U9343 : AOI22_X1 port map( A1 => n54219, A2 => n62135, B1 => n54171, B2 => 
                           n62133, ZN => n7292);
   U9344 : AOI22_X1 port map( A1 => n15749, A2 => n62139, B1 => n15748, B2 => 
                           n62137, ZN => n7293);
   U9345 : AOI22_X1 port map( A1 => n16538, A2 => n61831, B1 => n15750, B2 => 
                           n61828, ZN => n7291);
   U9346 : AOI22_X1 port map( A1 => n54363, A2 => n61852, B1 => n54339, B2 => 
                           n61849, ZN => n7284);
   U9347 : AOI22_X1 port map( A1 => n54479, A2 => n61840, B1 => n54623, B2 => 
                           n61837, ZN => n7285);
   U9348 : AOI22_X1 port map( A1 => n52175, A2 => n61765, B1 => n52199, B2 => 
                           n61762, ZN => n7308);
   U9349 : AOI22_X1 port map( A1 => n15504, A2 => n61753, B1 => n15448, B2 => 
                           n61750, ZN => n7309);
   U9350 : AOI22_X1 port map( A1 => n53931, A2 => n61810, B1 => n53979, B2 => 
                           n61807, ZN => n7299);
   U9351 : AOI22_X1 port map( A1 => n3018, A2 => n61804, B1 => n2994, B2 => 
                           n61801, ZN => n7300);
   U9352 : AOI22_X1 port map( A1 => n16660, A2 => n61882, B1 => n16506, B2 => 
                           n61879, ZN => n7887);
   U9353 : AOI22_X1 port map( A1 => n15827, A2 => n61894, B1 => n15803, B2 => 
                           n61891, ZN => n7884);
   U9354 : AOI22_X1 port map( A1 => n711, A2 => n62169, B1 => n735, B2 => 
                           n62167, ZN => n7898);
   U9355 : AOI22_X1 port map( A1 => n16320, A2 => n61873, B1 => n16684, B2 => 
                           n61870, ZN => n7897);
   U9356 : AOI22_X1 port map( A1 => n16612, A2 => n61927, B1 => n16588, B2 => 
                           n61924, ZN => n7871);
   U9357 : AOI22_X1 port map( A1 => n15879, A2 => n61915, B1 => n15880, B2 => 
                           n61912, ZN => n7874);
   U9358 : AOI22_X1 port map( A1 => n2486, A2 => n61792, B1 => n2462, B2 => 
                           n61789, ZN => n7847);
   U9359 : AOI22_X1 port map( A1 => n53499, A2 => n61942, B1 => n61941, B2 => 
                           n4575, ZN => n7858);
   U9360 : AOI22_X1 port map( A1 => n54227, A2 => n62135, B1 => n54179, B2 => 
                           n62133, ZN => n7921);
   U9361 : AOI22_X1 port map( A1 => n15877, A2 => n62139, B1 => n15876, B2 => 
                           n62137, ZN => n7922);
   U9362 : AOI22_X1 port map( A1 => n16530, A2 => n61831, B1 => n15878, B2 => 
                           n61828, ZN => n7919);
   U9363 : AOI22_X1 port map( A1 => n54371, A2 => n61852, B1 => n54347, B2 => 
                           n61849, ZN => n7909);
   U9364 : AOI22_X1 port map( A1 => n54495, A2 => n61840, B1 => n54639, B2 => 
                           n61837, ZN => n7911);
   U9365 : AOI22_X1 port map( A1 => n52183, A2 => n61765, B1 => n52207, B2 => 
                           n61762, ZN => n7940);
   U9366 : AOI22_X1 port map( A1 => n15464, A2 => n61753, B1 => n15440, B2 => 
                           n61750, ZN => n7941);
   U9367 : AOI22_X1 port map( A1 => n53939, A2 => n61810, B1 => n53987, B2 => 
                           n61807, ZN => n7929);
   U9368 : AOI22_X1 port map( A1 => n3026, A2 => n61804, B1 => n3002, B2 => 
                           n61801, ZN => n7930);
   U9369 : AOI22_X1 port map( A1 => n16661, A2 => n61882, B1 => n16507, B2 => 
                           n61879, ZN => n7790);
   U9370 : AOI22_X1 port map( A1 => n15828, A2 => n61894, B1 => n15804, B2 => 
                           n61891, ZN => n7789);
   U9371 : AOI22_X1 port map( A1 => n710, A2 => n62169, B1 => n734, B2 => 
                           n62167, ZN => n7798);
   U9372 : AOI22_X1 port map( A1 => n16322, A2 => n61873, B1 => n16685, B2 => 
                           n61870, ZN => n7797);
   U9373 : AOI22_X1 port map( A1 => n16613, A2 => n61927, B1 => n16589, B2 => 
                           n61924, ZN => n7781);
   U9374 : AOI22_X1 port map( A1 => n15884, A2 => n61915, B1 => n15885, B2 => 
                           n61912, ZN => n7782);
   U9375 : AOI22_X1 port map( A1 => n2485, A2 => n61792, B1 => n2461, B2 => 
                           n61789, ZN => n7772);
   U9376 : AOI22_X1 port map( A1 => n53498, A2 => n61942, B1 => n61941, B2 => 
                           n4574, ZN => n7774);
   U9377 : AOI22_X1 port map( A1 => n54226, A2 => n62135, B1 => n54178, B2 => 
                           n62133, ZN => n7817);
   U9378 : AOI22_X1 port map( A1 => n15882, A2 => n62139, B1 => n15881, B2 => 
                           n62137, ZN => n7818);
   U9379 : AOI22_X1 port map( A1 => n16531, A2 => n61831, B1 => n15883, B2 => 
                           n61828, ZN => n7816);
   U9380 : AOI22_X1 port map( A1 => n54370, A2 => n61852, B1 => n54346, B2 => 
                           n61849, ZN => n7809);
   U9381 : AOI22_X1 port map( A1 => n54496, A2 => n61840, B1 => n54640, B2 => 
                           n61837, ZN => n7810);
   U9382 : AOI22_X1 port map( A1 => n52182, A2 => n61765, B1 => n52206, B2 => 
                           n61762, ZN => n7833);
   U9383 : AOI22_X1 port map( A1 => n15465, A2 => n61753, B1 => n15441, B2 => 
                           n61750, ZN => n7834);
   U9384 : AOI22_X1 port map( A1 => n53938, A2 => n61810, B1 => n53986, B2 => 
                           n61807, ZN => n7824);
   U9385 : AOI22_X1 port map( A1 => n3025, A2 => n61804, B1 => n3001, B2 => 
                           n61801, ZN => n7825);
   U9386 : AOI22_X1 port map( A1 => n16662, A2 => n61882, B1 => n16508, B2 => 
                           n61879, ZN => n7715);
   U9387 : AOI22_X1 port map( A1 => n15829, A2 => n61894, B1 => n15805, B2 => 
                           n61891, ZN => n7714);
   U9388 : AOI22_X1 port map( A1 => n709, A2 => n62169, B1 => n733, B2 => 
                           n62167, ZN => n7723);
   U9389 : AOI22_X1 port map( A1 => n16324, A2 => n61873, B1 => n16686, B2 => 
                           n61870, ZN => n7722);
   U9390 : AOI22_X1 port map( A1 => n16614, A2 => n61927, B1 => n16590, B2 => 
                           n61924, ZN => n7706);
   U9391 : AOI22_X1 port map( A1 => n15914, A2 => n61915, B1 => n15915, B2 => 
                           n61912, ZN => n7707);
   U9392 : AOI22_X1 port map( A1 => n2484, A2 => n61792, B1 => n2460, B2 => 
                           n61789, ZN => n7697);
   U9393 : AOI22_X1 port map( A1 => n53497, A2 => n61942, B1 => n61941, B2 => 
                           n4573, ZN => n7699);
   U9394 : AOI22_X1 port map( A1 => n54225, A2 => n62135, B1 => n54177, B2 => 
                           n62133, ZN => n7742);
   U9395 : AOI22_X1 port map( A1 => n15887, A2 => n62139, B1 => n15886, B2 => 
                           n62137, ZN => n7743);
   U9396 : AOI22_X1 port map( A1 => n16532, A2 => n61831, B1 => n15888, B2 => 
                           n61828, ZN => n7741);
   U9397 : AOI22_X1 port map( A1 => n54369, A2 => n61852, B1 => n54345, B2 => 
                           n61849, ZN => n7734);
   U9398 : AOI22_X1 port map( A1 => n54497, A2 => n61840, B1 => n54641, B2 => 
                           n61837, ZN => n7735);
   U9399 : AOI22_X1 port map( A1 => n52181, A2 => n61765, B1 => n52205, B2 => 
                           n61762, ZN => n7758);
   U9400 : AOI22_X1 port map( A1 => n15466, A2 => n61753, B1 => n15442, B2 => 
                           n61750, ZN => n7759);
   U9401 : AOI22_X1 port map( A1 => n53937, A2 => n61810, B1 => n53985, B2 => 
                           n61807, ZN => n7749);
   U9402 : AOI22_X1 port map( A1 => n3024, A2 => n61804, B1 => n3000, B2 => 
                           n61801, ZN => n7750);
   U9403 : AOI22_X1 port map( A1 => n16663, A2 => n61882, B1 => n16509, B2 => 
                           n61879, ZN => n7640);
   U9404 : AOI22_X1 port map( A1 => n15830, A2 => n61894, B1 => n15806, B2 => 
                           n61891, ZN => n7639);
   U9405 : AOI22_X1 port map( A1 => n708, A2 => n62169, B1 => n732, B2 => 
                           n62167, ZN => n7648);
   U9406 : AOI22_X1 port map( A1 => n16326, A2 => n61873, B1 => n16687, B2 => 
                           n61870, ZN => n7647);
   U9407 : AOI22_X1 port map( A1 => n16615, A2 => n61927, B1 => n16591, B2 => 
                           n61924, ZN => n7631);
   U9408 : AOI22_X1 port map( A1 => n15892, A2 => n61915, B1 => n15893, B2 => 
                           n61912, ZN => n7632);
   U9409 : AOI22_X1 port map( A1 => n2483, A2 => n61792, B1 => n2459, B2 => 
                           n61789, ZN => n7622);
   U9410 : AOI22_X1 port map( A1 => n53496, A2 => n61942, B1 => n61941, B2 => 
                           n4572, ZN => n7624);
   U9411 : AOI22_X1 port map( A1 => n54224, A2 => n62135, B1 => n54176, B2 => 
                           n62133, ZN => n7667);
   U9412 : AOI22_X1 port map( A1 => n15890, A2 => n62139, B1 => n15889, B2 => 
                           n62137, ZN => n7668);
   U9413 : AOI22_X1 port map( A1 => n16533, A2 => n61831, B1 => n15891, B2 => 
                           n61828, ZN => n7666);
   U9414 : AOI22_X1 port map( A1 => n54368, A2 => n61852, B1 => n54344, B2 => 
                           n61849, ZN => n7659);
   U9415 : AOI22_X1 port map( A1 => n54498, A2 => n61840, B1 => n54642, B2 => 
                           n61837, ZN => n7660);
   U9416 : AOI22_X1 port map( A1 => n52180, A2 => n61765, B1 => n52204, B2 => 
                           n61762, ZN => n7683);
   U9417 : AOI22_X1 port map( A1 => n15499, A2 => n61753, B1 => n15443, B2 => 
                           n61750, ZN => n7684);
   U9418 : AOI22_X1 port map( A1 => n53936, A2 => n61810, B1 => n53984, B2 => 
                           n61807, ZN => n7674);
   U9419 : AOI22_X1 port map( A1 => n3023, A2 => n61804, B1 => n2999, B2 => 
                           n61801, ZN => n7675);
   U9420 : AOI22_X1 port map( A1 => n519, A2 => n61906, B1 => n61905, B2 => 
                           n5021, ZN => n7563);
   U9421 : AOI22_X1 port map( A1 => n16664, A2 => n61882, B1 => n16510, B2 => 
                           n61879, ZN => n7565);
   U9422 : AOI22_X1 port map( A1 => n15831, A2 => n61894, B1 => n15807, B2 => 
                           n61891, ZN => n7564);
   U9423 : AOI22_X1 port map( A1 => n707, A2 => n62169, B1 => n731, B2 => 
                           n62167, ZN => n7573);
   U9424 : AOI22_X1 port map( A1 => n16328, A2 => n61873, B1 => n16688, B2 => 
                           n61870, ZN => n7572);
   U9425 : AOI22_X1 port map( A1 => n16616, A2 => n61927, B1 => n16592, B2 => 
                           n61924, ZN => n7556);
   U9426 : AOI22_X1 port map( A1 => n15897, A2 => n61915, B1 => n15898, B2 => 
                           n61912, ZN => n7557);
   U9427 : AOI22_X1 port map( A1 => n2906, A2 => n61792, B1 => n2458, B2 => 
                           n61789, ZN => n7547);
   U9428 : AOI22_X1 port map( A1 => n53495, A2 => n61942, B1 => n61941, B2 => 
                           n4571, ZN => n7549);
   U9429 : AOI22_X1 port map( A1 => n54223, A2 => n62135, B1 => n54175, B2 => 
                           n62133, ZN => n7592);
   U9430 : AOI22_X1 port map( A1 => n15895, A2 => n62139, B1 => n15894, B2 => 
                           n62137, ZN => n7593);
   U9431 : AOI22_X1 port map( A1 => n16534, A2 => n61831, B1 => n15896, B2 => 
                           n61828, ZN => n7591);
   U9432 : AOI22_X1 port map( A1 => n54367, A2 => n61852, B1 => n54343, B2 => 
                           n61849, ZN => n7584);
   U9433 : AOI22_X1 port map( A1 => n54499, A2 => n61840, B1 => n54643, B2 => 
                           n61837, ZN => n7585);
   U9434 : AOI22_X1 port map( A1 => n52179, A2 => n61765, B1 => n52203, B2 => 
                           n61762, ZN => n7608);
   U9435 : AOI22_X1 port map( A1 => n15500, A2 => n61753, B1 => n15444, B2 => 
                           n61750, ZN => n7609);
   U9436 : AOI22_X1 port map( A1 => n53935, A2 => n61810, B1 => n53983, B2 => 
                           n61807, ZN => n7599);
   U9437 : AOI22_X1 port map( A1 => n3022, A2 => n61804, B1 => n2998, B2 => 
                           n61801, ZN => n7600);
   U9438 : AOI22_X1 port map( A1 => n16665, A2 => n61882, B1 => n16511, B2 => 
                           n61879, ZN => n7490);
   U9439 : AOI22_X1 port map( A1 => n15832, A2 => n61894, B1 => n15808, B2 => 
                           n61891, ZN => n7489);
   U9440 : AOI22_X1 port map( A1 => n706, A2 => n62169, B1 => n730, B2 => 
                           n62167, ZN => n7498);
   U9441 : AOI22_X1 port map( A1 => n16330, A2 => n61873, B1 => n16689, B2 => 
                           n61870, ZN => n7497);
   U9442 : AOI22_X1 port map( A1 => n16617, A2 => n61927, B1 => n16593, B2 => 
                           n61924, ZN => n7481);
   U9443 : AOI22_X1 port map( A1 => n15902, A2 => n61915, B1 => n15903, B2 => 
                           n61912, ZN => n7482);
   U9444 : AOI22_X1 port map( A1 => n2905, A2 => n61792, B1 => n2457, B2 => 
                           n61789, ZN => n7472);
   U9445 : AOI22_X1 port map( A1 => n53494, A2 => n61942, B1 => n61941, B2 => 
                           n4570, ZN => n7474);
   U9446 : AOI22_X1 port map( A1 => n54222, A2 => n62135, B1 => n54174, B2 => 
                           n62133, ZN => n7517);
   U9447 : AOI22_X1 port map( A1 => n15900, A2 => n62139, B1 => n15899, B2 => 
                           n62137, ZN => n7518);
   U9448 : AOI22_X1 port map( A1 => n16535, A2 => n61831, B1 => n15901, B2 => 
                           n61828, ZN => n7516);
   U9449 : AOI22_X1 port map( A1 => n54366, A2 => n61852, B1 => n54342, B2 => 
                           n61849, ZN => n7509);
   U9450 : AOI22_X1 port map( A1 => n54500, A2 => n61840, B1 => n54644, B2 => 
                           n61837, ZN => n7510);
   U9451 : AOI22_X1 port map( A1 => n52178, A2 => n61765, B1 => n52202, B2 => 
                           n61762, ZN => n7533);
   U9452 : AOI22_X1 port map( A1 => n15501, A2 => n61753, B1 => n15445, B2 => 
                           n61750, ZN => n7534);
   U9453 : AOI22_X1 port map( A1 => n53934, A2 => n61810, B1 => n53982, B2 => 
                           n61807, ZN => n7524);
   U9454 : AOI22_X1 port map( A1 => n3021, A2 => n61804, B1 => n2997, B2 => 
                           n61801, ZN => n7525);
   U9455 : AOI22_X1 port map( A1 => n16666, A2 => n61882, B1 => n16512, B2 => 
                           n61879, ZN => n7415);
   U9456 : AOI22_X1 port map( A1 => n15833, A2 => n61894, B1 => n15809, B2 => 
                           n61891, ZN => n7414);
   U9457 : AOI22_X1 port map( A1 => n705, A2 => n62169, B1 => n729, B2 => 
                           n62167, ZN => n7423);
   U9458 : AOI22_X1 port map( A1 => n16332, A2 => n61873, B1 => n16690, B2 => 
                           n61870, ZN => n7422);
   U9459 : AOI22_X1 port map( A1 => n16618, A2 => n61927, B1 => n16594, B2 => 
                           n61924, ZN => n7406);
   U9460 : AOI22_X1 port map( A1 => n15907, A2 => n61915, B1 => n15908, B2 => 
                           n61912, ZN => n7407);
   U9461 : AOI22_X1 port map( A1 => n2904, A2 => n61792, B1 => n2456, B2 => 
                           n61789, ZN => n7397);
   U9462 : AOI22_X1 port map( A1 => n53493, A2 => n61942, B1 => n61941, B2 => 
                           n4569, ZN => n7399);
   U9463 : AOI22_X1 port map( A1 => n54221, A2 => n62135, B1 => n54173, B2 => 
                           n62133, ZN => n7442);
   U9464 : AOI22_X1 port map( A1 => n15905, A2 => n62139, B1 => n15904, B2 => 
                           n62137, ZN => n7443);
   U9465 : AOI22_X1 port map( A1 => n16536, A2 => n61831, B1 => n15906, B2 => 
                           n61828, ZN => n7441);
   U9466 : AOI22_X1 port map( A1 => n54365, A2 => n61852, B1 => n54341, B2 => 
                           n61849, ZN => n7434);
   U9467 : AOI22_X1 port map( A1 => n54501, A2 => n61840, B1 => n54645, B2 => 
                           n61837, ZN => n7435);
   U9468 : AOI22_X1 port map( A1 => n52177, A2 => n61765, B1 => n52201, B2 => 
                           n61762, ZN => n7458);
   U9469 : AOI22_X1 port map( A1 => n15502, A2 => n61753, B1 => n15446, B2 => 
                           n61750, ZN => n7459);
   U9470 : AOI22_X1 port map( A1 => n53933, A2 => n61810, B1 => n53981, B2 => 
                           n61807, ZN => n7449);
   U9471 : AOI22_X1 port map( A1 => n3020, A2 => n61804, B1 => n2996, B2 => 
                           n61801, ZN => n7450);
   U9472 : AOI22_X1 port map( A1 => n16667, A2 => n61882, B1 => n16513, B2 => 
                           n61879, ZN => n7340);
   U9473 : AOI22_X1 port map( A1 => n15834, A2 => n61894, B1 => n15810, B2 => 
                           n61891, ZN => n7339);
   U9474 : AOI22_X1 port map( A1 => n704, A2 => n62169, B1 => n728, B2 => 
                           n62167, ZN => n7348);
   U9475 : AOI22_X1 port map( A1 => n16334, A2 => n61873, B1 => n16691, B2 => 
                           n61870, ZN => n7347);
   U9476 : AOI22_X1 port map( A1 => n16619, A2 => n61927, B1 => n16595, B2 => 
                           n61924, ZN => n7331);
   U9477 : AOI22_X1 port map( A1 => n15912, A2 => n61915, B1 => n15913, B2 => 
                           n61912, ZN => n7332);
   U9478 : AOI22_X1 port map( A1 => n2903, A2 => n61792, B1 => n2455, B2 => 
                           n61789, ZN => n7322);
   U9479 : AOI22_X1 port map( A1 => n53492, A2 => n61942, B1 => n61940, B2 => 
                           n4568, ZN => n7324);
   U9480 : AOI22_X1 port map( A1 => n54220, A2 => n62135, B1 => n54172, B2 => 
                           n62133, ZN => n7367);
   U9481 : AOI22_X1 port map( A1 => n15910, A2 => n62139, B1 => n15909, B2 => 
                           n62137, ZN => n7368);
   U9482 : AOI22_X1 port map( A1 => n16537, A2 => n61831, B1 => n15911, B2 => 
                           n61828, ZN => n7366);
   U9483 : AOI22_X1 port map( A1 => n54364, A2 => n61852, B1 => n54340, B2 => 
                           n61849, ZN => n7359);
   U9484 : AOI22_X1 port map( A1 => n54502, A2 => n61840, B1 => n54646, B2 => 
                           n61837, ZN => n7360);
   U9485 : AOI22_X1 port map( A1 => n52176, A2 => n61765, B1 => n52200, B2 => 
                           n61762, ZN => n7383);
   U9486 : AOI22_X1 port map( A1 => n15503, A2 => n61753, B1 => n15447, B2 => 
                           n61750, ZN => n7384);
   U9487 : AOI22_X1 port map( A1 => n53932, A2 => n61810, B1 => n53980, B2 => 
                           n61807, ZN => n7374);
   U9488 : AOI22_X1 port map( A1 => n3019, A2 => n61804, B1 => n2995, B2 => 
                           n61801, ZN => n7375);
   U9489 : AOI22_X1 port map( A1 => n16669, A2 => n61882, B1 => n16515, B2 => 
                           n61879, ZN => n7190);
   U9490 : AOI22_X1 port map( A1 => n15836, A2 => n61894, B1 => n15812, B2 => 
                           n61891, ZN => n7189);
   U9491 : AOI22_X1 port map( A1 => n702, A2 => n62169, B1 => n726, B2 => 
                           n62167, ZN => n7198);
   U9492 : AOI22_X1 port map( A1 => n16300, A2 => n61873, B1 => n16693, B2 => 
                           n61870, ZN => n7197);
   U9493 : AOI22_X1 port map( A1 => n16621, A2 => n61927, B1 => n16597, B2 => 
                           n61924, ZN => n7181);
   U9494 : AOI22_X1 port map( A1 => n15756, A2 => n61915, B1 => n15757, B2 => 
                           n61912, ZN => n7182);
   U9495 : AOI22_X1 port map( A1 => n2901, A2 => n61792, B1 => n2453, B2 => 
                           n61789, ZN => n7172);
   U9496 : AOI22_X1 port map( A1 => n53490, A2 => n61942, B1 => n61940, B2 => 
                           n4566, ZN => n7174);
   U9497 : AOI22_X1 port map( A1 => n54218, A2 => n62135, B1 => n54170, B2 => 
                           n62133, ZN => n7217);
   U9498 : AOI22_X1 port map( A1 => n15754, A2 => n62139, B1 => n15753, B2 => 
                           n62137, ZN => n7218);
   U9499 : AOI22_X1 port map( A1 => n16539, A2 => n61831, B1 => n15755, B2 => 
                           n61828, ZN => n7216);
   U9500 : AOI22_X1 port map( A1 => n54362, A2 => n61852, B1 => n54338, B2 => 
                           n61849, ZN => n7209);
   U9501 : AOI22_X1 port map( A1 => n54480, A2 => n61840, B1 => n54624, B2 => 
                           n61837, ZN => n7210);
   U9502 : AOI22_X1 port map( A1 => n52174, A2 => n61765, B1 => n52198, B2 => 
                           n61762, ZN => n7233);
   U9503 : AOI22_X1 port map( A1 => n15505, A2 => n61753, B1 => n15449, B2 => 
                           n61750, ZN => n7234);
   U9504 : AOI22_X1 port map( A1 => n53930, A2 => n61810, B1 => n53978, B2 => 
                           n61807, ZN => n7224);
   U9505 : AOI22_X1 port map( A1 => n3017, A2 => n61804, B1 => n2993, B2 => 
                           n61801, ZN => n7225);
   U9506 : AOI22_X1 port map( A1 => n61556, A2 => n16644, B1 => n61554, B2 => 
                           n16490, ZN => n14392);
   U9507 : AOI22_X1 port map( A1 => n61532, A2 => n16668, B1 => n61530, B2 => 
                           n16514, ZN => n14394);
   U9508 : AOI22_X1 port map( A1 => n61607, A2 => n1778, B1 => n61605, B2 => 
                           n1754, ZN => n14384);
   U9509 : AOI22_X1 port map( A1 => n61595, A2 => n15751, B1 => n61593, B2 => 
                           n15752, ZN => n14385);
   U9510 : AOI22_X1 port map( A1 => n61583, A2 => n4347, B1 => n61581, B2 => 
                           n4371, ZN => n14386);
   U9511 : AOI22_X1 port map( A1 => n61493, A2 => n655, B1 => n61491, B2 => 
                           n679, ZN => n14401);
   U9512 : AOI22_X1 port map( A1 => n61481, A2 => n607, B1 => n61479, B2 => 
                           n631, ZN => n14402);
   U9513 : AOI22_X1 port map( A1 => n61658, A2 => n963, B1 => n61656, B2 => 
                           n951, ZN => n14376);
   U9514 : AOI22_X1 port map( A1 => n61634, A2 => n53491, B1 => n61632, B2 => 
                           n4567, ZN => n14378);
   U9515 : AOI22_X1 port map( A1 => n61352, A2 => n3018, B1 => n61350, B2 => 
                           n2994, ZN => n14428);
   U9516 : AOI22_X1 port map( A1 => n61340, A2 => n15685, B1 => n61338, B2 => 
                           n16556, ZN => n14429);
   U9517 : AOI22_X1 port map( A1 => n61328, A2 => n2902, B1 => n61326, B2 => 
                           n2454, ZN => n14430);
   U9518 : AOI22_X1 port map( A1 => n61379, A2 => n16128, B1 => n61377, B2 => 
                           n16129, ZN => n14422);
   U9519 : AOI22_X1 port map( A1 => n61403, A2 => n15750, B1 => n61401, B2 => 
                           n16538, ZN => n14420);
   U9520 : AOI22_X1 port map( A1 => n61391, A2 => n59649, B1 => n61389, B2 => 
                           n59694, ZN => n14421);
   U9521 : AOI22_X1 port map( A1 => n61289, A2 => n2310, B1 => n61287, B2 => 
                           n2334, ZN => n14437);
   U9522 : AOI22_X1 port map( A1 => n61277, A2 => n15504, B1 => n61275, B2 => 
                           n15448, ZN => n14438);
   U9523 : AOI22_X1 port map( A1 => n61454, A2 => n54339, B1 => n61452, B2 => 
                           n54363, ZN => n14412);
   U9524 : AOI22_X1 port map( A1 => n61442, A2 => n54479, B1 => n61440, B2 => 
                           n54623, ZN => n14413);
   U9525 : AOI22_X1 port map( A1 => n61430, A2 => n54243, B1 => n61428, B2 => 
                           n54267, ZN => n14414);
   U9526 : AOI22_X1 port map( A1 => n61556, A2 => n16645, B1 => n61554, B2 => 
                           n16491, ZN => n9901);
   U9527 : AOI22_X1 port map( A1 => n61532, A2 => n16669, B1 => n61530, B2 => 
                           n16515, ZN => n9903);
   U9528 : AOI22_X1 port map( A1 => n61607, A2 => n1777, B1 => n61605, B2 => 
                           n1753, ZN => n9893);
   U9529 : AOI22_X1 port map( A1 => n61595, A2 => n15756, B1 => n61593, B2 => 
                           n15757, ZN => n9894);
   U9530 : AOI22_X1 port map( A1 => n61583, A2 => n4346, B1 => n61581, B2 => 
                           n4370, ZN => n9895);
   U9531 : AOI22_X1 port map( A1 => n61493, A2 => n654, B1 => n61491, B2 => 
                           n678, ZN => n9910);
   U9532 : AOI22_X1 port map( A1 => n61481, A2 => n606, B1 => n61479, B2 => 
                           n630, ZN => n9911);
   U9533 : AOI22_X1 port map( A1 => n61658, A2 => n4713, B1 => n61656, B2 => 
                           n950, ZN => n9885);
   U9534 : AOI22_X1 port map( A1 => n61634, A2 => n53490, B1 => n61632, B2 => 
                           n4566, ZN => n9887);
   U9535 : AOI22_X1 port map( A1 => n61352, A2 => n3017, B1 => n61350, B2 => 
                           n2993, ZN => n14353);
   U9536 : AOI22_X1 port map( A1 => n61340, A2 => n15688, B1 => n61338, B2 => 
                           n16557, ZN => n14354);
   U9537 : AOI22_X1 port map( A1 => n61328, A2 => n2901, B1 => n61326, B2 => 
                           n2453, ZN => n14355);
   U9538 : AOI22_X1 port map( A1 => n61379, A2 => n16132, B1 => n61377, B2 => 
                           n16133, ZN => n14347);
   U9539 : AOI22_X1 port map( A1 => n61403, A2 => n15755, B1 => n61401, B2 => 
                           n16539, ZN => n14345);
   U9540 : AOI22_X1 port map( A1 => n61391, A2 => n59650, B1 => n61389, B2 => 
                           n59695, ZN => n14346);
   U9541 : AOI22_X1 port map( A1 => n61289, A2 => n2309, B1 => n61287, B2 => 
                           n2333, ZN => n14362);
   U9542 : AOI22_X1 port map( A1 => n61277, A2 => n15505, B1 => n61275, B2 => 
                           n15449, ZN => n14363);
   U9543 : AOI22_X1 port map( A1 => n61454, A2 => n54338, B1 => n61452, B2 => 
                           n54362, ZN => n9921);
   U9544 : AOI22_X1 port map( A1 => n61442, A2 => n54480, B1 => n61440, B2 => 
                           n54624, ZN => n9922);
   U9545 : AOI22_X1 port map( A1 => n61430, A2 => n54242, B1 => n61428, B2 => 
                           n54266, ZN => n9923);
   U9546 : AOI22_X1 port map( A1 => n61556, A2 => n16646, B1 => n61554, B2 => 
                           n16492, ZN => n9826);
   U9547 : AOI22_X1 port map( A1 => n61532, A2 => n16670, B1 => n61530, B2 => 
                           n16516, ZN => n9828);
   U9548 : AOI22_X1 port map( A1 => n61607, A2 => n1776, B1 => n61605, B2 => 
                           n1752, ZN => n9818);
   U9549 : AOI22_X1 port map( A1 => n61595, A2 => n15761, B1 => n61593, B2 => 
                           n15762, ZN => n9819);
   U9550 : AOI22_X1 port map( A1 => n61583, A2 => n4345, B1 => n61581, B2 => 
                           n4369, ZN => n9820);
   U9551 : AOI22_X1 port map( A1 => n61493, A2 => n653, B1 => n61491, B2 => 
                           n677, ZN => n9835);
   U9552 : AOI22_X1 port map( A1 => n61481, A2 => n605, B1 => n61479, B2 => 
                           n629, ZN => n9836);
   U9553 : AOI22_X1 port map( A1 => n61658, A2 => n4712, B1 => n61656, B2 => 
                           n949, ZN => n9746);
   U9554 : AOI22_X1 port map( A1 => n61634, A2 => n53489, B1 => n61632, B2 => 
                           n4565, ZN => n9812);
   U9555 : AOI22_X1 port map( A1 => n61352, A2 => n3016, B1 => n61350, B2 => 
                           n2992, ZN => n9862);
   U9556 : AOI22_X1 port map( A1 => n61340, A2 => n15691, B1 => n61338, B2 => 
                           n16558, ZN => n9863);
   U9557 : AOI22_X1 port map( A1 => n61328, A2 => n2900, B1 => n61326, B2 => 
                           n2452, ZN => n9864);
   U9558 : AOI22_X1 port map( A1 => n61379, A2 => n16134, B1 => n61377, B2 => 
                           n16135, ZN => n9856);
   U9559 : AOI22_X1 port map( A1 => n61403, A2 => n15760, B1 => n61401, B2 => 
                           n16540, ZN => n9854);
   U9560 : AOI22_X1 port map( A1 => n61391, A2 => n59651, B1 => n61389, B2 => 
                           n59696, ZN => n9855);
   U9561 : AOI22_X1 port map( A1 => n61289, A2 => n2308, B1 => n61287, B2 => 
                           n2332, ZN => n9871);
   U9562 : AOI22_X1 port map( A1 => n61277, A2 => n15506, B1 => n61275, B2 => 
                           n15450, ZN => n9872);
   U9563 : AOI22_X1 port map( A1 => n61454, A2 => n54337, B1 => n61452, B2 => 
                           n54361, ZN => n9846);
   U9564 : AOI22_X1 port map( A1 => n61442, A2 => n54481, B1 => n61440, B2 => 
                           n54625, ZN => n9847);
   U9565 : AOI22_X1 port map( A1 => n61430, A2 => n54241, B1 => n61428, B2 => 
                           n54265, ZN => n9848);
   U9566 : AOI22_X1 port map( A1 => n61556, A2 => n16647, B1 => n61554, B2 => 
                           n16493, ZN => n9687);
   U9567 : AOI22_X1 port map( A1 => n61532, A2 => n16671, B1 => n61530, B2 => 
                           n16517, ZN => n9689);
   U9568 : AOI22_X1 port map( A1 => n61607, A2 => n1775, B1 => n61605, B2 => 
                           n1751, ZN => n9679);
   U9569 : AOI22_X1 port map( A1 => n61595, A2 => n15766, B1 => n61593, B2 => 
                           n15767, ZN => n9680);
   U9570 : AOI22_X1 port map( A1 => n61583, A2 => n4344, B1 => n61581, B2 => 
                           n4368, ZN => n9681);
   U9571 : AOI22_X1 port map( A1 => n61493, A2 => n652, B1 => n61491, B2 => 
                           n676, ZN => n9696);
   U9572 : AOI22_X1 port map( A1 => n61481, A2 => n604, B1 => n61479, B2 => 
                           n628, ZN => n9697);
   U9573 : AOI22_X1 port map( A1 => n61658, A2 => n4711, B1 => n61656, B2 => 
                           n948, ZN => n9671);
   U9574 : AOI22_X1 port map( A1 => n61634, A2 => n53488, B1 => n61632, B2 => 
                           n4564, ZN => n9673);
   U9575 : AOI22_X1 port map( A1 => n61352, A2 => n3015, B1 => n61350, B2 => 
                           n2991, ZN => n9723);
   U9576 : AOI22_X1 port map( A1 => n61340, A2 => n15694, B1 => n61338, B2 => 
                           n16559, ZN => n9724);
   U9577 : AOI22_X1 port map( A1 => n61328, A2 => n2899, B1 => n61326, B2 => 
                           n2451, ZN => n9725);
   U9578 : AOI22_X1 port map( A1 => n61379, A2 => n16136, B1 => n61377, B2 => 
                           n16137, ZN => n9717);
   U9579 : AOI22_X1 port map( A1 => n61403, A2 => n15765, B1 => n61401, B2 => 
                           n16541, ZN => n9715);
   U9580 : AOI22_X1 port map( A1 => n61391, A2 => n59652, B1 => n61389, B2 => 
                           n59697, ZN => n9716);
   U9581 : AOI22_X1 port map( A1 => n61289, A2 => n2307, B1 => n61287, B2 => 
                           n2331, ZN => n9732);
   U9582 : AOI22_X1 port map( A1 => n61277, A2 => n15507, B1 => n61275, B2 => 
                           n15451, ZN => n9733);
   U9583 : AOI22_X1 port map( A1 => n61454, A2 => n54336, B1 => n61452, B2 => 
                           n54360, ZN => n9707);
   U9584 : AOI22_X1 port map( A1 => n61442, A2 => n54482, B1 => n61440, B2 => 
                           n54626, ZN => n9708);
   U9585 : AOI22_X1 port map( A1 => n61430, A2 => n54240, B1 => n61428, B2 => 
                           n54264, ZN => n9709);
   U9586 : AOI22_X1 port map( A1 => n61557, A2 => n16648, B1 => n61554, B2 => 
                           n16494, ZN => n9596);
   U9587 : AOI22_X1 port map( A1 => n61533, A2 => n16672, B1 => n61530, B2 => 
                           n16518, ZN => n9598);
   U9588 : AOI22_X1 port map( A1 => n61608, A2 => n1774, B1 => n61605, B2 => 
                           n1750, ZN => n9588);
   U9589 : AOI22_X1 port map( A1 => n61596, A2 => n15771, B1 => n61593, B2 => 
                           n15772, ZN => n9589);
   U9590 : AOI22_X1 port map( A1 => n61584, A2 => n4343, B1 => n61581, B2 => 
                           n4367, ZN => n9590);
   U9591 : AOI22_X1 port map( A1 => n61494, A2 => n651, B1 => n61491, B2 => 
                           n675, ZN => n9621);
   U9592 : AOI22_X1 port map( A1 => n61482, A2 => n603, B1 => n61479, B2 => 
                           n627, ZN => n9622);
   U9593 : AOI22_X1 port map( A1 => n61659, A2 => n4710, B1 => n61656, B2 => 
                           n947, ZN => n9580);
   U9594 : AOI22_X1 port map( A1 => n61635, A2 => n53487, B1 => n61632, B2 => 
                           n4563, ZN => n9582);
   U9595 : AOI22_X1 port map( A1 => n61353, A2 => n3014, B1 => n61350, B2 => 
                           n2990, ZN => n9648);
   U9596 : AOI22_X1 port map( A1 => n61341, A2 => n15386, B1 => n61338, B2 => 
                           n15432, ZN => n9649);
   U9597 : AOI22_X1 port map( A1 => n61329, A2 => n2898, B1 => n61326, B2 => 
                           n2450, ZN => n9650);
   U9598 : AOI22_X1 port map( A1 => n61380, A2 => n16108, B1 => n61377, B2 => 
                           n16109, ZN => n9642);
   U9599 : AOI22_X1 port map( A1 => n61404, A2 => n15770, B1 => n61401, B2 => 
                           n16542, ZN => n9640);
   U9600 : AOI22_X1 port map( A1 => n61392, A2 => n59653, B1 => n61389, B2 => 
                           n59698, ZN => n9641);
   U9601 : AOI22_X1 port map( A1 => n61290, A2 => n2306, B1 => n61287, B2 => 
                           n2330, ZN => n9657);
   U9602 : AOI22_X1 port map( A1 => n61278, A2 => n15508, B1 => n61275, B2 => 
                           n15452, ZN => n9658);
   U9603 : AOI22_X1 port map( A1 => n61455, A2 => n54335, B1 => n61452, B2 => 
                           n54359, ZN => n9632);
   U9604 : AOI22_X1 port map( A1 => n61443, A2 => n54483, B1 => n61440, B2 => 
                           n54627, ZN => n9633);
   U9605 : AOI22_X1 port map( A1 => n61431, A2 => n54239, B1 => n61428, B2 => 
                           n54263, ZN => n9634);
   U9606 : AOI22_X1 port map( A1 => n61557, A2 => n16649, B1 => n61554, B2 => 
                           n16495, ZN => n9521);
   U9607 : AOI22_X1 port map( A1 => n61533, A2 => n16673, B1 => n61530, B2 => 
                           n16519, ZN => n9523);
   U9608 : AOI22_X1 port map( A1 => n61608, A2 => n1773, B1 => n61605, B2 => 
                           n1749, ZN => n9513);
   U9609 : AOI22_X1 port map( A1 => n61596, A2 => n15776, B1 => n61593, B2 => 
                           n15777, ZN => n9514);
   U9610 : AOI22_X1 port map( A1 => n61584, A2 => n4342, B1 => n61581, B2 => 
                           n4366, ZN => n9515);
   U9611 : AOI22_X1 port map( A1 => n61494, A2 => n650, B1 => n61491, B2 => 
                           n674, ZN => n9530);
   U9612 : AOI22_X1 port map( A1 => n61482, A2 => n602, B1 => n61479, B2 => 
                           n626, ZN => n9531);
   U9613 : AOI22_X1 port map( A1 => n61659, A2 => n4709, B1 => n61656, B2 => 
                           n946, ZN => n9505);
   U9614 : AOI22_X1 port map( A1 => n61635, A2 => n53486, B1 => n61632, B2 => 
                           n4562, ZN => n9507);
   U9615 : AOI22_X1 port map( A1 => n61353, A2 => n3013, B1 => n61350, B2 => 
                           n2989, ZN => n9557);
   U9616 : AOI22_X1 port map( A1 => n61341, A2 => n15395, B1 => n61338, B2 => 
                           n15433, ZN => n9558);
   U9617 : AOI22_X1 port map( A1 => n61329, A2 => n2897, B1 => n61326, B2 => 
                           n2449, ZN => n9559);
   U9618 : AOI22_X1 port map( A1 => n61380, A2 => n16120, B1 => n61377, B2 => 
                           n16121, ZN => n9551);
   U9619 : AOI22_X1 port map( A1 => n61404, A2 => n15775, B1 => n61401, B2 => 
                           n16543, ZN => n9549);
   U9620 : AOI22_X1 port map( A1 => n61392, A2 => n59654, B1 => n61389, B2 => 
                           n59699, ZN => n9550);
   U9621 : AOI22_X1 port map( A1 => n61290, A2 => n2305, B1 => n61287, B2 => 
                           n2329, ZN => n9566);
   U9622 : AOI22_X1 port map( A1 => n61278, A2 => n15509, B1 => n61275, B2 => 
                           n15453, ZN => n9567);
   U9623 : AOI22_X1 port map( A1 => n61455, A2 => n54334, B1 => n61452, B2 => 
                           n54358, ZN => n9541);
   U9624 : AOI22_X1 port map( A1 => n61443, A2 => n54484, B1 => n61440, B2 => 
                           n54628, ZN => n9542);
   U9625 : AOI22_X1 port map( A1 => n61431, A2 => n54238, B1 => n61428, B2 => 
                           n54262, ZN => n9543);
   U9626 : AOI22_X1 port map( A1 => n61557, A2 => n16650, B1 => n61554, B2 => 
                           n16496, ZN => n9446);
   U9627 : AOI22_X1 port map( A1 => n61533, A2 => n16674, B1 => n61530, B2 => 
                           n16520, ZN => n9448);
   U9628 : AOI22_X1 port map( A1 => n61608, A2 => n1772, B1 => n61605, B2 => 
                           n1748, ZN => n9438);
   U9629 : AOI22_X1 port map( A1 => n61596, A2 => n15781, B1 => n61593, B2 => 
                           n15782, ZN => n9439);
   U9630 : AOI22_X1 port map( A1 => n61584, A2 => n4341, B1 => n61581, B2 => 
                           n4365, ZN => n9440);
   U9631 : AOI22_X1 port map( A1 => n61494, A2 => n649, B1 => n61491, B2 => 
                           n673, ZN => n9455);
   U9632 : AOI22_X1 port map( A1 => n61482, A2 => n601, B1 => n61479, B2 => 
                           n625, ZN => n9456);
   U9633 : AOI22_X1 port map( A1 => n61659, A2 => n4708, B1 => n61656, B2 => 
                           n945, ZN => n9430);
   U9634 : AOI22_X1 port map( A1 => n61635, A2 => n53485, B1 => n61632, B2 => 
                           n4561, ZN => n9432);
   U9635 : AOI22_X1 port map( A1 => n61353, A2 => n3012, B1 => n61350, B2 => 
                           n2988, ZN => n9482);
   U9636 : AOI22_X1 port map( A1 => n61341, A2 => n15396, B1 => n61338, B2 => 
                           n15434, ZN => n9483);
   U9637 : AOI22_X1 port map( A1 => n61329, A2 => n2896, B1 => n61326, B2 => 
                           n2448, ZN => n9484);
   U9638 : AOI22_X1 port map( A1 => n61380, A2 => n16122, B1 => n61377, B2 => 
                           n16123, ZN => n9476);
   U9639 : AOI22_X1 port map( A1 => n61404, A2 => n15780, B1 => n61401, B2 => 
                           n16544, ZN => n9474);
   U9640 : AOI22_X1 port map( A1 => n61392, A2 => n59655, B1 => n61389, B2 => 
                           n59700, ZN => n9475);
   U9641 : AOI22_X1 port map( A1 => n61290, A2 => n2304, B1 => n61287, B2 => 
                           n2328, ZN => n9491);
   U9642 : AOI22_X1 port map( A1 => n61278, A2 => n15510, B1 => n61275, B2 => 
                           n15454, ZN => n9492);
   U9643 : AOI22_X1 port map( A1 => n61455, A2 => n54333, B1 => n61452, B2 => 
                           n54357, ZN => n9466);
   U9644 : AOI22_X1 port map( A1 => n61443, A2 => n54485, B1 => n61440, B2 => 
                           n54629, ZN => n9467);
   U9645 : AOI22_X1 port map( A1 => n61431, A2 => n54237, B1 => n61428, B2 => 
                           n54261, ZN => n9468);
   U9646 : AOI22_X1 port map( A1 => n61557, A2 => n16651, B1 => n61554, B2 => 
                           n16497, ZN => n9371);
   U9647 : AOI22_X1 port map( A1 => n61533, A2 => n16675, B1 => n61530, B2 => 
                           n16521, ZN => n9373);
   U9648 : AOI22_X1 port map( A1 => n61608, A2 => n1771, B1 => n61605, B2 => 
                           n1747, ZN => n9363);
   U9649 : AOI22_X1 port map( A1 => n61596, A2 => n15786, B1 => n61593, B2 => 
                           n15787, ZN => n9364);
   U9650 : AOI22_X1 port map( A1 => n61584, A2 => n4340, B1 => n61581, B2 => 
                           n4364, ZN => n9365);
   U9651 : AOI22_X1 port map( A1 => n61494, A2 => n648, B1 => n61491, B2 => 
                           n672, ZN => n9380);
   U9652 : AOI22_X1 port map( A1 => n61482, A2 => n600, B1 => n61479, B2 => 
                           n624, ZN => n9381);
   U9653 : AOI22_X1 port map( A1 => n61659, A2 => n4707, B1 => n61656, B2 => 
                           n944, ZN => n9355);
   U9654 : AOI22_X1 port map( A1 => n61635, A2 => n53484, B1 => n61632, B2 => 
                           n4560, ZN => n9357);
   U9655 : AOI22_X1 port map( A1 => n61353, A2 => n3011, B1 => n61350, B2 => 
                           n2987, ZN => n9407);
   U9656 : AOI22_X1 port map( A1 => n61341, A2 => n15397, B1 => n61338, B2 => 
                           n15435, ZN => n9408);
   U9657 : AOI22_X1 port map( A1 => n61329, A2 => n2895, B1 => n61326, B2 => 
                           n2447, ZN => n9409);
   U9658 : AOI22_X1 port map( A1 => n61380, A2 => n16110, B1 => n61377, B2 => 
                           n16111, ZN => n9401);
   U9659 : AOI22_X1 port map( A1 => n61404, A2 => n15785, B1 => n61401, B2 => 
                           n16545, ZN => n9399);
   U9660 : AOI22_X1 port map( A1 => n61392, A2 => n59656, B1 => n61389, B2 => 
                           n59701, ZN => n9400);
   U9661 : AOI22_X1 port map( A1 => n61290, A2 => n2303, B1 => n61287, B2 => 
                           n2327, ZN => n9416);
   U9662 : AOI22_X1 port map( A1 => n61278, A2 => n15511, B1 => n61275, B2 => 
                           n15455, ZN => n9417);
   U9663 : AOI22_X1 port map( A1 => n61455, A2 => n54332, B1 => n61452, B2 => 
                           n54356, ZN => n9391);
   U9664 : AOI22_X1 port map( A1 => n61443, A2 => n54486, B1 => n61440, B2 => 
                           n54630, ZN => n9392);
   U9665 : AOI22_X1 port map( A1 => n61431, A2 => n54236, B1 => n61428, B2 => 
                           n54260, ZN => n9393);
   U9666 : AOI22_X1 port map( A1 => n61557, A2 => n16652, B1 => n61554, B2 => 
                           n16498, ZN => n9232);
   U9667 : AOI22_X1 port map( A1 => n61533, A2 => n16676, B1 => n61530, B2 => 
                           n16522, ZN => n9234);
   U9668 : AOI22_X1 port map( A1 => n61608, A2 => n1770, B1 => n61605, B2 => 
                           n1746, ZN => n9224);
   U9669 : AOI22_X1 port map( A1 => n61596, A2 => n15791, B1 => n61593, B2 => 
                           n15792, ZN => n9225);
   U9670 : AOI22_X1 port map( A1 => n61584, A2 => n4339, B1 => n61581, B2 => 
                           n4363, ZN => n9226);
   U9671 : AOI22_X1 port map( A1 => n61494, A2 => n647, B1 => n61491, B2 => 
                           n671, ZN => n9241);
   U9672 : AOI22_X1 port map( A1 => n61482, A2 => n599, B1 => n61479, B2 => 
                           n623, ZN => n9242);
   U9673 : AOI22_X1 port map( A1 => n61659, A2 => n4706, B1 => n61656, B2 => 
                           n943, ZN => n9216);
   U9674 : AOI22_X1 port map( A1 => n61635, A2 => n53483, B1 => n61632, B2 => 
                           n4559, ZN => n9218);
   U9675 : AOI22_X1 port map( A1 => n61353, A2 => n3010, B1 => n61350, B2 => 
                           n2986, ZN => n9268);
   U9676 : AOI22_X1 port map( A1 => n61341, A2 => n15398, B1 => n61338, B2 => 
                           n15436, ZN => n9269);
   U9677 : AOI22_X1 port map( A1 => n61329, A2 => n2894, B1 => n61326, B2 => 
                           n2446, ZN => n9270);
   U9678 : AOI22_X1 port map( A1 => n61380, A2 => n16112, B1 => n61377, B2 => 
                           n16113, ZN => n9262);
   U9679 : AOI22_X1 port map( A1 => n61404, A2 => n15790, B1 => n61401, B2 => 
                           n16546, ZN => n9260);
   U9680 : AOI22_X1 port map( A1 => n61392, A2 => n59657, B1 => n61389, B2 => 
                           n59702, ZN => n9261);
   U9681 : AOI22_X1 port map( A1 => n61290, A2 => n2302, B1 => n61287, B2 => 
                           n2326, ZN => n9277);
   U9682 : AOI22_X1 port map( A1 => n61278, A2 => n15512, B1 => n61275, B2 => 
                           n15456, ZN => n9278);
   U9683 : AOI22_X1 port map( A1 => n61455, A2 => n54331, B1 => n61452, B2 => 
                           n54355, ZN => n9252);
   U9684 : AOI22_X1 port map( A1 => n61443, A2 => n54487, B1 => n61440, B2 => 
                           n54631, ZN => n9253);
   U9685 : AOI22_X1 port map( A1 => n61431, A2 => n54235, B1 => n61428, B2 => 
                           n54259, ZN => n9254);
   U9686 : AOI22_X1 port map( A1 => n61557, A2 => n16653, B1 => n61554, B2 => 
                           n16499, ZN => n9157);
   U9687 : AOI22_X1 port map( A1 => n61533, A2 => n16677, B1 => n61530, B2 => 
                           n16523, ZN => n9159);
   U9688 : AOI22_X1 port map( A1 => n61608, A2 => n1769, B1 => n61605, B2 => 
                           n1745, ZN => n9149);
   U9689 : AOI22_X1 port map( A1 => n61596, A2 => n15796, B1 => n61593, B2 => 
                           n15797, ZN => n9150);
   U9690 : AOI22_X1 port map( A1 => n61584, A2 => n4338, B1 => n61581, B2 => 
                           n4362, ZN => n9151);
   U9691 : AOI22_X1 port map( A1 => n61494, A2 => n646, B1 => n61491, B2 => 
                           n670, ZN => n9166);
   U9692 : AOI22_X1 port map( A1 => n61482, A2 => n598, B1 => n61479, B2 => 
                           n622, ZN => n9167);
   U9693 : AOI22_X1 port map( A1 => n61659, A2 => n4705, B1 => n61656, B2 => 
                           n942, ZN => n9141);
   U9694 : AOI22_X1 port map( A1 => n61635, A2 => n53482, B1 => n61632, B2 => 
                           n4558, ZN => n9143);
   U9695 : AOI22_X1 port map( A1 => n61353, A2 => n3009, B1 => n61350, B2 => 
                           n2985, ZN => n9193);
   U9696 : AOI22_X1 port map( A1 => n61341, A2 => n15399, B1 => n61338, B2 => 
                           n15437, ZN => n9194);
   U9697 : AOI22_X1 port map( A1 => n61329, A2 => n2893, B1 => n61326, B2 => 
                           n2445, ZN => n9195);
   U9698 : AOI22_X1 port map( A1 => n61380, A2 => n16114, B1 => n61377, B2 => 
                           n16115, ZN => n9187);
   U9699 : AOI22_X1 port map( A1 => n61404, A2 => n15795, B1 => n61401, B2 => 
                           n16547, ZN => n9185);
   U9700 : AOI22_X1 port map( A1 => n61392, A2 => n59658, B1 => n61389, B2 => 
                           n59703, ZN => n9186);
   U9701 : AOI22_X1 port map( A1 => n61290, A2 => n2301, B1 => n61287, B2 => 
                           n2325, ZN => n9202);
   U9702 : AOI22_X1 port map( A1 => n61278, A2 => n15513, B1 => n61275, B2 => 
                           n15457, ZN => n9203);
   U9703 : AOI22_X1 port map( A1 => n61455, A2 => n54330, B1 => n61452, B2 => 
                           n54354, ZN => n9177);
   U9704 : AOI22_X1 port map( A1 => n61443, A2 => n54488, B1 => n61440, B2 => 
                           n54632, ZN => n9178);
   U9705 : AOI22_X1 port map( A1 => n61431, A2 => n54234, B1 => n61428, B2 => 
                           n54258, ZN => n9179);
   U9706 : AOI22_X1 port map( A1 => n61557, A2 => n16654, B1 => n61554, B2 => 
                           n16500, ZN => n9082);
   U9707 : AOI22_X1 port map( A1 => n61533, A2 => n16678, B1 => n61530, B2 => 
                           n16524, ZN => n9084);
   U9708 : AOI22_X1 port map( A1 => n61608, A2 => n1768, B1 => n61605, B2 => 
                           n1744, ZN => n9074);
   U9709 : AOI22_X1 port map( A1 => n61596, A2 => n15801, B1 => n61593, B2 => 
                           n15802, ZN => n9075);
   U9710 : AOI22_X1 port map( A1 => n61584, A2 => n4337, B1 => n61581, B2 => 
                           n4361, ZN => n9076);
   U9711 : AOI22_X1 port map( A1 => n61494, A2 => n645, B1 => n61491, B2 => 
                           n669, ZN => n9091);
   U9712 : AOI22_X1 port map( A1 => n61482, A2 => n597, B1 => n61479, B2 => 
                           n621, ZN => n9092);
   U9713 : AOI22_X1 port map( A1 => n61659, A2 => n4704, B1 => n61656, B2 => 
                           n941, ZN => n9066);
   U9714 : AOI22_X1 port map( A1 => n61635, A2 => n53481, B1 => n61632, B2 => 
                           n4557, ZN => n9068);
   U9715 : AOI22_X1 port map( A1 => n61353, A2 => n3008, B1 => n61350, B2 => 
                           n2984, ZN => n9118);
   U9716 : AOI22_X1 port map( A1 => n61341, A2 => n15400, B1 => n61338, B2 => 
                           n15438, ZN => n9119);
   U9717 : AOI22_X1 port map( A1 => n61329, A2 => n2892, B1 => n61326, B2 => 
                           n2444, ZN => n9120);
   U9718 : AOI22_X1 port map( A1 => n61380, A2 => n16116, B1 => n61377, B2 => 
                           n16117, ZN => n9112);
   U9719 : AOI22_X1 port map( A1 => n61404, A2 => n15800, B1 => n61401, B2 => 
                           n16548, ZN => n9110);
   U9720 : AOI22_X1 port map( A1 => n61392, A2 => n59659, B1 => n61389, B2 => 
                           n59704, ZN => n9111);
   U9721 : AOI22_X1 port map( A1 => n61290, A2 => n2300, B1 => n61287, B2 => 
                           n2324, ZN => n9127);
   U9722 : AOI22_X1 port map( A1 => n61278, A2 => n15514, B1 => n61275, B2 => 
                           n15458, ZN => n9128);
   U9723 : AOI22_X1 port map( A1 => n61455, A2 => n54329, B1 => n61452, B2 => 
                           n54353, ZN => n9102);
   U9724 : AOI22_X1 port map( A1 => n61443, A2 => n54489, B1 => n61440, B2 => 
                           n54633, ZN => n9103);
   U9725 : AOI22_X1 port map( A1 => n61431, A2 => n54233, B1 => n61428, B2 => 
                           n54257, ZN => n9104);
   U9726 : AOI22_X1 port map( A1 => n61557, A2 => n16655, B1 => n61554, B2 => 
                           n16501, ZN => n9007);
   U9727 : AOI22_X1 port map( A1 => n61533, A2 => n16679, B1 => n61530, B2 => 
                           n16525, ZN => n9009);
   U9728 : AOI22_X1 port map( A1 => n61608, A2 => n1767, B1 => n61605, B2 => 
                           n1743, ZN => n8999);
   U9729 : AOI22_X1 port map( A1 => n61596, A2 => n15854, B1 => n61593, B2 => 
                           n15855, ZN => n9000);
   U9730 : AOI22_X1 port map( A1 => n61584, A2 => n4336, B1 => n61581, B2 => 
                           n4360, ZN => n9001);
   U9731 : AOI22_X1 port map( A1 => n61494, A2 => n644, B1 => n61491, B2 => 
                           n668, ZN => n9016);
   U9732 : AOI22_X1 port map( A1 => n61482, A2 => n596, B1 => n61479, B2 => 
                           n620, ZN => n9017);
   U9733 : AOI22_X1 port map( A1 => n61659, A2 => n4703, B1 => n61656, B2 => 
                           n940, ZN => n8991);
   U9734 : AOI22_X1 port map( A1 => n61635, A2 => n53480, B1 => n61632, B2 => 
                           n4556, ZN => n8993);
   U9735 : AOI22_X1 port map( A1 => n61353, A2 => n3007, B1 => n61350, B2 => 
                           n2983, ZN => n9043);
   U9736 : AOI22_X1 port map( A1 => n61341, A2 => n15401, B1 => n61338, B2 => 
                           n15439, ZN => n9044);
   U9737 : AOI22_X1 port map( A1 => n61329, A2 => n2891, B1 => n61326, B2 => 
                           n2443, ZN => n9045);
   U9738 : AOI22_X1 port map( A1 => n61380, A2 => n16118, B1 => n61377, B2 => 
                           n16119, ZN => n9037);
   U9739 : AOI22_X1 port map( A1 => n61404, A2 => n15853, B1 => n61401, B2 => 
                           n16549, ZN => n9035);
   U9740 : AOI22_X1 port map( A1 => n61392, A2 => n59660, B1 => n61389, B2 => 
                           n59705, ZN => n9036);
   U9741 : AOI22_X1 port map( A1 => n61290, A2 => n2299, B1 => n61287, B2 => 
                           n2323, ZN => n9052);
   U9742 : AOI22_X1 port map( A1 => n61278, A2 => n15515, B1 => n61275, B2 => 
                           n15459, ZN => n9053);
   U9743 : AOI22_X1 port map( A1 => n61455, A2 => n54328, B1 => n61452, B2 => 
                           n54352, ZN => n9027);
   U9744 : AOI22_X1 port map( A1 => n61443, A2 => n54490, B1 => n61440, B2 => 
                           n54634, ZN => n9028);
   U9745 : AOI22_X1 port map( A1 => n61431, A2 => n54232, B1 => n61428, B2 => 
                           n54256, ZN => n9029);
   U9746 : AOI22_X1 port map( A1 => n61557, A2 => n16656, B1 => n61553, B2 => 
                           n16502, ZN => n8932);
   U9747 : AOI22_X1 port map( A1 => n61533, A2 => n16680, B1 => n61529, B2 => 
                           n16526, ZN => n8934);
   U9748 : AOI22_X1 port map( A1 => n61608, A2 => n1766, B1 => n61604, B2 => 
                           n1742, ZN => n8924);
   U9749 : AOI22_X1 port map( A1 => n61596, A2 => n15859, B1 => n61592, B2 => 
                           n15860, ZN => n8925);
   U9750 : AOI22_X1 port map( A1 => n61584, A2 => n4335, B1 => n61580, B2 => 
                           n4359, ZN => n8926);
   U9751 : AOI22_X1 port map( A1 => n61494, A2 => n643, B1 => n61490, B2 => 
                           n667, ZN => n8941);
   U9752 : AOI22_X1 port map( A1 => n61482, A2 => n595, B1 => n61478, B2 => 
                           n619, ZN => n8942);
   U9753 : AOI22_X1 port map( A1 => n61659, A2 => n4702, B1 => n61655, B2 => 
                           n939, ZN => n8916);
   U9754 : AOI22_X1 port map( A1 => n61635, A2 => n53479, B1 => n61631, B2 => 
                           n4555, ZN => n8918);
   U9755 : AOI22_X1 port map( A1 => n61353, A2 => n3006, B1 => n61349, B2 => 
                           n2982, ZN => n8968);
   U9756 : AOI22_X1 port map( A1 => n61341, A2 => n15697, B1 => n61337, B2 => 
                           n16560, ZN => n8969);
   U9757 : AOI22_X1 port map( A1 => n61329, A2 => n2890, B1 => n61325, B2 => 
                           n2442, ZN => n8970);
   U9758 : AOI22_X1 port map( A1 => n61380, A2 => n16100, B1 => n61376, B2 => 
                           n16101, ZN => n8962);
   U9759 : AOI22_X1 port map( A1 => n61404, A2 => n15858, B1 => n61400, B2 => 
                           n16550, ZN => n8960);
   U9760 : AOI22_X1 port map( A1 => n61392, A2 => n59661, B1 => n61388, B2 => 
                           n59706, ZN => n8961);
   U9761 : AOI22_X1 port map( A1 => n61290, A2 => n999, B1 => n61286, B2 => 
                           n2322, ZN => n8977);
   U9762 : AOI22_X1 port map( A1 => n61278, A2 => n15516, B1 => n61274, B2 => 
                           n15460, ZN => n8978);
   U9763 : AOI22_X1 port map( A1 => n61455, A2 => n54327, B1 => n61451, B2 => 
                           n54351, ZN => n8952);
   U9764 : AOI22_X1 port map( A1 => n61443, A2 => n54491, B1 => n61439, B2 => 
                           n54635, ZN => n8953);
   U9765 : AOI22_X1 port map( A1 => n61431, A2 => n54231, B1 => n61427, B2 => 
                           n54255, ZN => n8954);
   U9766 : AOI22_X1 port map( A1 => n61557, A2 => n16657, B1 => n61553, B2 => 
                           n16503, ZN => n8857);
   U9767 : AOI22_X1 port map( A1 => n61533, A2 => n16681, B1 => n61529, B2 => 
                           n16527, ZN => n8859);
   U9768 : AOI22_X1 port map( A1 => n61608, A2 => n1765, B1 => n61604, B2 => 
                           n1741, ZN => n8849);
   U9769 : AOI22_X1 port map( A1 => n61596, A2 => n15864, B1 => n61592, B2 => 
                           n15865, ZN => n8850);
   U9770 : AOI22_X1 port map( A1 => n61584, A2 => n4334, B1 => n61580, B2 => 
                           n4358, ZN => n8851);
   U9771 : AOI22_X1 port map( A1 => n61494, A2 => n642, B1 => n61490, B2 => 
                           n666, ZN => n8866);
   U9772 : AOI22_X1 port map( A1 => n61482, A2 => n594, B1 => n61478, B2 => 
                           n618, ZN => n8867);
   U9773 : AOI22_X1 port map( A1 => n61659, A2 => n4701, B1 => n61655, B2 => 
                           n938, ZN => n8841);
   U9774 : AOI22_X1 port map( A1 => n61635, A2 => n53478, B1 => n61631, B2 => 
                           n4554, ZN => n8843);
   U9775 : AOI22_X1 port map( A1 => n61353, A2 => n3005, B1 => n61349, B2 => 
                           n2981, ZN => n8893);
   U9776 : AOI22_X1 port map( A1 => n61341, A2 => n15700, B1 => n61337, B2 => 
                           n16561, ZN => n8894);
   U9777 : AOI22_X1 port map( A1 => n61329, A2 => n2889, B1 => n61325, B2 => 
                           n2441, ZN => n8895);
   U9778 : AOI22_X1 port map( A1 => n61380, A2 => n16102, B1 => n61376, B2 => 
                           n16103, ZN => n8887);
   U9779 : AOI22_X1 port map( A1 => n61404, A2 => n15863, B1 => n61400, B2 => 
                           n16551, ZN => n8885);
   U9780 : AOI22_X1 port map( A1 => n61392, A2 => n59662, B1 => n61388, B2 => 
                           n59707, ZN => n8886);
   U9781 : AOI22_X1 port map( A1 => n61290, A2 => n998, B1 => n61286, B2 => 
                           n2321, ZN => n8902);
   U9782 : AOI22_X1 port map( A1 => n61278, A2 => n15517, B1 => n61274, B2 => 
                           n15461, ZN => n8903);
   U9783 : AOI22_X1 port map( A1 => n61455, A2 => n54326, B1 => n61451, B2 => 
                           n54350, ZN => n8877);
   U9784 : AOI22_X1 port map( A1 => n61443, A2 => n54492, B1 => n61439, B2 => 
                           n54636, ZN => n8878);
   U9785 : AOI22_X1 port map( A1 => n61431, A2 => n54230, B1 => n61427, B2 => 
                           n54254, ZN => n8879);
   U9786 : AOI22_X1 port map( A1 => n61557, A2 => n16658, B1 => n61553, B2 => 
                           n16504, ZN => n8782);
   U9787 : AOI22_X1 port map( A1 => n61533, A2 => n16682, B1 => n61529, B2 => 
                           n16528, ZN => n8784);
   U9788 : AOI22_X1 port map( A1 => n61608, A2 => n1764, B1 => n61604, B2 => 
                           n1740, ZN => n8774);
   U9789 : AOI22_X1 port map( A1 => n61596, A2 => n15869, B1 => n61592, B2 => 
                           n15870, ZN => n8775);
   U9790 : AOI22_X1 port map( A1 => n61584, A2 => n4333, B1 => n61580, B2 => 
                           n4357, ZN => n8776);
   U9791 : AOI22_X1 port map( A1 => n61494, A2 => n641, B1 => n61490, B2 => 
                           n665, ZN => n8791);
   U9792 : AOI22_X1 port map( A1 => n61482, A2 => n593, B1 => n61478, B2 => 
                           n617, ZN => n8792);
   U9793 : AOI22_X1 port map( A1 => n61659, A2 => n4700, B1 => n61655, B2 => 
                           n937, ZN => n8766);
   U9794 : AOI22_X1 port map( A1 => n61635, A2 => n53477, B1 => n61631, B2 => 
                           n4553, ZN => n8768);
   U9795 : AOI22_X1 port map( A1 => n61353, A2 => n3004, B1 => n61349, B2 => 
                           n2980, ZN => n8818);
   U9796 : AOI22_X1 port map( A1 => n61341, A2 => n15703, B1 => n61337, B2 => 
                           n16562, ZN => n8819);
   U9797 : AOI22_X1 port map( A1 => n61329, A2 => n2888, B1 => n61325, B2 => 
                           n2440, ZN => n8820);
   U9798 : AOI22_X1 port map( A1 => n61380, A2 => n16104, B1 => n61376, B2 => 
                           n16105, ZN => n8812);
   U9799 : AOI22_X1 port map( A1 => n61404, A2 => n15868, B1 => n61400, B2 => 
                           n16552, ZN => n8810);
   U9800 : AOI22_X1 port map( A1 => n61392, A2 => n59663, B1 => n61388, B2 => 
                           n59708, ZN => n8811);
   U9801 : AOI22_X1 port map( A1 => n61290, A2 => n997, B1 => n61286, B2 => 
                           n2320, ZN => n8827);
   U9802 : AOI22_X1 port map( A1 => n61278, A2 => n15518, B1 => n61274, B2 => 
                           n15462, ZN => n8828);
   U9803 : AOI22_X1 port map( A1 => n61455, A2 => n54325, B1 => n61451, B2 => 
                           n54349, ZN => n8802);
   U9804 : AOI22_X1 port map( A1 => n61443, A2 => n54493, B1 => n61439, B2 => 
                           n54637, ZN => n8803);
   U9805 : AOI22_X1 port map( A1 => n61431, A2 => n54229, B1 => n61427, B2 => 
                           n54253, ZN => n8804);
   U9806 : AOI22_X1 port map( A1 => n61557, A2 => n16659, B1 => n61553, B2 => 
                           n16505, ZN => n8707);
   U9807 : AOI22_X1 port map( A1 => n61533, A2 => n16683, B1 => n61529, B2 => 
                           n16529, ZN => n8709);
   U9808 : AOI22_X1 port map( A1 => n61608, A2 => n1763, B1 => n61604, B2 => 
                           n1739, ZN => n8699);
   U9809 : AOI22_X1 port map( A1 => n61596, A2 => n15874, B1 => n61592, B2 => 
                           n15875, ZN => n8700);
   U9810 : AOI22_X1 port map( A1 => n61584, A2 => n4332, B1 => n61580, B2 => 
                           n4356, ZN => n8701);
   U9811 : AOI22_X1 port map( A1 => n61494, A2 => n640, B1 => n61490, B2 => 
                           n664, ZN => n8716);
   U9812 : AOI22_X1 port map( A1 => n61482, A2 => n592, B1 => n61478, B2 => 
                           n616, ZN => n8717);
   U9813 : AOI22_X1 port map( A1 => n61659, A2 => n4699, B1 => n61655, B2 => 
                           n936, ZN => n8691);
   U9814 : AOI22_X1 port map( A1 => n61635, A2 => n53476, B1 => n61631, B2 => 
                           n4552, ZN => n8693);
   U9815 : AOI22_X1 port map( A1 => n61353, A2 => n3003, B1 => n61349, B2 => 
                           n2979, ZN => n8743);
   U9816 : AOI22_X1 port map( A1 => n61341, A2 => n15706, B1 => n61337, B2 => 
                           n16563, ZN => n8744);
   U9817 : AOI22_X1 port map( A1 => n61329, A2 => n2887, B1 => n61325, B2 => 
                           n2439, ZN => n8745);
   U9818 : AOI22_X1 port map( A1 => n61380, A2 => n16106, B1 => n61376, B2 => 
                           n16107, ZN => n8737);
   U9819 : AOI22_X1 port map( A1 => n61404, A2 => n15873, B1 => n61400, B2 => 
                           n16553, ZN => n8735);
   U9820 : AOI22_X1 port map( A1 => n61392, A2 => n59664, B1 => n61388, B2 => 
                           n59709, ZN => n8736);
   U9821 : AOI22_X1 port map( A1 => n61290, A2 => n996, B1 => n61286, B2 => 
                           n2319, ZN => n8752);
   U9822 : AOI22_X1 port map( A1 => n61278, A2 => n15519, B1 => n61274, B2 => 
                           n15463, ZN => n8753);
   U9823 : AOI22_X1 port map( A1 => n61455, A2 => n54324, B1 => n61451, B2 => 
                           n54348, ZN => n8727);
   U9824 : AOI22_X1 port map( A1 => n61443, A2 => n54494, B1 => n61439, B2 => 
                           n54638, ZN => n8728);
   U9825 : AOI22_X1 port map( A1 => n61431, A2 => n54228, B1 => n61427, B2 => 
                           n54252, ZN => n8729);
   U9826 : AOI22_X1 port map( A1 => n61558, A2 => n16830, B1 => n61553, B2 => 
                           n16831, ZN => n8632);
   U9827 : AOI22_X1 port map( A1 => n61546, A2 => n4272, B1 => n61541, B2 => 
                           n4264, ZN => n8633);
   U9828 : AOI22_X1 port map( A1 => n61534, A2 => n16437, B1 => n61529, B2 => 
                           n16445, ZN => n8634);
   U9829 : AOI22_X1 port map( A1 => n61609, A2 => n127, B1 => n61604, B2 => 
                           n119, ZN => n8624);
   U9830 : AOI22_X1 port map( A1 => n61597, A2 => n15918, B1 => n61592, B2 => 
                           n15919, ZN => n8625);
   U9831 : AOI22_X1 port map( A1 => n61585, A2 => n3963, B1 => n61580, B2 => 
                           n3995, ZN => n8626);
   U9832 : AOI22_X1 port map( A1 => n61495, A2 => n530, B1 => n61490, B2 => 
                           n538, ZN => n8641);
   U9833 : AOI22_X1 port map( A1 => n61483, A2 => n513, B1 => n61478, B2 => 
                           n522, ZN => n8642);
   U9834 : AOI22_X1 port map( A1 => n61660, A2 => n4179, B1 => n61655, B2 => 
                           n4171, ZN => n8616);
   U9835 : AOI22_X1 port map( A1 => n61648, A2 => n51631, B1 => n61643, B2 => 
                           n51655, ZN => n8617);
   U9836 : AOI22_X1 port map( A1 => n61636, A2 => n51623, B1 => n61631, B2 => 
                           n51615, ZN => n8618);
   U9837 : AOI22_X1 port map( A1 => n61354, A2 => n387, B1 => n61349, B2 => 
                           n379, ZN => n8668);
   U9838 : AOI22_X1 port map( A1 => n61342, A2 => n15316, B1 => n61337, B2 => 
                           n15324, ZN => n8669);
   U9839 : AOI22_X1 port map( A1 => n61330, A2 => n355, B1 => n61325, B2 => 
                           n347, ZN => n8670);
   U9840 : AOI22_X1 port map( A1 => n61381, A2 => n50971, B1 => n61376, B2 => 
                           n50939, ZN => n8662);
   U9841 : AOI22_X1 port map( A1 => n61405, A2 => n51719, B1 => n61400, B2 => 
                           n51727, ZN => n8660);
   U9842 : AOI22_X1 port map( A1 => n61393, A2 => n15467, B1 => n61388, B2 => 
                           n15475, ZN => n8661);
   U9843 : AOI22_X1 port map( A1 => n61291, A2 => n4296, B1 => n61286, B2 => 
                           n4304, ZN => n8677);
   U9844 : AOI22_X1 port map( A1 => n61279, A2 => n16469, B1 => n61274, B2 => 
                           n15675, ZN => n8678);
   U9845 : AOI22_X1 port map( A1 => n61456, A2 => n51767, B1 => n61451, B2 => 
                           n51775, ZN => n8652);
   U9846 : AOI22_X1 port map( A1 => n61444, A2 => n451, B1 => n61439, B2 => 
                           n443, ZN => n8653);
   U9847 : AOI22_X1 port map( A1 => n61432, A2 => n51735, B1 => n61427, B2 => 
                           n51743, ZN => n8654);
   U9848 : AOI22_X1 port map( A1 => n61558, A2 => n16832, B1 => n61553, B2 => 
                           n16833, ZN => n8557);
   U9849 : AOI22_X1 port map( A1 => n61546, A2 => n4271, B1 => n61541, B2 => 
                           n4263, ZN => n8558);
   U9850 : AOI22_X1 port map( A1 => n61534, A2 => n16438, B1 => n61529, B2 => 
                           n16446, ZN => n8559);
   U9851 : AOI22_X1 port map( A1 => n61609, A2 => n126, B1 => n61604, B2 => 
                           n118, ZN => n8549);
   U9852 : AOI22_X1 port map( A1 => n61597, A2 => n15922, B1 => n61592, B2 => 
                           n15947, ZN => n8550);
   U9853 : AOI22_X1 port map( A1 => n61585, A2 => n3962, B1 => n61580, B2 => 
                           n3994, ZN => n8551);
   U9854 : AOI22_X1 port map( A1 => n61495, A2 => n529, B1 => n61490, B2 => 
                           n537, ZN => n8566);
   U9855 : AOI22_X1 port map( A1 => n61483, A2 => n512, B1 => n61478, B2 => 
                           n521, ZN => n8567);
   U9856 : AOI22_X1 port map( A1 => n61660, A2 => n4178, B1 => n61655, B2 => 
                           n4170, ZN => n8541);
   U9857 : AOI22_X1 port map( A1 => n61648, A2 => n51630, B1 => n61643, B2 => 
                           n51654, ZN => n8542);
   U9858 : AOI22_X1 port map( A1 => n61636, A2 => n51622, B1 => n61631, B2 => 
                           n51614, ZN => n8543);
   U9859 : AOI22_X1 port map( A1 => n61354, A2 => n386, B1 => n61349, B2 => 
                           n378, ZN => n8593);
   U9860 : AOI22_X1 port map( A1 => n61342, A2 => n15317, B1 => n61337, B2 => 
                           n15325, ZN => n8594);
   U9861 : AOI22_X1 port map( A1 => n61330, A2 => n354, B1 => n61325, B2 => 
                           n346, ZN => n8595);
   U9862 : AOI22_X1 port map( A1 => n61381, A2 => n50970, B1 => n61376, B2 => 
                           n50938, ZN => n8587);
   U9863 : AOI22_X1 port map( A1 => n61405, A2 => n51718, B1 => n61400, B2 => 
                           n51726, ZN => n8585);
   U9864 : AOI22_X1 port map( A1 => n61393, A2 => n15468, B1 => n61388, B2 => 
                           n15476, ZN => n8586);
   U9865 : AOI22_X1 port map( A1 => n61291, A2 => n4295, B1 => n61286, B2 => 
                           n4303, ZN => n8602);
   U9866 : AOI22_X1 port map( A1 => n61279, A2 => n16470, B1 => n61274, B2 => 
                           n15678, ZN => n8603);
   U9867 : AOI22_X1 port map( A1 => n61456, A2 => n51766, B1 => n61451, B2 => 
                           n51774, ZN => n8577);
   U9868 : AOI22_X1 port map( A1 => n61444, A2 => n450, B1 => n61439, B2 => 
                           n442, ZN => n8578);
   U9869 : AOI22_X1 port map( A1 => n61432, A2 => n51734, B1 => n61427, B2 => 
                           n51742, ZN => n8579);
   U9870 : AOI22_X1 port map( A1 => n61558, A2 => n16834, B1 => n61553, B2 => 
                           n16835, ZN => n8482);
   U9871 : AOI22_X1 port map( A1 => n61546, A2 => n4270, B1 => n61541, B2 => 
                           n4262, ZN => n8483);
   U9872 : AOI22_X1 port map( A1 => n61534, A2 => n16439, B1 => n61529, B2 => 
                           n16447, ZN => n8484);
   U9873 : AOI22_X1 port map( A1 => n61609, A2 => n125, B1 => n61604, B2 => 
                           n117, ZN => n8474);
   U9874 : AOI22_X1 port map( A1 => n61597, A2 => n15950, B1 => n61592, B2 => 
                           n15951, ZN => n8475);
   U9875 : AOI22_X1 port map( A1 => n61585, A2 => n3961, B1 => n61580, B2 => 
                           n3993, ZN => n8476);
   U9876 : AOI22_X1 port map( A1 => n61495, A2 => n528, B1 => n61490, B2 => 
                           n536, ZN => n8491);
   U9877 : AOI22_X1 port map( A1 => n61483, A2 => n511, B1 => n61478, B2 => 
                           n520, ZN => n8492);
   U9878 : AOI22_X1 port map( A1 => n61660, A2 => n4177, B1 => n61655, B2 => 
                           n4169, ZN => n8466);
   U9879 : AOI22_X1 port map( A1 => n61648, A2 => n51629, B1 => n61643, B2 => 
                           n51653, ZN => n8467);
   U9880 : AOI22_X1 port map( A1 => n61636, A2 => n51621, B1 => n61631, B2 => 
                           n51613, ZN => n8468);
   U9881 : AOI22_X1 port map( A1 => n61354, A2 => n385, B1 => n61349, B2 => 
                           n377, ZN => n8518);
   U9882 : AOI22_X1 port map( A1 => n61342, A2 => n15318, B1 => n61337, B2 => 
                           n15326, ZN => n8519);
   U9883 : AOI22_X1 port map( A1 => n61330, A2 => n353, B1 => n61325, B2 => 
                           n345, ZN => n8520);
   U9884 : AOI22_X1 port map( A1 => n61381, A2 => n50969, B1 => n61376, B2 => 
                           n50937, ZN => n8512);
   U9885 : AOI22_X1 port map( A1 => n61405, A2 => n51717, B1 => n61400, B2 => 
                           n51725, ZN => n8510);
   U9886 : AOI22_X1 port map( A1 => n61393, A2 => n15469, B1 => n61388, B2 => 
                           n15477, ZN => n8511);
   U9887 : AOI22_X1 port map( A1 => n61291, A2 => n4294, B1 => n61286, B2 => 
                           n4302, ZN => n8527);
   U9888 : AOI22_X1 port map( A1 => n61279, A2 => n16471, B1 => n61274, B2 => 
                           n15681, ZN => n8528);
   U9889 : AOI22_X1 port map( A1 => n61456, A2 => n51765, B1 => n61451, B2 => 
                           n51773, ZN => n8502);
   U9890 : AOI22_X1 port map( A1 => n61444, A2 => n449, B1 => n61439, B2 => 
                           n441, ZN => n8503);
   U9891 : AOI22_X1 port map( A1 => n61432, A2 => n51733, B1 => n61427, B2 => 
                           n51741, ZN => n8504);
   U9892 : AOI22_X1 port map( A1 => n61558, A2 => n16836, B1 => n61553, B2 => 
                           n16837, ZN => n8407);
   U9893 : AOI22_X1 port map( A1 => n61546, A2 => n4269, B1 => n61541, B2 => 
                           n4261, ZN => n8408);
   U9894 : AOI22_X1 port map( A1 => n61534, A2 => n16440, B1 => n61529, B2 => 
                           n16448, ZN => n8409);
   U9895 : AOI22_X1 port map( A1 => n61609, A2 => n124, B1 => n61604, B2 => 
                           n116, ZN => n8399);
   U9896 : AOI22_X1 port map( A1 => n61597, A2 => n15954, B1 => n61592, B2 => 
                           n15955, ZN => n8400);
   U9897 : AOI22_X1 port map( A1 => n61585, A2 => n3960, B1 => n61580, B2 => 
                           n3992, ZN => n8401);
   U9898 : AOI22_X1 port map( A1 => n61495, A2 => n527, B1 => n61490, B2 => 
                           n535, ZN => n8416);
   U9899 : AOI22_X1 port map( A1 => n61483, A2 => n510, B1 => n61478, B2 => 
                           n518, ZN => n8417);
   U9900 : AOI22_X1 port map( A1 => n61660, A2 => n4176, B1 => n61655, B2 => 
                           n4168, ZN => n8391);
   U9901 : AOI22_X1 port map( A1 => n61648, A2 => n51628, B1 => n61643, B2 => 
                           n51652, ZN => n8392);
   U9902 : AOI22_X1 port map( A1 => n61636, A2 => n51620, B1 => n61631, B2 => 
                           n51612, ZN => n8393);
   U9903 : AOI22_X1 port map( A1 => n61354, A2 => n384, B1 => n61349, B2 => 
                           n376, ZN => n8443);
   U9904 : AOI22_X1 port map( A1 => n61342, A2 => n15319, B1 => n61337, B2 => 
                           n15327, ZN => n8444);
   U9905 : AOI22_X1 port map( A1 => n61330, A2 => n352, B1 => n61325, B2 => 
                           n344, ZN => n8445);
   U9906 : AOI22_X1 port map( A1 => n61381, A2 => n50968, B1 => n61376, B2 => 
                           n50936, ZN => n8437);
   U9907 : AOI22_X1 port map( A1 => n61405, A2 => n51716, B1 => n61400, B2 => 
                           n51724, ZN => n8435);
   U9908 : AOI22_X1 port map( A1 => n61393, A2 => n15470, B1 => n61388, B2 => 
                           n15478, ZN => n8436);
   U9909 : AOI22_X1 port map( A1 => n61291, A2 => n4293, B1 => n61286, B2 => 
                           n4301, ZN => n8452);
   U9910 : AOI22_X1 port map( A1 => n61279, A2 => n16472, B1 => n61274, B2 => 
                           n15684, ZN => n8453);
   U9911 : AOI22_X1 port map( A1 => n61456, A2 => n51764, B1 => n61451, B2 => 
                           n51772, ZN => n8427);
   U9912 : AOI22_X1 port map( A1 => n61444, A2 => n448, B1 => n61439, B2 => 
                           n440, ZN => n8428);
   U9913 : AOI22_X1 port map( A1 => n61432, A2 => n51732, B1 => n61427, B2 => 
                           n51740, ZN => n8429);
   U9914 : AOI22_X1 port map( A1 => n61558, A2 => n16838, B1 => n61553, B2 => 
                           n16839, ZN => n8332);
   U9915 : AOI22_X1 port map( A1 => n61546, A2 => n4268, B1 => n61541, B2 => 
                           n4260, ZN => n8333);
   U9916 : AOI22_X1 port map( A1 => n61534, A2 => n16441, B1 => n61529, B2 => 
                           n16449, ZN => n8334);
   U9917 : AOI22_X1 port map( A1 => n61609, A2 => n123, B1 => n61604, B2 => 
                           n115, ZN => n8324);
   U9918 : AOI22_X1 port map( A1 => n61597, A2 => n15958, B1 => n61592, B2 => 
                           n15959, ZN => n8325);
   U9919 : AOI22_X1 port map( A1 => n61585, A2 => n3959, B1 => n61580, B2 => 
                           n3991, ZN => n8326);
   U9920 : AOI22_X1 port map( A1 => n61495, A2 => n526, B1 => n61490, B2 => 
                           n534, ZN => n8341);
   U9921 : AOI22_X1 port map( A1 => n61483, A2 => n509, B1 => n61478, B2 => 
                           n517, ZN => n8342);
   U9922 : AOI22_X1 port map( A1 => n61660, A2 => n4175, B1 => n61655, B2 => 
                           n4167, ZN => n8316);
   U9923 : AOI22_X1 port map( A1 => n61648, A2 => n51627, B1 => n61643, B2 => 
                           n51651, ZN => n8317);
   U9924 : AOI22_X1 port map( A1 => n61636, A2 => n51619, B1 => n61631, B2 => 
                           n51611, ZN => n8318);
   U9925 : AOI22_X1 port map( A1 => n61354, A2 => n383, B1 => n61349, B2 => 
                           n375, ZN => n8368);
   U9926 : AOI22_X1 port map( A1 => n61342, A2 => n15320, B1 => n61337, B2 => 
                           n15328, ZN => n8369);
   U9927 : AOI22_X1 port map( A1 => n61330, A2 => n351, B1 => n61325, B2 => 
                           n343, ZN => n8370);
   U9928 : AOI22_X1 port map( A1 => n61381, A2 => n50967, B1 => n61376, B2 => 
                           n50935, ZN => n8362);
   U9929 : AOI22_X1 port map( A1 => n61405, A2 => n51715, B1 => n61400, B2 => 
                           n51723, ZN => n8360);
   U9930 : AOI22_X1 port map( A1 => n61393, A2 => n15471, B1 => n61388, B2 => 
                           n15479, ZN => n8361);
   U9931 : AOI22_X1 port map( A1 => n61291, A2 => n4292, B1 => n61286, B2 => 
                           n4300, ZN => n8377);
   U9932 : AOI22_X1 port map( A1 => n61279, A2 => n16473, B1 => n61274, B2 => 
                           n15663, ZN => n8378);
   U9933 : AOI22_X1 port map( A1 => n61456, A2 => n51763, B1 => n61451, B2 => 
                           n51771, ZN => n8352);
   U9934 : AOI22_X1 port map( A1 => n61444, A2 => n447, B1 => n61439, B2 => 
                           n439, ZN => n8353);
   U9935 : AOI22_X1 port map( A1 => n61432, A2 => n51731, B1 => n61427, B2 => 
                           n51739, ZN => n8354);
   U9936 : AOI22_X1 port map( A1 => n61558, A2 => n16840, B1 => n61553, B2 => 
                           n16841, ZN => n8257);
   U9937 : AOI22_X1 port map( A1 => n61546, A2 => n4267, B1 => n61541, B2 => 
                           n4259, ZN => n8258);
   U9938 : AOI22_X1 port map( A1 => n61534, A2 => n16442, B1 => n61529, B2 => 
                           n16450, ZN => n8259);
   U9939 : AOI22_X1 port map( A1 => n61609, A2 => n122, B1 => n61604, B2 => 
                           n114, ZN => n8249);
   U9940 : AOI22_X1 port map( A1 => n61597, A2 => n15962, B1 => n61592, B2 => 
                           n15963, ZN => n8250);
   U9941 : AOI22_X1 port map( A1 => n61585, A2 => n3958, B1 => n61580, B2 => 
                           n3966, ZN => n8251);
   U9942 : AOI22_X1 port map( A1 => n61495, A2 => n525, B1 => n61490, B2 => 
                           n533, ZN => n8266);
   U9943 : AOI22_X1 port map( A1 => n61483, A2 => n508, B1 => n61478, B2 => 
                           n516, ZN => n8267);
   U9944 : AOI22_X1 port map( A1 => n61660, A2 => n4174, B1 => n61655, B2 => 
                           n4166, ZN => n8241);
   U9945 : AOI22_X1 port map( A1 => n61648, A2 => n51626, B1 => n61643, B2 => 
                           n51650, ZN => n8242);
   U9946 : AOI22_X1 port map( A1 => n61636, A2 => n51618, B1 => n61631, B2 => 
                           n51610, ZN => n8243);
   U9947 : AOI22_X1 port map( A1 => n61354, A2 => n382, B1 => n61349, B2 => 
                           n374, ZN => n8293);
   U9948 : AOI22_X1 port map( A1 => n61342, A2 => n15321, B1 => n61337, B2 => 
                           n15329, ZN => n8294);
   U9949 : AOI22_X1 port map( A1 => n61330, A2 => n350, B1 => n61325, B2 => 
                           n342, ZN => n8295);
   U9950 : AOI22_X1 port map( A1 => n61381, A2 => n50966, B1 => n61376, B2 => 
                           n50934, ZN => n8287);
   U9951 : AOI22_X1 port map( A1 => n61405, A2 => n51714, B1 => n61400, B2 => 
                           n51722, ZN => n8285);
   U9952 : AOI22_X1 port map( A1 => n61393, A2 => n15472, B1 => n61388, B2 => 
                           n15480, ZN => n8286);
   U9953 : AOI22_X1 port map( A1 => n61291, A2 => n4291, B1 => n61286, B2 => 
                           n4299, ZN => n8302);
   U9954 : AOI22_X1 port map( A1 => n61279, A2 => n16474, B1 => n61274, B2 => 
                           n15666, ZN => n8303);
   U9955 : AOI22_X1 port map( A1 => n61456, A2 => n51762, B1 => n61451, B2 => 
                           n51770, ZN => n8277);
   U9956 : AOI22_X1 port map( A1 => n61444, A2 => n446, B1 => n61439, B2 => 
                           n438, ZN => n8278);
   U9957 : AOI22_X1 port map( A1 => n61432, A2 => n51730, B1 => n61427, B2 => 
                           n51738, ZN => n8279);
   U9958 : AOI22_X1 port map( A1 => n61558, A2 => n16842, B1 => n61553, B2 => 
                           n16843, ZN => n8182);
   U9959 : AOI22_X1 port map( A1 => n61546, A2 => n4266, B1 => n61541, B2 => 
                           n4258, ZN => n8183);
   U9960 : AOI22_X1 port map( A1 => n61534, A2 => n16443, B1 => n61529, B2 => 
                           n16451, ZN => n8184);
   U9961 : AOI22_X1 port map( A1 => n61609, A2 => n121, B1 => n61604, B2 => 
                           n113, ZN => n8174);
   U9962 : AOI22_X1 port map( A1 => n61597, A2 => n15966, B1 => n61592, B2 => 
                           n15967, ZN => n8175);
   U9963 : AOI22_X1 port map( A1 => n61585, A2 => n3957, B1 => n61580, B2 => 
                           n3965, ZN => n8176);
   U9964 : AOI22_X1 port map( A1 => n61495, A2 => n524, B1 => n61490, B2 => 
                           n532, ZN => n8191);
   U9965 : AOI22_X1 port map( A1 => n61483, A2 => n507, B1 => n61478, B2 => 
                           n515, ZN => n8192);
   U9966 : AOI22_X1 port map( A1 => n61660, A2 => n4173, B1 => n61655, B2 => 
                           n4165, ZN => n8166);
   U9967 : AOI22_X1 port map( A1 => n61648, A2 => n51625, B1 => n61643, B2 => 
                           n51649, ZN => n8167);
   U9968 : AOI22_X1 port map( A1 => n61636, A2 => n51617, B1 => n61631, B2 => 
                           n51609, ZN => n8168);
   U9969 : AOI22_X1 port map( A1 => n61354, A2 => n381, B1 => n61349, B2 => 
                           n373, ZN => n8218);
   U9970 : AOI22_X1 port map( A1 => n61342, A2 => n15322, B1 => n61337, B2 => 
                           n15330, ZN => n8219);
   U9971 : AOI22_X1 port map( A1 => n61330, A2 => n349, B1 => n61325, B2 => 
                           n341, ZN => n8220);
   U9972 : AOI22_X1 port map( A1 => n61381, A2 => n50965, B1 => n61376, B2 => 
                           n50933, ZN => n8212);
   U9973 : AOI22_X1 port map( A1 => n61405, A2 => n51713, B1 => n61400, B2 => 
                           n51721, ZN => n8210);
   U9974 : AOI22_X1 port map( A1 => n61393, A2 => n15473, B1 => n61388, B2 => 
                           n15481, ZN => n8211);
   U9975 : AOI22_X1 port map( A1 => n61291, A2 => n4290, B1 => n61286, B2 => 
                           n4298, ZN => n8227);
   U9976 : AOI22_X1 port map( A1 => n61279, A2 => n16475, B1 => n61274, B2 => 
                           n15669, ZN => n8228);
   U9977 : AOI22_X1 port map( A1 => n61456, A2 => n51761, B1 => n61451, B2 => 
                           n51769, ZN => n8202);
   U9978 : AOI22_X1 port map( A1 => n61444, A2 => n445, B1 => n61439, B2 => 
                           n437, ZN => n8203);
   U9979 : AOI22_X1 port map( A1 => n61432, A2 => n51729, B1 => n61427, B2 => 
                           n51737, ZN => n8204);
   U9980 : AOI22_X1 port map( A1 => n61558, A2 => n16844, B1 => n61553, B2 => 
                           n16845, ZN => n8007);
   U9981 : AOI22_X1 port map( A1 => n61546, A2 => n4265, B1 => n61541, B2 => 
                           n4257, ZN => n8012);
   U9982 : AOI22_X1 port map( A1 => n61534, A2 => n16444, B1 => n61529, B2 => 
                           n16452, ZN => n8017);
   U9983 : AOI22_X1 port map( A1 => n61609, A2 => n120, B1 => n61604, B2 => 
                           n112, ZN => n7982);
   U9984 : AOI22_X1 port map( A1 => n61597, A2 => n15970, B1 => n61592, B2 => 
                           n15971, ZN => n7987);
   U9985 : AOI22_X1 port map( A1 => n61585, A2 => n3956, B1 => n61580, B2 => 
                           n3964, ZN => n7992);
   U9986 : AOI22_X1 port map( A1 => n61495, A2 => n523, B1 => n61490, B2 => 
                           n531, ZN => n8037);
   U9987 : AOI22_X1 port map( A1 => n61483, A2 => n506, B1 => n61478, B2 => 
                           n514, ZN => n8042);
   U9988 : AOI22_X1 port map( A1 => n61660, A2 => n4172, B1 => n61655, B2 => 
                           n4164, ZN => n7957);
   U9989 : AOI22_X1 port map( A1 => n61648, A2 => n51624, B1 => n61643, B2 => 
                           n51648, ZN => n7962);
   U9990 : AOI22_X1 port map( A1 => n61636, A2 => n51616, B1 => n61631, B2 => 
                           n51608, ZN => n7967);
   U9991 : AOI22_X1 port map( A1 => n61354, A2 => n380, B1 => n61349, B2 => 
                           n372, ZN => n8111);
   U9992 : AOI22_X1 port map( A1 => n61342, A2 => n15323, B1 => n61337, B2 => 
                           n15343, ZN => n8116);
   U9993 : AOI22_X1 port map( A1 => n61330, A2 => n348, B1 => n61325, B2 => 
                           n340, ZN => n8121);
   U9994 : AOI22_X1 port map( A1 => n61381, A2 => n50964, B1 => n61376, B2 => 
                           n50932, ZN => n8096);
   U9995 : AOI22_X1 port map( A1 => n61405, A2 => n51712, B1 => n61400, B2 => 
                           n51720, ZN => n8086);
   U9996 : AOI22_X1 port map( A1 => n61393, A2 => n15474, B1 => n61388, B2 => 
                           n15482, ZN => n8091);
   U9997 : AOI22_X1 port map( A1 => n61291, A2 => n4289, B1 => n61286, B2 => 
                           n4297, ZN => n8141);
   U9998 : AOI22_X1 port map( A1 => n61279, A2 => n16476, B1 => n61274, B2 => 
                           n15672, ZN => n8146);
   U9999 : AOI22_X1 port map( A1 => n61456, A2 => n51760, B1 => n61451, B2 => 
                           n51768, ZN => n8061);
   U10000 : AOI22_X1 port map( A1 => n61444, A2 => n444, B1 => n61439, B2 => 
                           n436, ZN => n8066);
   U10001 : AOI22_X1 port map( A1 => n61432, A2 => n51728, B1 => n61427, B2 => 
                           n51736, ZN => n8071);
   U10002 : AOI22_X1 port map( A1 => n61556, A2 => n16636, B1 => n61555, B2 => 
                           n16482, ZN => n15010);
   U10003 : AOI22_X1 port map( A1 => n61532, A2 => n16660, B1 => n61531, B2 => 
                           n16506, ZN => n15014);
   U10004 : AOI22_X1 port map( A1 => n61607, A2 => n1786, B1 => n61606, B2 => 
                           n1762, ZN => n14998);
   U10005 : AOI22_X1 port map( A1 => n61595, A2 => n15879, B1 => n61594, B2 => 
                           n15880, ZN => n14999);
   U10006 : AOI22_X1 port map( A1 => n61583, A2 => n4355, B1 => n61582, B2 => 
                           n4378, ZN => n15002);
   U10007 : AOI22_X1 port map( A1 => n61493, A2 => n663, B1 => n61492, B2 => 
                           n687, ZN => n15022);
   U10008 : AOI22_X1 port map( A1 => n61481, A2 => n615, B1 => n61480, B2 => 
                           n639, ZN => n15024);
   U10009 : AOI22_X1 port map( A1 => n61658, A2 => n971, B1 => n61657, B2 => 
                           n4698, ZN => n14976);
   U10010 : AOI22_X1 port map( A1 => n61634, A2 => n53499, B1 => n61633, B2 => 
                           n4575, ZN => n14989);
   U10011 : AOI22_X1 port map( A1 => n61352, A2 => n3026, B1 => n61351, B2 => 
                           n3002, ZN => n15056);
   U10012 : AOI22_X1 port map( A1 => n61340, A2 => n15380, B1 => n61339, B2 => 
                           n15402, ZN => n15059);
   U10013 : AOI22_X1 port map( A1 => n61328, A2 => n2486, B1 => n61327, B2 => 
                           n2462, ZN => n15060);
   U10014 : AOI22_X1 port map( A1 => n61379, A2 => n16140, B1 => n61378, B2 => 
                           n16477, ZN => n15049);
   U10015 : AOI22_X1 port map( A1 => n61403, A2 => n15878, B1 => n61402, B2 => 
                           n16530, ZN => n15046);
   U10016 : AOI22_X1 port map( A1 => n61391, A2 => n59665, B1 => n61390, B2 => 
                           n59710, ZN => n15048);
   U10017 : AOI22_X1 port map( A1 => n61289, A2 => n2318, B1 => n61288, B2 => 
                           n2342, ZN => n15069);
   U10018 : AOI22_X1 port map( A1 => n61277, A2 => n15464, B1 => n61276, B2 => 
                           n15440, ZN => n15070);
   U10019 : AOI22_X1 port map( A1 => n61454, A2 => n54347, B1 => n61453, B2 => 
                           n54371, ZN => n15035);
   U10020 : AOI22_X1 port map( A1 => n61442, A2 => n54495, B1 => n61441, B2 => 
                           n54639, ZN => n15037);
   U10021 : AOI22_X1 port map( A1 => n61430, A2 => n54251, B1 => n61429, B2 => 
                           n54275, ZN => n15039);
   U10022 : AOI22_X1 port map( A1 => n61556, A2 => n16637, B1 => n61555, B2 => 
                           n16483, ZN => n14917);
   U10023 : AOI22_X1 port map( A1 => n61532, A2 => n16661, B1 => n61531, B2 => 
                           n16507, ZN => n14919);
   U10024 : AOI22_X1 port map( A1 => n61607, A2 => n1785, B1 => n61606, B2 => 
                           n1761, ZN => n14909);
   U10025 : AOI22_X1 port map( A1 => n61595, A2 => n15884, B1 => n61594, B2 => 
                           n15885, ZN => n14910);
   U10026 : AOI22_X1 port map( A1 => n61583, A2 => n4354, B1 => n61582, B2 => 
                           n4377, ZN => n14911);
   U10027 : AOI22_X1 port map( A1 => n61493, A2 => n662, B1 => n61492, B2 => 
                           n686, ZN => n14926);
   U10028 : AOI22_X1 port map( A1 => n61481, A2 => n614, B1 => n61480, B2 => 
                           n638, ZN => n14927);
   U10029 : AOI22_X1 port map( A1 => n61658, A2 => n970, B1 => n61657, B2 => 
                           n4697, ZN => n14901);
   U10030 : AOI22_X1 port map( A1 => n61634, A2 => n53498, B1 => n61633, B2 => 
                           n4574, ZN => n14903);
   U10031 : AOI22_X1 port map( A1 => n61352, A2 => n3025, B1 => n61351, B2 => 
                           n3001, ZN => n14953);
   U10032 : AOI22_X1 port map( A1 => n61340, A2 => n15381, B1 => n61339, B2 => 
                           n15427, ZN => n14954);
   U10033 : AOI22_X1 port map( A1 => n61328, A2 => n2485, B1 => n61327, B2 => 
                           n2461, ZN => n14955);
   U10034 : AOI22_X1 port map( A1 => n61379, A2 => n16141, B1 => n61378, B2 => 
                           n16478, ZN => n14947);
   U10035 : AOI22_X1 port map( A1 => n61403, A2 => n15883, B1 => n61402, B2 => 
                           n16531, ZN => n14945);
   U10036 : AOI22_X1 port map( A1 => n61391, A2 => n59666, B1 => n61390, B2 => 
                           n59711, ZN => n14946);
   U10037 : AOI22_X1 port map( A1 => n61289, A2 => n2317, B1 => n61288, B2 => 
                           n2341, ZN => n14962);
   U10038 : AOI22_X1 port map( A1 => n61277, A2 => n15465, B1 => n61276, B2 => 
                           n15441, ZN => n14963);
   U10039 : AOI22_X1 port map( A1 => n61454, A2 => n54346, B1 => n61453, B2 => 
                           n54370, ZN => n14937);
   U10040 : AOI22_X1 port map( A1 => n61442, A2 => n54496, B1 => n61441, B2 => 
                           n54640, ZN => n14938);
   U10041 : AOI22_X1 port map( A1 => n61430, A2 => n54250, B1 => n61429, B2 => 
                           n54274, ZN => n14939);
   U10042 : AOI22_X1 port map( A1 => n61556, A2 => n16638, B1 => n61555, B2 => 
                           n16484, ZN => n14842);
   U10043 : AOI22_X1 port map( A1 => n61532, A2 => n16662, B1 => n61531, B2 => 
                           n16508, ZN => n14844);
   U10044 : AOI22_X1 port map( A1 => n61607, A2 => n1784, B1 => n61606, B2 => 
                           n1760, ZN => n14834);
   U10045 : AOI22_X1 port map( A1 => n61595, A2 => n15914, B1 => n61594, B2 => 
                           n15915, ZN => n14835);
   U10046 : AOI22_X1 port map( A1 => n61583, A2 => n4353, B1 => n61582, B2 => 
                           n4376, ZN => n14836);
   U10047 : AOI22_X1 port map( A1 => n61493, A2 => n661, B1 => n61492, B2 => 
                           n685, ZN => n14851);
   U10048 : AOI22_X1 port map( A1 => n61481, A2 => n613, B1 => n61480, B2 => 
                           n637, ZN => n14852);
   U10049 : AOI22_X1 port map( A1 => n61658, A2 => n969, B1 => n61657, B2 => 
                           n4696, ZN => n14826);
   U10050 : AOI22_X1 port map( A1 => n61634, A2 => n53497, B1 => n61633, B2 => 
                           n4573, ZN => n14828);
   U10051 : AOI22_X1 port map( A1 => n61352, A2 => n3024, B1 => n61351, B2 => 
                           n3000, ZN => n14878);
   U10052 : AOI22_X1 port map( A1 => n61340, A2 => n15382, B1 => n61339, B2 => 
                           n15428, ZN => n14879);
   U10053 : AOI22_X1 port map( A1 => n61328, A2 => n2484, B1 => n61327, B2 => 
                           n2460, ZN => n14880);
   U10054 : AOI22_X1 port map( A1 => n61379, A2 => n16142, B1 => n61378, B2 => 
                           n16479, ZN => n14872);
   U10055 : AOI22_X1 port map( A1 => n61403, A2 => n15888, B1 => n61402, B2 => 
                           n16532, ZN => n14870);
   U10056 : AOI22_X1 port map( A1 => n61391, A2 => n59667, B1 => n61390, B2 => 
                           n59712, ZN => n14871);
   U10057 : AOI22_X1 port map( A1 => n61289, A2 => n2316, B1 => n61288, B2 => 
                           n2340, ZN => n14887);
   U10058 : AOI22_X1 port map( A1 => n61277, A2 => n15466, B1 => n61276, B2 => 
                           n15442, ZN => n14888);
   U10059 : AOI22_X1 port map( A1 => n61454, A2 => n54345, B1 => n61453, B2 => 
                           n54369, ZN => n14862);
   U10060 : AOI22_X1 port map( A1 => n61442, A2 => n54497, B1 => n61441, B2 => 
                           n54641, ZN => n14863);
   U10061 : AOI22_X1 port map( A1 => n61430, A2 => n54249, B1 => n61429, B2 => 
                           n54273, ZN => n14864);
   U10062 : AOI22_X1 port map( A1 => n61556, A2 => n16639, B1 => n61555, B2 => 
                           n16485, ZN => n14767);
   U10063 : AOI22_X1 port map( A1 => n61532, A2 => n16663, B1 => n61531, B2 => 
                           n16509, ZN => n14769);
   U10064 : AOI22_X1 port map( A1 => n61607, A2 => n1783, B1 => n61606, B2 => 
                           n1759, ZN => n14759);
   U10065 : AOI22_X1 port map( A1 => n61595, A2 => n15892, B1 => n61594, B2 => 
                           n15893, ZN => n14760);
   U10066 : AOI22_X1 port map( A1 => n61583, A2 => n4352, B1 => n61582, B2 => 
                           n4375, ZN => n14761);
   U10067 : AOI22_X1 port map( A1 => n61493, A2 => n660, B1 => n61492, B2 => 
                           n684, ZN => n14776);
   U10068 : AOI22_X1 port map( A1 => n61481, A2 => n612, B1 => n61480, B2 => 
                           n636, ZN => n14777);
   U10069 : AOI22_X1 port map( A1 => n61658, A2 => n968, B1 => n61657, B2 => 
                           n956, ZN => n14751);
   U10070 : AOI22_X1 port map( A1 => n61634, A2 => n53496, B1 => n61633, B2 => 
                           n4572, ZN => n14753);
   U10071 : AOI22_X1 port map( A1 => n61352, A2 => n3023, B1 => n61351, B2 => 
                           n2999, ZN => n14803);
   U10072 : AOI22_X1 port map( A1 => n61340, A2 => n15383, B1 => n61339, B2 => 
                           n15429, ZN => n14804);
   U10073 : AOI22_X1 port map( A1 => n61328, A2 => n2483, B1 => n61327, B2 => 
                           n2459, ZN => n14805);
   U10074 : AOI22_X1 port map( A1 => n61379, A2 => n16138, B1 => n61378, B2 => 
                           n16480, ZN => n14797);
   U10075 : AOI22_X1 port map( A1 => n61403, A2 => n15891, B1 => n61402, B2 => 
                           n16533, ZN => n14795);
   U10076 : AOI22_X1 port map( A1 => n61391, A2 => n59668, B1 => n61390, B2 => 
                           n59713, ZN => n14796);
   U10077 : AOI22_X1 port map( A1 => n61289, A2 => n2315, B1 => n61288, B2 => 
                           n2339, ZN => n14812);
   U10078 : AOI22_X1 port map( A1 => n61277, A2 => n15499, B1 => n61276, B2 => 
                           n15443, ZN => n14813);
   U10079 : AOI22_X1 port map( A1 => n61454, A2 => n54344, B1 => n61453, B2 => 
                           n54368, ZN => n14787);
   U10080 : AOI22_X1 port map( A1 => n61442, A2 => n54498, B1 => n61441, B2 => 
                           n54642, ZN => n14788);
   U10081 : AOI22_X1 port map( A1 => n61430, A2 => n54248, B1 => n61429, B2 => 
                           n54272, ZN => n14789);
   U10082 : AOI22_X1 port map( A1 => n61556, A2 => n16640, B1 => n61555, B2 => 
                           n16486, ZN => n14692);
   U10083 : AOI22_X1 port map( A1 => n61532, A2 => n16664, B1 => n61531, B2 => 
                           n16510, ZN => n14694);
   U10084 : AOI22_X1 port map( A1 => n61607, A2 => n1782, B1 => n61606, B2 => 
                           n1758, ZN => n14684);
   U10085 : AOI22_X1 port map( A1 => n61595, A2 => n15897, B1 => n61594, B2 => 
                           n15898, ZN => n14685);
   U10086 : AOI22_X1 port map( A1 => n61583, A2 => n4351, B1 => n61582, B2 => 
                           n519, ZN => n14686);
   U10087 : AOI22_X1 port map( A1 => n61493, A2 => n659, B1 => n61492, B2 => 
                           n683, ZN => n14701);
   U10088 : AOI22_X1 port map( A1 => n61481, A2 => n611, B1 => n61480, B2 => 
                           n635, ZN => n14702);
   U10089 : AOI22_X1 port map( A1 => n61658, A2 => n967, B1 => n61657, B2 => 
                           n955, ZN => n14676);
   U10090 : AOI22_X1 port map( A1 => n61634, A2 => n53495, B1 => n61633, B2 => 
                           n4571, ZN => n14678);
   U10091 : AOI22_X1 port map( A1 => n61352, A2 => n3022, B1 => n61351, B2 => 
                           n2998, ZN => n14728);
   U10092 : AOI22_X1 port map( A1 => n61340, A2 => n15384, B1 => n61339, B2 => 
                           n15430, ZN => n14729);
   U10093 : AOI22_X1 port map( A1 => n61328, A2 => n2906, B1 => n61327, B2 => 
                           n2458, ZN => n14730);
   U10094 : AOI22_X1 port map( A1 => n61379, A2 => n16139, B1 => n61378, B2 => 
                           n16481, ZN => n14722);
   U10095 : AOI22_X1 port map( A1 => n61403, A2 => n15896, B1 => n61402, B2 => 
                           n16534, ZN => n14720);
   U10096 : AOI22_X1 port map( A1 => n61391, A2 => n59669, B1 => n61390, B2 => 
                           n59714, ZN => n14721);
   U10097 : AOI22_X1 port map( A1 => n61289, A2 => n2314, B1 => n61288, B2 => 
                           n2338, ZN => n14737);
   U10098 : AOI22_X1 port map( A1 => n61277, A2 => n15500, B1 => n61276, B2 => 
                           n15444, ZN => n14738);
   U10099 : AOI22_X1 port map( A1 => n61454, A2 => n54343, B1 => n61453, B2 => 
                           n54367, ZN => n14712);
   U10100 : AOI22_X1 port map( A1 => n61442, A2 => n54499, B1 => n61441, B2 => 
                           n54643, ZN => n14713);
   U10101 : AOI22_X1 port map( A1 => n61430, A2 => n54247, B1 => n61429, B2 => 
                           n54271, ZN => n14714);
   U10102 : AOI22_X1 port map( A1 => n61556, A2 => n16641, B1 => n61555, B2 => 
                           n16487, ZN => n14617);
   U10103 : AOI22_X1 port map( A1 => n61532, A2 => n16665, B1 => n61531, B2 => 
                           n16511, ZN => n14619);
   U10104 : AOI22_X1 port map( A1 => n61607, A2 => n1781, B1 => n61606, B2 => 
                           n1757, ZN => n14609);
   U10105 : AOI22_X1 port map( A1 => n61595, A2 => n15902, B1 => n61594, B2 => 
                           n15903, ZN => n14610);
   U10106 : AOI22_X1 port map( A1 => n61583, A2 => n4350, B1 => n61582, B2 => 
                           n4374, ZN => n14611);
   U10107 : AOI22_X1 port map( A1 => n61493, A2 => n658, B1 => n61492, B2 => 
                           n682, ZN => n14626);
   U10108 : AOI22_X1 port map( A1 => n61481, A2 => n610, B1 => n61480, B2 => 
                           n634, ZN => n14627);
   U10109 : AOI22_X1 port map( A1 => n61658, A2 => n966, B1 => n61657, B2 => 
                           n954, ZN => n14601);
   U10110 : AOI22_X1 port map( A1 => n61634, A2 => n53494, B1 => n61633, B2 => 
                           n4570, ZN => n14603);
   U10111 : AOI22_X1 port map( A1 => n61352, A2 => n3021, B1 => n61351, B2 => 
                           n2997, ZN => n14653);
   U10112 : AOI22_X1 port map( A1 => n61340, A2 => n15385, B1 => n61339, B2 => 
                           n15431, ZN => n14654);
   U10113 : AOI22_X1 port map( A1 => n61328, A2 => n2905, B1 => n61327, B2 => 
                           n2457, ZN => n14655);
   U10114 : AOI22_X1 port map( A1 => n61379, A2 => n16124, B1 => n61378, B2 => 
                           n16125, ZN => n14647);
   U10115 : AOI22_X1 port map( A1 => n61403, A2 => n15901, B1 => n61402, B2 => 
                           n16535, ZN => n14645);
   U10116 : AOI22_X1 port map( A1 => n61391, A2 => n59670, B1 => n61390, B2 => 
                           n59715, ZN => n14646);
   U10117 : AOI22_X1 port map( A1 => n61289, A2 => n2313, B1 => n61288, B2 => 
                           n2337, ZN => n14662);
   U10118 : AOI22_X1 port map( A1 => n61277, A2 => n15501, B1 => n61276, B2 => 
                           n15445, ZN => n14663);
   U10119 : AOI22_X1 port map( A1 => n61454, A2 => n54342, B1 => n61453, B2 => 
                           n54366, ZN => n14637);
   U10120 : AOI22_X1 port map( A1 => n61442, A2 => n54500, B1 => n61441, B2 => 
                           n54644, ZN => n14638);
   U10121 : AOI22_X1 port map( A1 => n61430, A2 => n54246, B1 => n61429, B2 => 
                           n54270, ZN => n14639);
   U10122 : AOI22_X1 port map( A1 => n61556, A2 => n16642, B1 => n61555, B2 => 
                           n16488, ZN => n14542);
   U10123 : AOI22_X1 port map( A1 => n61532, A2 => n16666, B1 => n61531, B2 => 
                           n16512, ZN => n14544);
   U10124 : AOI22_X1 port map( A1 => n61607, A2 => n1780, B1 => n61606, B2 => 
                           n1756, ZN => n14534);
   U10125 : AOI22_X1 port map( A1 => n61595, A2 => n15907, B1 => n61594, B2 => 
                           n15908, ZN => n14535);
   U10126 : AOI22_X1 port map( A1 => n61583, A2 => n4349, B1 => n61582, B2 => 
                           n4373, ZN => n14536);
   U10127 : AOI22_X1 port map( A1 => n61493, A2 => n657, B1 => n61492, B2 => 
                           n681, ZN => n14551);
   U10128 : AOI22_X1 port map( A1 => n61481, A2 => n609, B1 => n61480, B2 => 
                           n633, ZN => n14552);
   U10129 : AOI22_X1 port map( A1 => n61658, A2 => n965, B1 => n61657, B2 => 
                           n953, ZN => n14526);
   U10130 : AOI22_X1 port map( A1 => n61634, A2 => n53493, B1 => n61633, B2 => 
                           n4569, ZN => n14528);
   U10131 : AOI22_X1 port map( A1 => n61352, A2 => n3020, B1 => n61351, B2 => 
                           n2996, ZN => n14578);
   U10132 : AOI22_X1 port map( A1 => n61340, A2 => n15726, B1 => n61339, B2 => 
                           n16554, ZN => n14579);
   U10133 : AOI22_X1 port map( A1 => n61328, A2 => n2904, B1 => n61327, B2 => 
                           n2456, ZN => n14580);
   U10134 : AOI22_X1 port map( A1 => n61379, A2 => n16126, B1 => n61378, B2 => 
                           n16127, ZN => n14572);
   U10135 : AOI22_X1 port map( A1 => n61403, A2 => n15906, B1 => n61402, B2 => 
                           n16536, ZN => n14570);
   U10136 : AOI22_X1 port map( A1 => n61391, A2 => n59671, B1 => n61390, B2 => 
                           n59716, ZN => n14571);
   U10137 : AOI22_X1 port map( A1 => n61289, A2 => n2312, B1 => n61288, B2 => 
                           n2336, ZN => n14587);
   U10138 : AOI22_X1 port map( A1 => n61277, A2 => n15502, B1 => n61276, B2 => 
                           n15446, ZN => n14588);
   U10139 : AOI22_X1 port map( A1 => n61454, A2 => n54341, B1 => n61453, B2 => 
                           n54365, ZN => n14562);
   U10140 : AOI22_X1 port map( A1 => n61442, A2 => n54501, B1 => n61441, B2 => 
                           n54645, ZN => n14563);
   U10141 : AOI22_X1 port map( A1 => n61430, A2 => n54245, B1 => n61429, B2 => 
                           n54269, ZN => n14564);
   U10142 : AOI22_X1 port map( A1 => n61556, A2 => n16643, B1 => n61555, B2 => 
                           n16489, ZN => n14467);
   U10143 : AOI22_X1 port map( A1 => n61532, A2 => n16667, B1 => n61531, B2 => 
                           n16513, ZN => n14469);
   U10144 : AOI22_X1 port map( A1 => n61607, A2 => n1779, B1 => n61606, B2 => 
                           n1755, ZN => n14459);
   U10145 : AOI22_X1 port map( A1 => n61595, A2 => n15912, B1 => n61594, B2 => 
                           n15913, ZN => n14460);
   U10146 : AOI22_X1 port map( A1 => n61583, A2 => n4348, B1 => n61582, B2 => 
                           n4372, ZN => n14461);
   U10147 : AOI22_X1 port map( A1 => n61493, A2 => n656, B1 => n61492, B2 => 
                           n680, ZN => n14476);
   U10148 : AOI22_X1 port map( A1 => n61481, A2 => n608, B1 => n61480, B2 => 
                           n632, ZN => n14477);
   U10149 : AOI22_X1 port map( A1 => n61658, A2 => n964, B1 => n61657, B2 => 
                           n952, ZN => n14451);
   U10150 : AOI22_X1 port map( A1 => n61634, A2 => n53492, B1 => n61633, B2 => 
                           n4568, ZN => n14453);
   U10151 : AOI22_X1 port map( A1 => n61352, A2 => n3019, B1 => n61351, B2 => 
                           n2995, ZN => n14503);
   U10152 : AOI22_X1 port map( A1 => n61340, A2 => n15729, B1 => n61339, B2 => 
                           n16555, ZN => n14504);
   U10153 : AOI22_X1 port map( A1 => n61328, A2 => n2903, B1 => n61327, B2 => 
                           n2455, ZN => n14505);
   U10154 : AOI22_X1 port map( A1 => n61379, A2 => n16130, B1 => n61378, B2 => 
                           n16131, ZN => n14497);
   U10155 : AOI22_X1 port map( A1 => n61403, A2 => n15911, B1 => n61402, B2 => 
                           n16537, ZN => n14495);
   U10156 : AOI22_X1 port map( A1 => n61391, A2 => n59672, B1 => n61390, B2 => 
                           n59717, ZN => n14496);
   U10157 : AOI22_X1 port map( A1 => n61289, A2 => n2311, B1 => n61288, B2 => 
                           n2335, ZN => n14512);
   U10158 : AOI22_X1 port map( A1 => n61277, A2 => n15503, B1 => n61276, B2 => 
                           n15447, ZN => n14513);
   U10159 : AOI22_X1 port map( A1 => n61454, A2 => n54340, B1 => n61453, B2 => 
                           n54364, ZN => n14487);
   U10160 : AOI22_X1 port map( A1 => n61442, A2 => n54502, B1 => n61441, B2 => 
                           n54646, ZN => n14488);
   U10161 : AOI22_X1 port map( A1 => n61430, A2 => n54244, B1 => n61429, B2 => 
                           n54268, ZN => n14489);
   U10162 : AOI22_X1 port map( A1 => n16672, A2 => n61883, B1 => n16518, B2 => 
                           n61880, ZN => n6965);
   U10163 : AOI22_X1 port map( A1 => n15839, A2 => n61895, B1 => n15815, B2 => 
                           n61892, ZN => n6964);
   U10164 : AOI22_X1 port map( A1 => n699, A2 => n62168, B1 => n723, B2 => 
                           n62166, ZN => n6973);
   U10165 : AOI22_X1 port map( A1 => n16306, A2 => n61874, B1 => n16696, B2 => 
                           n61871, ZN => n6972);
   U10166 : AOI22_X1 port map( A1 => n16624, A2 => n61928, B1 => n16600, B2 => 
                           n61925, ZN => n6956);
   U10167 : AOI22_X1 port map( A1 => n15771, A2 => n61916, B1 => n15772, B2 => 
                           n61913, ZN => n6957);
   U10168 : AOI22_X1 port map( A1 => n2898, A2 => n61793, B1 => n2450, B2 => 
                           n61790, ZN => n6947);
   U10169 : AOI22_X1 port map( A1 => n53487, A2 => n61943, B1 => n61940, B2 => 
                           n4563, ZN => n6949);
   U10170 : AOI22_X1 port map( A1 => n54215, A2 => n62134, B1 => n54167, B2 => 
                           n62132, ZN => n6992);
   U10171 : AOI22_X1 port map( A1 => n15769, A2 => n62138, B1 => n15768, B2 => 
                           n62136, ZN => n6993);
   U10172 : AOI22_X1 port map( A1 => n16542, A2 => n61832, B1 => n15770, B2 => 
                           n61829, ZN => n6991);
   U10173 : AOI22_X1 port map( A1 => n54359, A2 => n61853, B1 => n54335, B2 => 
                           n61850, ZN => n6984);
   U10174 : AOI22_X1 port map( A1 => n54483, A2 => n61841, B1 => n54627, B2 => 
                           n61838, ZN => n6985);
   U10175 : AOI22_X1 port map( A1 => n52171, A2 => n61766, B1 => n52195, B2 => 
                           n61763, ZN => n7008);
   U10176 : AOI22_X1 port map( A1 => n15508, A2 => n61754, B1 => n15452, B2 => 
                           n61751, ZN => n7009);
   U10177 : AOI22_X1 port map( A1 => n53927, A2 => n61811, B1 => n53975, B2 => 
                           n61808, ZN => n6999);
   U10178 : AOI22_X1 port map( A1 => n3014, A2 => n61805, B1 => n2990, B2 => 
                           n61802, ZN => n7000);
   U10179 : OAI22_X1 port map( A1 => n60795, A2 => n61966, B1 => n52979, B2 => 
                           n60794, ZN => n13733);
   U10180 : OAI22_X1 port map( A1 => n60795, A2 => n61980, B1 => n52978, B2 => 
                           n60794, ZN => n13734);
   U10181 : OAI22_X1 port map( A1 => n60795, A2 => n61994, B1 => n52977, B2 => 
                           n60794, ZN => n13735);
   U10182 : OAI22_X1 port map( A1 => n60795, A2 => n62008, B1 => n52976, B2 => 
                           n60794, ZN => n13736);
   U10183 : OAI22_X1 port map( A1 => n60795, A2 => n62022, B1 => n52975, B2 => 
                           n60794, ZN => n13737);
   U10184 : OAI22_X1 port map( A1 => n60796, A2 => n62036, B1 => n52974, B2 => 
                           n60794, ZN => n13738);
   U10185 : OAI22_X1 port map( A1 => n60796, A2 => n62050, B1 => n52973, B2 => 
                           n60794, ZN => n13739);
   U10186 : OAI22_X1 port map( A1 => n60796, A2 => n62064, B1 => n52972, B2 => 
                           n60794, ZN => n13740);
   U10187 : OAI22_X1 port map( A1 => n60796, A2 => n62078, B1 => n52971, B2 => 
                           n60794, ZN => n13741);
   U10188 : OAI22_X1 port map( A1 => n60796, A2 => n62092, B1 => n52970, B2 => 
                           n60794, ZN => n13742);
   U10189 : OAI22_X1 port map( A1 => n60797, A2 => n62106, B1 => n52969, B2 => 
                           n60794, ZN => n13743);
   U10190 : OAI22_X1 port map( A1 => n60797, A2 => n60959, B1 => n52968, B2 => 
                           n60794, ZN => n13744);
   U10191 : OAI22_X1 port map( A1 => n60797, A2 => n60973, B1 => n52967, B2 => 
                           n15131, ZN => n13745);
   U10192 : OAI22_X1 port map( A1 => n60797, A2 => n60987, B1 => n52966, B2 => 
                           n15131, ZN => n13746);
   U10193 : OAI22_X1 port map( A1 => n60797, A2 => n61001, B1 => n52965, B2 => 
                           n15131, ZN => n13747);
   U10194 : OAI22_X1 port map( A1 => n60798, A2 => n61015, B1 => n52964, B2 => 
                           n15131, ZN => n13748);
   U10195 : OAI22_X1 port map( A1 => n60798, A2 => n61029, B1 => n52963, B2 => 
                           n15131, ZN => n13749);
   U10196 : OAI22_X1 port map( A1 => n60798, A2 => n61043, B1 => n52962, B2 => 
                           n15131, ZN => n13750);
   U10197 : OAI22_X1 port map( A1 => n60798, A2 => n61057, B1 => n52961, B2 => 
                           n15131, ZN => n13751);
   U10198 : OAI22_X1 port map( A1 => n60798, A2 => n61071, B1 => n52960, B2 => 
                           n60794, ZN => n13752);
   U10199 : OAI22_X1 port map( A1 => n60799, A2 => n61085, B1 => n52959, B2 => 
                           n60794, ZN => n13753);
   U10200 : OAI22_X1 port map( A1 => n60799, A2 => n61099, B1 => n52958, B2 => 
                           n60794, ZN => n13754);
   U10201 : OAI22_X1 port map( A1 => n60799, A2 => n61113, B1 => n52957, B2 => 
                           n60794, ZN => n13755);
   U10202 : OAI22_X1 port map( A1 => n60799, A2 => n61127, B1 => n52956, B2 => 
                           n60794, ZN => n13756);
   U10203 : OAI22_X1 port map( A1 => n59976, A2 => n61974, B1 => n2510, B2 => 
                           n59975, ZN => n10821);
   U10204 : OAI22_X1 port map( A1 => n59976, A2 => n61988, B1 => n2509, B2 => 
                           n59975, ZN => n10822);
   U10205 : OAI22_X1 port map( A1 => n59976, A2 => n62002, B1 => n2508, B2 => 
                           n59975, ZN => n10823);
   U10206 : OAI22_X1 port map( A1 => n59976, A2 => n62016, B1 => n2507, B2 => 
                           n59975, ZN => n10824);
   U10207 : OAI22_X1 port map( A1 => n59976, A2 => n62030, B1 => n2506, B2 => 
                           n59975, ZN => n10825);
   U10208 : OAI22_X1 port map( A1 => n59977, A2 => n62044, B1 => n2505, B2 => 
                           n59975, ZN => n10826);
   U10209 : OAI22_X1 port map( A1 => n59977, A2 => n62058, B1 => n2504, B2 => 
                           n59975, ZN => n10827);
   U10210 : OAI22_X1 port map( A1 => n59977, A2 => n62072, B1 => n2503, B2 => 
                           n59975, ZN => n10828);
   U10211 : OAI22_X1 port map( A1 => n59977, A2 => n62086, B1 => n2502, B2 => 
                           n59975, ZN => n10829);
   U10212 : OAI22_X1 port map( A1 => n59977, A2 => n62100, B1 => n2501, B2 => 
                           n59975, ZN => n10830);
   U10213 : OAI22_X1 port map( A1 => n59978, A2 => n62114, B1 => n2500, B2 => 
                           n59975, ZN => n10831);
   U10214 : OAI22_X1 port map( A1 => n59978, A2 => n60967, B1 => n2499, B2 => 
                           n59975, ZN => n10832);
   U10215 : OAI22_X1 port map( A1 => n59978, A2 => n60981, B1 => n2498, B2 => 
                           n15243, ZN => n10833);
   U10216 : OAI22_X1 port map( A1 => n59978, A2 => n60995, B1 => n2497, B2 => 
                           n15243, ZN => n10834);
   U10217 : OAI22_X1 port map( A1 => n59978, A2 => n61009, B1 => n2496, B2 => 
                           n15243, ZN => n10835);
   U10218 : OAI22_X1 port map( A1 => n59979, A2 => n61023, B1 => n2495, B2 => 
                           n15243, ZN => n10836);
   U10219 : OAI22_X1 port map( A1 => n59979, A2 => n61037, B1 => n2494, B2 => 
                           n15243, ZN => n10837);
   U10220 : OAI22_X1 port map( A1 => n59979, A2 => n61051, B1 => n2493, B2 => 
                           n15243, ZN => n10838);
   U10221 : OAI22_X1 port map( A1 => n59979, A2 => n61065, B1 => n2492, B2 => 
                           n15243, ZN => n10839);
   U10222 : OAI22_X1 port map( A1 => n59979, A2 => n61079, B1 => n2491, B2 => 
                           n59975, ZN => n10840);
   U10223 : OAI22_X1 port map( A1 => n59980, A2 => n61093, B1 => n2490, B2 => 
                           n59975, ZN => n10841);
   U10224 : OAI22_X1 port map( A1 => n59980, A2 => n61107, B1 => n2489, B2 => 
                           n59975, ZN => n10842);
   U10225 : OAI22_X1 port map( A1 => n59980, A2 => n61121, B1 => n2488, B2 => 
                           n59975, ZN => n10843);
   U10226 : OAI22_X1 port map( A1 => n59980, A2 => n61135, B1 => n2487, B2 => 
                           n59975, ZN => n10844);
   U10227 : OAI22_X1 port map( A1 => n60948, A2 => n61965, B1 => n2076, B2 => 
                           n60947, ZN => n14277);
   U10228 : OAI22_X1 port map( A1 => n60948, A2 => n61979, B1 => n2248, B2 => 
                           n60947, ZN => n14278);
   U10229 : OAI22_X1 port map( A1 => n60948, A2 => n61993, B1 => n2247, B2 => 
                           n60947, ZN => n14279);
   U10230 : OAI22_X1 port map( A1 => n60948, A2 => n62007, B1 => n2246, B2 => 
                           n60947, ZN => n14280);
   U10231 : OAI22_X1 port map( A1 => n60948, A2 => n62021, B1 => n2245, B2 => 
                           n60947, ZN => n14281);
   U10232 : OAI22_X1 port map( A1 => n60949, A2 => n62035, B1 => n2244, B2 => 
                           n60947, ZN => n14282);
   U10233 : OAI22_X1 port map( A1 => n60949, A2 => n62049, B1 => n2243, B2 => 
                           n60947, ZN => n14283);
   U10234 : OAI22_X1 port map( A1 => n60949, A2 => n62063, B1 => n2242, B2 => 
                           n60947, ZN => n14284);
   U10235 : OAI22_X1 port map( A1 => n60949, A2 => n62077, B1 => n2241, B2 => 
                           n60947, ZN => n14285);
   U10236 : OAI22_X1 port map( A1 => n60949, A2 => n62091, B1 => n2240, B2 => 
                           n60947, ZN => n14286);
   U10237 : OAI22_X1 port map( A1 => n60950, A2 => n62105, B1 => n2239, B2 => 
                           n60947, ZN => n14287);
   U10238 : OAI22_X1 port map( A1 => n60950, A2 => n60958, B1 => n2075, B2 => 
                           n60947, ZN => n14288);
   U10239 : OAI22_X1 port map( A1 => n60950, A2 => n60972, B1 => n2238, B2 => 
                           n15096, ZN => n14289);
   U10240 : OAI22_X1 port map( A1 => n60950, A2 => n60986, B1 => n2237, B2 => 
                           n15096, ZN => n14290);
   U10241 : OAI22_X1 port map( A1 => n60950, A2 => n61000, B1 => n2236, B2 => 
                           n15096, ZN => n14291);
   U10242 : OAI22_X1 port map( A1 => n60951, A2 => n61014, B1 => n2235, B2 => 
                           n15096, ZN => n14292);
   U10243 : OAI22_X1 port map( A1 => n60951, A2 => n61028, B1 => n2220, B2 => 
                           n15096, ZN => n14293);
   U10244 : OAI22_X1 port map( A1 => n60951, A2 => n61042, B1 => n2219, B2 => 
                           n15096, ZN => n14294);
   U10245 : OAI22_X1 port map( A1 => n60951, A2 => n61056, B1 => n2218, B2 => 
                           n15096, ZN => n14295);
   U10246 : OAI22_X1 port map( A1 => n60951, A2 => n61070, B1 => n2217, B2 => 
                           n60947, ZN => n14296);
   U10247 : OAI22_X1 port map( A1 => n60952, A2 => n61084, B1 => n2216, B2 => 
                           n60947, ZN => n14297);
   U10248 : OAI22_X1 port map( A1 => n60952, A2 => n61098, B1 => n2215, B2 => 
                           n60947, ZN => n14298);
   U10249 : OAI22_X1 port map( A1 => n60952, A2 => n61112, B1 => n2214, B2 => 
                           n60947, ZN => n14299);
   U10250 : OAI22_X1 port map( A1 => n60952, A2 => n61126, B1 => n2213, B2 => 
                           n60947, ZN => n14300);
   U10251 : OAI22_X1 port map( A1 => n60516, A2 => n61969, B1 => n53171, B2 => 
                           n60515, ZN => n12741);
   U10252 : OAI22_X1 port map( A1 => n60516, A2 => n61983, B1 => n53170, B2 => 
                           n60515, ZN => n12742);
   U10253 : OAI22_X1 port map( A1 => n60516, A2 => n61997, B1 => n53169, B2 => 
                           n60515, ZN => n12743);
   U10254 : OAI22_X1 port map( A1 => n60516, A2 => n62011, B1 => n53168, B2 => 
                           n60515, ZN => n12744);
   U10255 : OAI22_X1 port map( A1 => n60516, A2 => n62025, B1 => n53167, B2 => 
                           n60515, ZN => n12745);
   U10256 : OAI22_X1 port map( A1 => n60517, A2 => n62039, B1 => n53166, B2 => 
                           n60515, ZN => n12746);
   U10257 : OAI22_X1 port map( A1 => n60517, A2 => n62053, B1 => n53165, B2 => 
                           n60515, ZN => n12747);
   U10258 : OAI22_X1 port map( A1 => n60517, A2 => n62067, B1 => n53164, B2 => 
                           n60515, ZN => n12748);
   U10259 : OAI22_X1 port map( A1 => n60517, A2 => n62081, B1 => n53163, B2 => 
                           n60515, ZN => n12749);
   U10260 : OAI22_X1 port map( A1 => n60517, A2 => n62095, B1 => n53162, B2 => 
                           n60515, ZN => n12750);
   U10261 : OAI22_X1 port map( A1 => n60518, A2 => n62109, B1 => n53161, B2 => 
                           n60515, ZN => n12751);
   U10262 : OAI22_X1 port map( A1 => n60518, A2 => n60962, B1 => n53160, B2 => 
                           n60515, ZN => n12752);
   U10263 : OAI22_X1 port map( A1 => n60518, A2 => n60976, B1 => n53159, B2 => 
                           n15165, ZN => n12753);
   U10264 : OAI22_X1 port map( A1 => n60518, A2 => n60990, B1 => n53158, B2 => 
                           n15165, ZN => n12754);
   U10265 : OAI22_X1 port map( A1 => n60518, A2 => n61004, B1 => n53157, B2 => 
                           n15165, ZN => n12755);
   U10266 : OAI22_X1 port map( A1 => n60519, A2 => n61018, B1 => n53156, B2 => 
                           n15165, ZN => n12756);
   U10267 : OAI22_X1 port map( A1 => n60519, A2 => n61032, B1 => n53155, B2 => 
                           n15165, ZN => n12757);
   U10268 : OAI22_X1 port map( A1 => n60519, A2 => n61046, B1 => n53154, B2 => 
                           n15165, ZN => n12758);
   U10269 : OAI22_X1 port map( A1 => n60519, A2 => n61060, B1 => n53153, B2 => 
                           n15165, ZN => n12759);
   U10270 : OAI22_X1 port map( A1 => n60519, A2 => n61074, B1 => n53152, B2 => 
                           n60515, ZN => n12760);
   U10271 : OAI22_X1 port map( A1 => n60520, A2 => n61088, B1 => n53151, B2 => 
                           n60515, ZN => n12761);
   U10272 : OAI22_X1 port map( A1 => n60520, A2 => n61102, B1 => n53150, B2 => 
                           n60515, ZN => n12762);
   U10273 : OAI22_X1 port map( A1 => n60520, A2 => n61116, B1 => n53149, B2 => 
                           n60515, ZN => n12763);
   U10274 : OAI22_X1 port map( A1 => n60520, A2 => n61130, B1 => n53148, B2 => 
                           n60515, ZN => n12764);
   U10275 : OAI22_X1 port map( A1 => n60940, A2 => n62091, B1 => n962, B2 => 
                           n60938, ZN => n14254);
   U10276 : OAI22_X1 port map( A1 => n60941, A2 => n62105, B1 => n961, B2 => 
                           n60938, ZN => n14255);
   U10277 : OAI22_X1 port map( A1 => n60941, A2 => n60958, B1 => n960, B2 => 
                           n60938, ZN => n14256);
   U10278 : OAI22_X1 port map( A1 => n60941, A2 => n60972, B1 => n959, B2 => 
                           n15098, ZN => n14257);
   U10279 : OAI22_X1 port map( A1 => n60941, A2 => n60986, B1 => n958, B2 => 
                           n15098, ZN => n14258);
   U10280 : OAI22_X1 port map( A1 => n60943, A2 => n61112, B1 => n957, B2 => 
                           n15098, ZN => n14267);
   U10281 : OAI22_X1 port map( A1 => n60831, A2 => n61966, B1 => n911, B2 => 
                           n60830, ZN => n13861);
   U10282 : OAI22_X1 port map( A1 => n60831, A2 => n61980, B1 => n910, B2 => 
                           n60830, ZN => n13862);
   U10283 : OAI22_X1 port map( A1 => n60831, A2 => n61994, B1 => n909, B2 => 
                           n60830, ZN => n13863);
   U10284 : OAI22_X1 port map( A1 => n60831, A2 => n62008, B1 => n908, B2 => 
                           n60830, ZN => n13864);
   U10285 : OAI22_X1 port map( A1 => n60831, A2 => n62022, B1 => n907, B2 => 
                           n60830, ZN => n13865);
   U10286 : OAI22_X1 port map( A1 => n60832, A2 => n62036, B1 => n906, B2 => 
                           n60830, ZN => n13866);
   U10287 : OAI22_X1 port map( A1 => n60832, A2 => n62050, B1 => n905, B2 => 
                           n60830, ZN => n13867);
   U10288 : OAI22_X1 port map( A1 => n60832, A2 => n62064, B1 => n904, B2 => 
                           n60830, ZN => n13868);
   U10289 : OAI22_X1 port map( A1 => n60832, A2 => n62078, B1 => n903, B2 => 
                           n60830, ZN => n13869);
   U10290 : OAI22_X1 port map( A1 => n60832, A2 => n62092, B1 => n902, B2 => 
                           n60830, ZN => n13870);
   U10291 : OAI22_X1 port map( A1 => n60833, A2 => n62106, B1 => n901, B2 => 
                           n60830, ZN => n13871);
   U10292 : OAI22_X1 port map( A1 => n60833, A2 => n60959, B1 => n900, B2 => 
                           n60830, ZN => n13872);
   U10293 : OAI22_X1 port map( A1 => n60833, A2 => n60973, B1 => n899, B2 => 
                           n15122, ZN => n13873);
   U10294 : OAI22_X1 port map( A1 => n60833, A2 => n60987, B1 => n898, B2 => 
                           n15122, ZN => n13874);
   U10295 : OAI22_X1 port map( A1 => n60833, A2 => n61001, B1 => n897, B2 => 
                           n15122, ZN => n13875);
   U10296 : OAI22_X1 port map( A1 => n60834, A2 => n61015, B1 => n896, B2 => 
                           n15122, ZN => n13876);
   U10297 : OAI22_X1 port map( A1 => n60834, A2 => n61029, B1 => n895, B2 => 
                           n15122, ZN => n13877);
   U10298 : OAI22_X1 port map( A1 => n60834, A2 => n61043, B1 => n894, B2 => 
                           n15122, ZN => n13878);
   U10299 : OAI22_X1 port map( A1 => n60834, A2 => n61057, B1 => n893, B2 => 
                           n15122, ZN => n13879);
   U10300 : OAI22_X1 port map( A1 => n60834, A2 => n61071, B1 => n892, B2 => 
                           n60830, ZN => n13880);
   U10301 : OAI22_X1 port map( A1 => n60835, A2 => n61085, B1 => n891, B2 => 
                           n60830, ZN => n13881);
   U10302 : OAI22_X1 port map( A1 => n60835, A2 => n61099, B1 => n890, B2 => 
                           n60830, ZN => n13882);
   U10303 : OAI22_X1 port map( A1 => n60835, A2 => n61113, B1 => n889, B2 => 
                           n60830, ZN => n13883);
   U10304 : OAI22_X1 port map( A1 => n60835, A2 => n61127, B1 => n888, B2 => 
                           n60830, ZN => n13884);
   U10305 : OAI22_X1 port map( A1 => n60363, A2 => n61970, B1 => n91, B2 => 
                           n15190, ZN => n12197);
   U10306 : OAI22_X1 port map( A1 => n60363, A2 => n61984, B1 => n90, B2 => 
                           n15190, ZN => n12198);
   U10307 : OAI22_X1 port map( A1 => n60363, A2 => n61998, B1 => n89, B2 => 
                           n15190, ZN => n12199);
   U10308 : OAI22_X1 port map( A1 => n60363, A2 => n62012, B1 => n88, B2 => 
                           n15190, ZN => n12200);
   U10309 : OAI22_X1 port map( A1 => n60363, A2 => n62026, B1 => n87, B2 => 
                           n15190, ZN => n12201);
   U10310 : OAI22_X1 port map( A1 => n60364, A2 => n62040, B1 => n86, B2 => 
                           n15190, ZN => n12202);
   U10311 : OAI22_X1 port map( A1 => n60364, A2 => n62054, B1 => n85, B2 => 
                           n15190, ZN => n12203);
   U10312 : OAI22_X1 port map( A1 => n60364, A2 => n62068, B1 => n84, B2 => 
                           n60362, ZN => n12204);
   U10313 : OAI22_X1 port map( A1 => n60364, A2 => n62082, B1 => n83, B2 => 
                           n60362, ZN => n12205);
   U10314 : OAI22_X1 port map( A1 => n60364, A2 => n62096, B1 => n82, B2 => 
                           n60362, ZN => n12206);
   U10315 : OAI22_X1 port map( A1 => n60365, A2 => n62110, B1 => n81, B2 => 
                           n60362, ZN => n12207);
   U10316 : OAI22_X1 port map( A1 => n60365, A2 => n60963, B1 => n80, B2 => 
                           n60362, ZN => n12208);
   U10317 : OAI22_X1 port map( A1 => n60129, A2 => n61972, B1 => n188, B2 => 
                           n60128, ZN => n11365);
   U10318 : OAI22_X1 port map( A1 => n60129, A2 => n61986, B1 => n187, B2 => 
                           n60128, ZN => n11366);
   U10319 : OAI22_X1 port map( A1 => n60129, A2 => n62000, B1 => n186, B2 => 
                           n60128, ZN => n11367);
   U10320 : OAI22_X1 port map( A1 => n60129, A2 => n62014, B1 => n185, B2 => 
                           n60128, ZN => n11368);
   U10321 : OAI22_X1 port map( A1 => n60129, A2 => n62028, B1 => n184, B2 => 
                           n60128, ZN => n11369);
   U10322 : OAI22_X1 port map( A1 => n60130, A2 => n62042, B1 => n183, B2 => 
                           n60128, ZN => n11370);
   U10323 : OAI22_X1 port map( A1 => n60130, A2 => n62056, B1 => n182, B2 => 
                           n60128, ZN => n11371);
   U10324 : OAI22_X1 port map( A1 => n60130, A2 => n62070, B1 => n181, B2 => 
                           n60128, ZN => n11372);
   U10325 : OAI22_X1 port map( A1 => n60130, A2 => n62084, B1 => n180, B2 => 
                           n60128, ZN => n11373);
   U10326 : OAI22_X1 port map( A1 => n60130, A2 => n62098, B1 => n179, B2 => 
                           n60128, ZN => n11374);
   U10327 : OAI22_X1 port map( A1 => n60131, A2 => n62112, B1 => n178, B2 => 
                           n60128, ZN => n11375);
   U10328 : OAI22_X1 port map( A1 => n60131, A2 => n60965, B1 => n177, B2 => 
                           n60128, ZN => n11376);
   U10329 : OAI22_X1 port map( A1 => n60131, A2 => n60979, B1 => n176, B2 => 
                           n15225, ZN => n11377);
   U10330 : OAI22_X1 port map( A1 => n60131, A2 => n60993, B1 => n175, B2 => 
                           n15225, ZN => n11378);
   U10331 : OAI22_X1 port map( A1 => n60131, A2 => n61007, B1 => n174, B2 => 
                           n15225, ZN => n11379);
   U10332 : OAI22_X1 port map( A1 => n60132, A2 => n61021, B1 => n173, B2 => 
                           n15225, ZN => n11380);
   U10333 : OAI22_X1 port map( A1 => n60132, A2 => n61035, B1 => n172, B2 => 
                           n15225, ZN => n11381);
   U10334 : OAI22_X1 port map( A1 => n60132, A2 => n61049, B1 => n171, B2 => 
                           n15225, ZN => n11382);
   U10335 : OAI22_X1 port map( A1 => n60132, A2 => n61063, B1 => n170, B2 => 
                           n15225, ZN => n11383);
   U10336 : OAI22_X1 port map( A1 => n60132, A2 => n61077, B1 => n169, B2 => 
                           n60128, ZN => n11384);
   U10337 : OAI22_X1 port map( A1 => n60133, A2 => n61091, B1 => n168, B2 => 
                           n60128, ZN => n11385);
   U10338 : OAI22_X1 port map( A1 => n60133, A2 => n61105, B1 => n167, B2 => 
                           n60128, ZN => n11386);
   U10339 : OAI22_X1 port map( A1 => n60133, A2 => n61119, B1 => n166, B2 => 
                           n60128, ZN => n11387);
   U10340 : OAI22_X1 port map( A1 => n60133, A2 => n61133, B1 => n165, B2 => 
                           n60128, ZN => n11388);
   U10341 : OAI22_X1 port map( A1 => n60120, A2 => n61972, B1 => n164, B2 => 
                           n60119, ZN => n11333);
   U10342 : OAI22_X1 port map( A1 => n60120, A2 => n61986, B1 => n163, B2 => 
                           n60119, ZN => n11334);
   U10343 : OAI22_X1 port map( A1 => n60120, A2 => n62000, B1 => n162, B2 => 
                           n60119, ZN => n11335);
   U10344 : OAI22_X1 port map( A1 => n60120, A2 => n62014, B1 => n161, B2 => 
                           n60119, ZN => n11336);
   U10345 : OAI22_X1 port map( A1 => n60120, A2 => n62028, B1 => n160, B2 => 
                           n60119, ZN => n11337);
   U10346 : OAI22_X1 port map( A1 => n60777, A2 => n61966, B1 => n3432, B2 => 
                           n60776, ZN => n13669);
   U10347 : OAI22_X1 port map( A1 => n60777, A2 => n61980, B1 => n3431, B2 => 
                           n60776, ZN => n13670);
   U10348 : OAI22_X1 port map( A1 => n60777, A2 => n61994, B1 => n3430, B2 => 
                           n60776, ZN => n13671);
   U10349 : OAI22_X1 port map( A1 => n60777, A2 => n62008, B1 => n3429, B2 => 
                           n60776, ZN => n13672);
   U10350 : OAI22_X1 port map( A1 => n60777, A2 => n62022, B1 => n3428, B2 => 
                           n60776, ZN => n13673);
   U10351 : OAI22_X1 port map( A1 => n60778, A2 => n62036, B1 => n3427, B2 => 
                           n60776, ZN => n13674);
   U10352 : OAI22_X1 port map( A1 => n60778, A2 => n62050, B1 => n3426, B2 => 
                           n60776, ZN => n13675);
   U10353 : OAI22_X1 port map( A1 => n60778, A2 => n62064, B1 => n3425, B2 => 
                           n60776, ZN => n13676);
   U10354 : OAI22_X1 port map( A1 => n60778, A2 => n62078, B1 => n3424, B2 => 
                           n60776, ZN => n13677);
   U10355 : OAI22_X1 port map( A1 => n60778, A2 => n62092, B1 => n3423, B2 => 
                           n60776, ZN => n13678);
   U10356 : OAI22_X1 port map( A1 => n60779, A2 => n62106, B1 => n3422, B2 => 
                           n60776, ZN => n13679);
   U10357 : OAI22_X1 port map( A1 => n60779, A2 => n60959, B1 => n3421, B2 => 
                           n60776, ZN => n13680);
   U10358 : OAI22_X1 port map( A1 => n60779, A2 => n60973, B1 => n3420, B2 => 
                           n15133, ZN => n13681);
   U10359 : OAI22_X1 port map( A1 => n60779, A2 => n60987, B1 => n3419, B2 => 
                           n15133, ZN => n13682);
   U10360 : OAI22_X1 port map( A1 => n60779, A2 => n61001, B1 => n3418, B2 => 
                           n15133, ZN => n13683);
   U10361 : OAI22_X1 port map( A1 => n60780, A2 => n61015, B1 => n3417, B2 => 
                           n15133, ZN => n13684);
   U10362 : OAI22_X1 port map( A1 => n60780, A2 => n61029, B1 => n3416, B2 => 
                           n15133, ZN => n13685);
   U10363 : OAI22_X1 port map( A1 => n60780, A2 => n61043, B1 => n3415, B2 => 
                           n15133, ZN => n13686);
   U10364 : OAI22_X1 port map( A1 => n60780, A2 => n61057, B1 => n3414, B2 => 
                           n15133, ZN => n13687);
   U10365 : OAI22_X1 port map( A1 => n60780, A2 => n61071, B1 => n3413, B2 => 
                           n60776, ZN => n13688);
   U10366 : OAI22_X1 port map( A1 => n60781, A2 => n61085, B1 => n3412, B2 => 
                           n60776, ZN => n13689);
   U10367 : OAI22_X1 port map( A1 => n60781, A2 => n61099, B1 => n3411, B2 => 
                           n60776, ZN => n13690);
   U10368 : OAI22_X1 port map( A1 => n60781, A2 => n61113, B1 => n3410, B2 => 
                           n60776, ZN => n13691);
   U10369 : OAI22_X1 port map( A1 => n60781, A2 => n61127, B1 => n3409, B2 => 
                           n60776, ZN => n13692);
   U10370 : OAI22_X1 port map( A1 => n59995, A2 => n62058, B1 => n5131, B2 => 
                           n59993, ZN => n10891);
   U10371 : OAI22_X1 port map( A1 => n59995, A2 => n62072, B1 => n5130, B2 => 
                           n59993, ZN => n10892);
   U10372 : OAI22_X1 port map( A1 => n59995, A2 => n62086, B1 => n5129, B2 => 
                           n59993, ZN => n10893);
   U10373 : OAI22_X1 port map( A1 => n59995, A2 => n62100, B1 => n5128, B2 => 
                           n59993, ZN => n10894);
   U10374 : OAI22_X1 port map( A1 => n59996, A2 => n62114, B1 => n5127, B2 => 
                           n59993, ZN => n10895);
   U10375 : OAI22_X1 port map( A1 => n59996, A2 => n60966, B1 => n5126, B2 => 
                           n59993, ZN => n10896);
   U10376 : OAI22_X1 port map( A1 => n59998, A2 => n61092, B1 => n5125, B2 => 
                           n15241, ZN => n10905);
   U10377 : OAI22_X1 port map( A1 => n59998, A2 => n61106, B1 => n5124, B2 => 
                           n15241, ZN => n10906);
   U10378 : OAI22_X1 port map( A1 => n59998, A2 => n61120, B1 => n5123, B2 => 
                           n15241, ZN => n10907);
   U10379 : OAI22_X1 port map( A1 => n59998, A2 => n61134, B1 => n5122, B2 => 
                           n15241, ZN => n10908);
   U10380 : OAI22_X1 port map( A1 => n59967, A2 => n61974, B1 => n5121, B2 => 
                           n59966, ZN => n10789);
   U10381 : OAI22_X1 port map( A1 => n59967, A2 => n61988, B1 => n5120, B2 => 
                           n59966, ZN => n10790);
   U10382 : OAI22_X1 port map( A1 => n59967, A2 => n62002, B1 => n5119, B2 => 
                           n59966, ZN => n10791);
   U10383 : OAI22_X1 port map( A1 => n59967, A2 => n62016, B1 => n5118, B2 => 
                           n59966, ZN => n10792);
   U10384 : OAI22_X1 port map( A1 => n59958, A2 => n61974, B1 => n5117, B2 => 
                           n59957, ZN => n10757);
   U10385 : OAI22_X1 port map( A1 => n59958, A2 => n61988, B1 => n5116, B2 => 
                           n59957, ZN => n10758);
   U10386 : OAI22_X1 port map( A1 => n59958, A2 => n62002, B1 => n5115, B2 => 
                           n59957, ZN => n10759);
   U10387 : OAI22_X1 port map( A1 => n59958, A2 => n62016, B1 => n5114, B2 => 
                           n59957, ZN => n10760);
   U10388 : OAI22_X1 port map( A1 => n59958, A2 => n62030, B1 => n5113, B2 => 
                           n59957, ZN => n10761);
   U10389 : OAI22_X1 port map( A1 => n59959, A2 => n62044, B1 => n5112, B2 => 
                           n59957, ZN => n10762);
   U10390 : OAI22_X1 port map( A1 => n59959, A2 => n62058, B1 => n5111, B2 => 
                           n59957, ZN => n10763);
   U10391 : OAI22_X1 port map( A1 => n59959, A2 => n62072, B1 => n5110, B2 => 
                           n59957, ZN => n10764);
   U10392 : OAI22_X1 port map( A1 => n59959, A2 => n62086, B1 => n5109, B2 => 
                           n59957, ZN => n10765);
   U10393 : OAI22_X1 port map( A1 => n59959, A2 => n62100, B1 => n5108, B2 => 
                           n59957, ZN => n10766);
   U10394 : OAI22_X1 port map( A1 => n59960, A2 => n62114, B1 => n5107, B2 => 
                           n59957, ZN => n10767);
   U10395 : OAI22_X1 port map( A1 => n59960, A2 => n60967, B1 => n5106, B2 => 
                           n59957, ZN => n10768);
   U10396 : OAI22_X1 port map( A1 => n59960, A2 => n60981, B1 => n5105, B2 => 
                           n15245, ZN => n10769);
   U10397 : OAI22_X1 port map( A1 => n59960, A2 => n60995, B1 => n5104, B2 => 
                           n15245, ZN => n10770);
   U10398 : OAI22_X1 port map( A1 => n59960, A2 => n61009, B1 => n5103, B2 => 
                           n15245, ZN => n10771);
   U10399 : OAI22_X1 port map( A1 => n59961, A2 => n61023, B1 => n5102, B2 => 
                           n15245, ZN => n10772);
   U10400 : OAI22_X1 port map( A1 => n59961, A2 => n61037, B1 => n5101, B2 => 
                           n15245, ZN => n10773);
   U10401 : OAI22_X1 port map( A1 => n59961, A2 => n61051, B1 => n5100, B2 => 
                           n15245, ZN => n10774);
   U10402 : OAI22_X1 port map( A1 => n59961, A2 => n61065, B1 => n5099, B2 => 
                           n15245, ZN => n10775);
   U10403 : OAI22_X1 port map( A1 => n59961, A2 => n61079, B1 => n5098, B2 => 
                           n59957, ZN => n10776);
   U10404 : OAI22_X1 port map( A1 => n59962, A2 => n61093, B1 => n5097, B2 => 
                           n59957, ZN => n10777);
   U10405 : OAI22_X1 port map( A1 => n59962, A2 => n61107, B1 => n5096, B2 => 
                           n59957, ZN => n10778);
   U10406 : OAI22_X1 port map( A1 => n59962, A2 => n61121, B1 => n5095, B2 => 
                           n59957, ZN => n10779);
   U10407 : OAI22_X1 port map( A1 => n59962, A2 => n61135, B1 => n5094, B2 => 
                           n59957, ZN => n10780);
   U10408 : OAI22_X1 port map( A1 => n59832, A2 => n61975, B1 => n5093, B2 => 
                           n59831, ZN => n10309);
   U10409 : OAI22_X1 port map( A1 => n59832, A2 => n61989, B1 => n5092, B2 => 
                           n59831, ZN => n10310);
   U10410 : OAI22_X1 port map( A1 => n59832, A2 => n62003, B1 => n5091, B2 => 
                           n59831, ZN => n10311);
   U10411 : OAI22_X1 port map( A1 => n59832, A2 => n62017, B1 => n5090, B2 => 
                           n59831, ZN => n10312);
   U10412 : OAI22_X1 port map( A1 => n59832, A2 => n62031, B1 => n5089, B2 => 
                           n59831, ZN => n10313);
   U10413 : OAI22_X1 port map( A1 => n59833, A2 => n62045, B1 => n5088, B2 => 
                           n59831, ZN => n10314);
   U10414 : OAI22_X1 port map( A1 => n59833, A2 => n62059, B1 => n5087, B2 => 
                           n59831, ZN => n10315);
   U10415 : OAI22_X1 port map( A1 => n59833, A2 => n62073, B1 => n5086, B2 => 
                           n59831, ZN => n10316);
   U10416 : OAI22_X1 port map( A1 => n59833, A2 => n62087, B1 => n5085, B2 => 
                           n59831, ZN => n10317);
   U10417 : OAI22_X1 port map( A1 => n59833, A2 => n62101, B1 => n5084, B2 => 
                           n59831, ZN => n10318);
   U10418 : OAI22_X1 port map( A1 => n59834, A2 => n62115, B1 => n5083, B2 => 
                           n59831, ZN => n10319);
   U10419 : OAI22_X1 port map( A1 => n59834, A2 => n60968, B1 => n5082, B2 => 
                           n59831, ZN => n10320);
   U10420 : OAI22_X1 port map( A1 => n59834, A2 => n60982, B1 => n5081, B2 => 
                           n15266, ZN => n10321);
   U10421 : OAI22_X1 port map( A1 => n59834, A2 => n60996, B1 => n5080, B2 => 
                           n15266, ZN => n10322);
   U10422 : OAI22_X1 port map( A1 => n59834, A2 => n61010, B1 => n5079, B2 => 
                           n15266, ZN => n10323);
   U10423 : OAI22_X1 port map( A1 => n59835, A2 => n61024, B1 => n5078, B2 => 
                           n15266, ZN => n10324);
   U10424 : OAI22_X1 port map( A1 => n59835, A2 => n61038, B1 => n5077, B2 => 
                           n15266, ZN => n10325);
   U10425 : OAI22_X1 port map( A1 => n59835, A2 => n61052, B1 => n5076, B2 => 
                           n15266, ZN => n10326);
   U10426 : OAI22_X1 port map( A1 => n59835, A2 => n61066, B1 => n5075, B2 => 
                           n15266, ZN => n10327);
   U10427 : OAI22_X1 port map( A1 => n59835, A2 => n61080, B1 => n5074, B2 => 
                           n59831, ZN => n10328);
   U10428 : OAI22_X1 port map( A1 => n59836, A2 => n61094, B1 => n5073, B2 => 
                           n59831, ZN => n10329);
   U10429 : OAI22_X1 port map( A1 => n59836, A2 => n61108, B1 => n5072, B2 => 
                           n59831, ZN => n10330);
   U10430 : OAI22_X1 port map( A1 => n59836, A2 => n61122, B1 => n5071, B2 => 
                           n59831, ZN => n10331);
   U10431 : OAI22_X1 port map( A1 => n59836, A2 => n61136, B1 => n5070, B2 => 
                           n59831, ZN => n10332);
   U10432 : OAI22_X1 port map( A1 => n59823, A2 => n61975, B1 => n5069, B2 => 
                           n59822, ZN => n10277);
   U10433 : OAI22_X1 port map( A1 => n59823, A2 => n61989, B1 => n5068, B2 => 
                           n59822, ZN => n10278);
   U10434 : OAI22_X1 port map( A1 => n59823, A2 => n62003, B1 => n5067, B2 => 
                           n59822, ZN => n10279);
   U10435 : OAI22_X1 port map( A1 => n59823, A2 => n62017, B1 => n5066, B2 => 
                           n59822, ZN => n10280);
   U10436 : OAI22_X1 port map( A1 => n59823, A2 => n62031, B1 => n5065, B2 => 
                           n59822, ZN => n10281);
   U10437 : OAI22_X1 port map( A1 => n59824, A2 => n62045, B1 => n5064, B2 => 
                           n59822, ZN => n10282);
   U10438 : OAI22_X1 port map( A1 => n59824, A2 => n62059, B1 => n5063, B2 => 
                           n59822, ZN => n10283);
   U10439 : OAI22_X1 port map( A1 => n59824, A2 => n62073, B1 => n5062, B2 => 
                           n59822, ZN => n10284);
   U10440 : OAI22_X1 port map( A1 => n59824, A2 => n62087, B1 => n5061, B2 => 
                           n59822, ZN => n10285);
   U10441 : OAI22_X1 port map( A1 => n59824, A2 => n62101, B1 => n5060, B2 => 
                           n59822, ZN => n10286);
   U10442 : OAI22_X1 port map( A1 => n59825, A2 => n62115, B1 => n5059, B2 => 
                           n59822, ZN => n10287);
   U10443 : OAI22_X1 port map( A1 => n59825, A2 => n60968, B1 => n5058, B2 => 
                           n59822, ZN => n10288);
   U10444 : OAI22_X1 port map( A1 => n59825, A2 => n60982, B1 => n5057, B2 => 
                           n15267, ZN => n10289);
   U10445 : OAI22_X1 port map( A1 => n59825, A2 => n60996, B1 => n5056, B2 => 
                           n15267, ZN => n10290);
   U10446 : OAI22_X1 port map( A1 => n59825, A2 => n61010, B1 => n5055, B2 => 
                           n15267, ZN => n10291);
   U10447 : OAI22_X1 port map( A1 => n59826, A2 => n61024, B1 => n5054, B2 => 
                           n15267, ZN => n10292);
   U10448 : OAI22_X1 port map( A1 => n59826, A2 => n61038, B1 => n5053, B2 => 
                           n15267, ZN => n10293);
   U10449 : OAI22_X1 port map( A1 => n59826, A2 => n61052, B1 => n5052, B2 => 
                           n15267, ZN => n10294);
   U10450 : OAI22_X1 port map( A1 => n59826, A2 => n61066, B1 => n5051, B2 => 
                           n15267, ZN => n10295);
   U10451 : OAI22_X1 port map( A1 => n59826, A2 => n61080, B1 => n5050, B2 => 
                           n59822, ZN => n10296);
   U10452 : OAI22_X1 port map( A1 => n60669, A2 => n61967, B1 => n53403, B2 => 
                           n60668, ZN => n13285);
   U10453 : OAI22_X1 port map( A1 => n60669, A2 => n61981, B1 => n53402, B2 => 
                           n60668, ZN => n13286);
   U10454 : OAI22_X1 port map( A1 => n60669, A2 => n61995, B1 => n53401, B2 => 
                           n60668, ZN => n13287);
   U10455 : OAI22_X1 port map( A1 => n60669, A2 => n62009, B1 => n53400, B2 => 
                           n60668, ZN => n13288);
   U10456 : OAI22_X1 port map( A1 => n60669, A2 => n62023, B1 => n53399, B2 => 
                           n60668, ZN => n13289);
   U10457 : OAI22_X1 port map( A1 => n60670, A2 => n62037, B1 => n53398, B2 => 
                           n60668, ZN => n13290);
   U10458 : OAI22_X1 port map( A1 => n60670, A2 => n62051, B1 => n53397, B2 => 
                           n60668, ZN => n13291);
   U10459 : OAI22_X1 port map( A1 => n60670, A2 => n62065, B1 => n53396, B2 => 
                           n60668, ZN => n13292);
   U10460 : OAI22_X1 port map( A1 => n60670, A2 => n62079, B1 => n53395, B2 => 
                           n60668, ZN => n13293);
   U10461 : OAI22_X1 port map( A1 => n60670, A2 => n62093, B1 => n53394, B2 => 
                           n60668, ZN => n13294);
   U10462 : OAI22_X1 port map( A1 => n60671, A2 => n62107, B1 => n53393, B2 => 
                           n60668, ZN => n13295);
   U10463 : OAI22_X1 port map( A1 => n60671, A2 => n60960, B1 => n53392, B2 => 
                           n60668, ZN => n13296);
   U10464 : OAI22_X1 port map( A1 => n60671, A2 => n60974, B1 => n53391, B2 => 
                           n15146, ZN => n13297);
   U10465 : OAI22_X1 port map( A1 => n60671, A2 => n60988, B1 => n53390, B2 => 
                           n15146, ZN => n13298);
   U10466 : OAI22_X1 port map( A1 => n60671, A2 => n61002, B1 => n53389, B2 => 
                           n15146, ZN => n13299);
   U10467 : OAI22_X1 port map( A1 => n60672, A2 => n61016, B1 => n53388, B2 => 
                           n15146, ZN => n13300);
   U10468 : OAI22_X1 port map( A1 => n60672, A2 => n61030, B1 => n53387, B2 => 
                           n15146, ZN => n13301);
   U10469 : OAI22_X1 port map( A1 => n60672, A2 => n61044, B1 => n53386, B2 => 
                           n15146, ZN => n13302);
   U10470 : OAI22_X1 port map( A1 => n60672, A2 => n61058, B1 => n53385, B2 => 
                           n15146, ZN => n13303);
   U10471 : OAI22_X1 port map( A1 => n60672, A2 => n61072, B1 => n53384, B2 => 
                           n60668, ZN => n13304);
   U10472 : OAI22_X1 port map( A1 => n60673, A2 => n61086, B1 => n53383, B2 => 
                           n60668, ZN => n13305);
   U10473 : OAI22_X1 port map( A1 => n60673, A2 => n61100, B1 => n53382, B2 => 
                           n60668, ZN => n13306);
   U10474 : OAI22_X1 port map( A1 => n60673, A2 => n61114, B1 => n53381, B2 => 
                           n60668, ZN => n13307);
   U10475 : OAI22_X1 port map( A1 => n60673, A2 => n61128, B1 => n53380, B2 => 
                           n60668, ZN => n13308);
   U10476 : OAI22_X1 port map( A1 => n60660, A2 => n61970, B1 => n53379, B2 => 
                           n60659, ZN => n13253);
   U10477 : OAI22_X1 port map( A1 => n60660, A2 => n61984, B1 => n53378, B2 => 
                           n60659, ZN => n13254);
   U10478 : OAI22_X1 port map( A1 => n60660, A2 => n61998, B1 => n53377, B2 => 
                           n60659, ZN => n13255);
   U10479 : OAI22_X1 port map( A1 => n60660, A2 => n62012, B1 => n53376, B2 => 
                           n60659, ZN => n13256);
   U10480 : OAI22_X1 port map( A1 => n60660, A2 => n62026, B1 => n53375, B2 => 
                           n60659, ZN => n13257);
   U10481 : OAI22_X1 port map( A1 => n60661, A2 => n62040, B1 => n53374, B2 => 
                           n60659, ZN => n13258);
   U10482 : OAI22_X1 port map( A1 => n60661, A2 => n62054, B1 => n53373, B2 => 
                           n60659, ZN => n13259);
   U10483 : OAI22_X1 port map( A1 => n60661, A2 => n62068, B1 => n53372, B2 => 
                           n60659, ZN => n13260);
   U10484 : OAI22_X1 port map( A1 => n60661, A2 => n62082, B1 => n53371, B2 => 
                           n60659, ZN => n13261);
   U10485 : OAI22_X1 port map( A1 => n60661, A2 => n62096, B1 => n53370, B2 => 
                           n60659, ZN => n13262);
   U10486 : OAI22_X1 port map( A1 => n60662, A2 => n62110, B1 => n53369, B2 => 
                           n60659, ZN => n13263);
   U10487 : OAI22_X1 port map( A1 => n60662, A2 => n60960, B1 => n53368, B2 => 
                           n60659, ZN => n13264);
   U10488 : OAI22_X1 port map( A1 => n60662, A2 => n60974, B1 => n53367, B2 => 
                           n15148, ZN => n13265);
   U10489 : OAI22_X1 port map( A1 => n60662, A2 => n60988, B1 => n53366, B2 => 
                           n15148, ZN => n13266);
   U10490 : OAI22_X1 port map( A1 => n60662, A2 => n61002, B1 => n53365, B2 => 
                           n15148, ZN => n13267);
   U10491 : OAI22_X1 port map( A1 => n60663, A2 => n61016, B1 => n53364, B2 => 
                           n15148, ZN => n13268);
   U10492 : OAI22_X1 port map( A1 => n60663, A2 => n61030, B1 => n53363, B2 => 
                           n15148, ZN => n13269);
   U10493 : OAI22_X1 port map( A1 => n60663, A2 => n61044, B1 => n53362, B2 => 
                           n15148, ZN => n13270);
   U10494 : OAI22_X1 port map( A1 => n60663, A2 => n61058, B1 => n53361, B2 => 
                           n15148, ZN => n13271);
   U10495 : OAI22_X1 port map( A1 => n60663, A2 => n61072, B1 => n53360, B2 => 
                           n60659, ZN => n13272);
   U10496 : OAI22_X1 port map( A1 => n60664, A2 => n61086, B1 => n53359, B2 => 
                           n60659, ZN => n13273);
   U10497 : OAI22_X1 port map( A1 => n60664, A2 => n61100, B1 => n53358, B2 => 
                           n60659, ZN => n13274);
   U10498 : OAI22_X1 port map( A1 => n60664, A2 => n61114, B1 => n53357, B2 => 
                           n60659, ZN => n13275);
   U10499 : OAI22_X1 port map( A1 => n60664, A2 => n61128, B1 => n53356, B2 => 
                           n60659, ZN => n13276);
   U10500 : OAI22_X1 port map( A1 => n60651, A2 => n61967, B1 => n5001, B2 => 
                           n60650, ZN => n13221);
   U10501 : OAI22_X1 port map( A1 => n60651, A2 => n61981, B1 => n5000, B2 => 
                           n60650, ZN => n13222);
   U10502 : OAI22_X1 port map( A1 => n60651, A2 => n61995, B1 => n4999, B2 => 
                           n60650, ZN => n13223);
   U10503 : OAI22_X1 port map( A1 => n60651, A2 => n62009, B1 => n4998, B2 => 
                           n60650, ZN => n13224);
   U10504 : OAI22_X1 port map( A1 => n60651, A2 => n62023, B1 => n4997, B2 => 
                           n60650, ZN => n13225);
   U10505 : OAI22_X1 port map( A1 => n60652, A2 => n62037, B1 => n4996, B2 => 
                           n60650, ZN => n13226);
   U10506 : OAI22_X1 port map( A1 => n60652, A2 => n62051, B1 => n4995, B2 => 
                           n60650, ZN => n13227);
   U10507 : OAI22_X1 port map( A1 => n60652, A2 => n62065, B1 => n4994, B2 => 
                           n60650, ZN => n13228);
   U10508 : OAI22_X1 port map( A1 => n60652, A2 => n62079, B1 => n4993, B2 => 
                           n60650, ZN => n13229);
   U10509 : OAI22_X1 port map( A1 => n60652, A2 => n62093, B1 => n4992, B2 => 
                           n60650, ZN => n13230);
   U10510 : OAI22_X1 port map( A1 => n60653, A2 => n62107, B1 => n4991, B2 => 
                           n60650, ZN => n13231);
   U10511 : OAI22_X1 port map( A1 => n60653, A2 => n60960, B1 => n4990, B2 => 
                           n60650, ZN => n13232);
   U10512 : OAI22_X1 port map( A1 => n60653, A2 => n60974, B1 => n4989, B2 => 
                           n15149, ZN => n13233);
   U10513 : OAI22_X1 port map( A1 => n60653, A2 => n60988, B1 => n4988, B2 => 
                           n15149, ZN => n13234);
   U10514 : OAI22_X1 port map( A1 => n60653, A2 => n61002, B1 => n4987, B2 => 
                           n15149, ZN => n13235);
   U10515 : OAI22_X1 port map( A1 => n60654, A2 => n61016, B1 => n4986, B2 => 
                           n15149, ZN => n13236);
   U10516 : OAI22_X1 port map( A1 => n60654, A2 => n61030, B1 => n4985, B2 => 
                           n15149, ZN => n13237);
   U10517 : OAI22_X1 port map( A1 => n60654, A2 => n61044, B1 => n4984, B2 => 
                           n15149, ZN => n13238);
   U10518 : OAI22_X1 port map( A1 => n60654, A2 => n61058, B1 => n4983, B2 => 
                           n15149, ZN => n13239);
   U10519 : OAI22_X1 port map( A1 => n60654, A2 => n61072, B1 => n4982, B2 => 
                           n60650, ZN => n13240);
   U10520 : OAI22_X1 port map( A1 => n60655, A2 => n61086, B1 => n4981, B2 => 
                           n60650, ZN => n13241);
   U10521 : OAI22_X1 port map( A1 => n60655, A2 => n61100, B1 => n4980, B2 => 
                           n60650, ZN => n13242);
   U10522 : OAI22_X1 port map( A1 => n60655, A2 => n61114, B1 => n4979, B2 => 
                           n60650, ZN => n13243);
   U10523 : OAI22_X1 port map( A1 => n60655, A2 => n61128, B1 => n4978, B2 => 
                           n60650, ZN => n13244);
   U10524 : OAI22_X1 port map( A1 => n60642, A2 => n61967, B1 => n4977, B2 => 
                           n60641, ZN => n13189);
   U10525 : OAI22_X1 port map( A1 => n60642, A2 => n61981, B1 => n4976, B2 => 
                           n60641, ZN => n13190);
   U10526 : OAI22_X1 port map( A1 => n60642, A2 => n61995, B1 => n4975, B2 => 
                           n60641, ZN => n13191);
   U10527 : OAI22_X1 port map( A1 => n60642, A2 => n62009, B1 => n4974, B2 => 
                           n60641, ZN => n13192);
   U10528 : OAI22_X1 port map( A1 => n60642, A2 => n62023, B1 => n4973, B2 => 
                           n60641, ZN => n13193);
   U10529 : OAI22_X1 port map( A1 => n60643, A2 => n62037, B1 => n4972, B2 => 
                           n60641, ZN => n13194);
   U10530 : OAI22_X1 port map( A1 => n60643, A2 => n62051, B1 => n4971, B2 => 
                           n60641, ZN => n13195);
   U10531 : OAI22_X1 port map( A1 => n60643, A2 => n62065, B1 => n4970, B2 => 
                           n60641, ZN => n13196);
   U10532 : OAI22_X1 port map( A1 => n60643, A2 => n62079, B1 => n4969, B2 => 
                           n60641, ZN => n13197);
   U10533 : OAI22_X1 port map( A1 => n60643, A2 => n62093, B1 => n4968, B2 => 
                           n60641, ZN => n13198);
   U10534 : OAI22_X1 port map( A1 => n60644, A2 => n62107, B1 => n4967, B2 => 
                           n60641, ZN => n13199);
   U10535 : OAI22_X1 port map( A1 => n60644, A2 => n60960, B1 => n4966, B2 => 
                           n60641, ZN => n13200);
   U10536 : OAI22_X1 port map( A1 => n60644, A2 => n60974, B1 => n4965, B2 => 
                           n15150, ZN => n13201);
   U10537 : OAI22_X1 port map( A1 => n60644, A2 => n60988, B1 => n4964, B2 => 
                           n15150, ZN => n13202);
   U10538 : OAI22_X1 port map( A1 => n60644, A2 => n61002, B1 => n4963, B2 => 
                           n15150, ZN => n13203);
   U10539 : OAI22_X1 port map( A1 => n60645, A2 => n61016, B1 => n4962, B2 => 
                           n15150, ZN => n13204);
   U10540 : OAI22_X1 port map( A1 => n60645, A2 => n61030, B1 => n4961, B2 => 
                           n15150, ZN => n13205);
   U10541 : OAI22_X1 port map( A1 => n60645, A2 => n61044, B1 => n4960, B2 => 
                           n15150, ZN => n13206);
   U10542 : OAI22_X1 port map( A1 => n60645, A2 => n61058, B1 => n4959, B2 => 
                           n15150, ZN => n13207);
   U10543 : OAI22_X1 port map( A1 => n60645, A2 => n61072, B1 => n4958, B2 => 
                           n60641, ZN => n13208);
   U10544 : OAI22_X1 port map( A1 => n60646, A2 => n61086, B1 => n4957, B2 => 
                           n60641, ZN => n13209);
   U10545 : OAI22_X1 port map( A1 => n60646, A2 => n61100, B1 => n4956, B2 => 
                           n60641, ZN => n13210);
   U10546 : OAI22_X1 port map( A1 => n60646, A2 => n61114, B1 => n4955, B2 => 
                           n60641, ZN => n13211);
   U10547 : OAI22_X1 port map( A1 => n60646, A2 => n61128, B1 => n4954, B2 => 
                           n60641, ZN => n13212);
   U10548 : OAI22_X1 port map( A1 => n60615, A2 => n61968, B1 => n9778, B2 => 
                           n60614, ZN => n13093);
   U10549 : OAI22_X1 port map( A1 => n60615, A2 => n61982, B1 => n9777, B2 => 
                           n60614, ZN => n13094);
   U10550 : OAI22_X1 port map( A1 => n60615, A2 => n61996, B1 => n9776, B2 => 
                           n60614, ZN => n13095);
   U10551 : OAI22_X1 port map( A1 => n60615, A2 => n62010, B1 => n9775, B2 => 
                           n60614, ZN => n13096);
   U10552 : OAI22_X1 port map( A1 => n60615, A2 => n62024, B1 => n9774, B2 => 
                           n60614, ZN => n13097);
   U10553 : OAI22_X1 port map( A1 => n60616, A2 => n62038, B1 => n9773, B2 => 
                           n60614, ZN => n13098);
   U10554 : OAI22_X1 port map( A1 => n60616, A2 => n62052, B1 => n9772, B2 => 
                           n60614, ZN => n13099);
   U10555 : OAI22_X1 port map( A1 => n60616, A2 => n62066, B1 => n9771, B2 => 
                           n60614, ZN => n13100);
   U10556 : OAI22_X1 port map( A1 => n60616, A2 => n62080, B1 => n9770, B2 => 
                           n60614, ZN => n13101);
   U10557 : OAI22_X1 port map( A1 => n60616, A2 => n62094, B1 => n9769, B2 => 
                           n60614, ZN => n13102);
   U10558 : OAI22_X1 port map( A1 => n60617, A2 => n62108, B1 => n9768, B2 => 
                           n60614, ZN => n13103);
   U10559 : OAI22_X1 port map( A1 => n60617, A2 => n60961, B1 => n9767, B2 => 
                           n60614, ZN => n13104);
   U10560 : OAI22_X1 port map( A1 => n60617, A2 => n60975, B1 => n9766, B2 => 
                           n15153, ZN => n13105);
   U10561 : OAI22_X1 port map( A1 => n60617, A2 => n60989, B1 => n9765, B2 => 
                           n15153, ZN => n13106);
   U10562 : OAI22_X1 port map( A1 => n60617, A2 => n61003, B1 => n9764, B2 => 
                           n15153, ZN => n13107);
   U10563 : OAI22_X1 port map( A1 => n60618, A2 => n61017, B1 => n9763, B2 => 
                           n15153, ZN => n13108);
   U10564 : OAI22_X1 port map( A1 => n60618, A2 => n61031, B1 => n9762, B2 => 
                           n15153, ZN => n13109);
   U10565 : OAI22_X1 port map( A1 => n60618, A2 => n61045, B1 => n9761, B2 => 
                           n15153, ZN => n13110);
   U10566 : OAI22_X1 port map( A1 => n60618, A2 => n61059, B1 => n9760, B2 => 
                           n15153, ZN => n13111);
   U10567 : OAI22_X1 port map( A1 => n60618, A2 => n61073, B1 => n9759, B2 => 
                           n60614, ZN => n13112);
   U10568 : OAI22_X1 port map( A1 => n60619, A2 => n61087, B1 => n9758, B2 => 
                           n60614, ZN => n13113);
   U10569 : OAI22_X1 port map( A1 => n60619, A2 => n61101, B1 => n9757, B2 => 
                           n60614, ZN => n13114);
   U10570 : OAI22_X1 port map( A1 => n60619, A2 => n61115, B1 => n9756, B2 => 
                           n60614, ZN => n13115);
   U10571 : OAI22_X1 port map( A1 => n60619, A2 => n61129, B1 => n9755, B2 => 
                           n60614, ZN => n13116);
   U10572 : OAI22_X1 port map( A1 => n60606, A2 => n61968, B1 => n9810, B2 => 
                           n60605, ZN => n13061);
   U10573 : OAI22_X1 port map( A1 => n60606, A2 => n61982, B1 => n9809, B2 => 
                           n60605, ZN => n13062);
   U10574 : OAI22_X1 port map( A1 => n60606, A2 => n61996, B1 => n9808, B2 => 
                           n60605, ZN => n13063);
   U10575 : OAI22_X1 port map( A1 => n60606, A2 => n62010, B1 => n9807, B2 => 
                           n60605, ZN => n13064);
   U10576 : OAI22_X1 port map( A1 => n60606, A2 => n62024, B1 => n9806, B2 => 
                           n60605, ZN => n13065);
   U10577 : OAI22_X1 port map( A1 => n60607, A2 => n62038, B1 => n9805, B2 => 
                           n60605, ZN => n13066);
   U10578 : OAI22_X1 port map( A1 => n60607, A2 => n62052, B1 => n9804, B2 => 
                           n60605, ZN => n13067);
   U10579 : OAI22_X1 port map( A1 => n60607, A2 => n62066, B1 => n9803, B2 => 
                           n60605, ZN => n13068);
   U10580 : OAI22_X1 port map( A1 => n60607, A2 => n62080, B1 => n9802, B2 => 
                           n60605, ZN => n13069);
   U10581 : OAI22_X1 port map( A1 => n60607, A2 => n62094, B1 => n9801, B2 => 
                           n60605, ZN => n13070);
   U10582 : OAI22_X1 port map( A1 => n60608, A2 => n62108, B1 => n9800, B2 => 
                           n60605, ZN => n13071);
   U10583 : OAI22_X1 port map( A1 => n60608, A2 => n60961, B1 => n9799, B2 => 
                           n60605, ZN => n13072);
   U10584 : OAI22_X1 port map( A1 => n60608, A2 => n60975, B1 => n9798, B2 => 
                           n15154, ZN => n13073);
   U10585 : OAI22_X1 port map( A1 => n60608, A2 => n60989, B1 => n9797, B2 => 
                           n15154, ZN => n13074);
   U10586 : OAI22_X1 port map( A1 => n60608, A2 => n61003, B1 => n9796, B2 => 
                           n15154, ZN => n13075);
   U10587 : OAI22_X1 port map( A1 => n60609, A2 => n61017, B1 => n9795, B2 => 
                           n15154, ZN => n13076);
   U10588 : OAI22_X1 port map( A1 => n60609, A2 => n61031, B1 => n9794, B2 => 
                           n15154, ZN => n13077);
   U10589 : OAI22_X1 port map( A1 => n60609, A2 => n61045, B1 => n9793, B2 => 
                           n15154, ZN => n13078);
   U10590 : OAI22_X1 port map( A1 => n60609, A2 => n61059, B1 => n9792, B2 => 
                           n15154, ZN => n13079);
   U10591 : OAI22_X1 port map( A1 => n60609, A2 => n61073, B1 => n9791, B2 => 
                           n60605, ZN => n13080);
   U10592 : OAI22_X1 port map( A1 => n60610, A2 => n61087, B1 => n9790, B2 => 
                           n60605, ZN => n13081);
   U10593 : OAI22_X1 port map( A1 => n60610, A2 => n61101, B1 => n9789, B2 => 
                           n60605, ZN => n13082);
   U10594 : OAI22_X1 port map( A1 => n60610, A2 => n61115, B1 => n9788, B2 => 
                           n60605, ZN => n13083);
   U10595 : OAI22_X1 port map( A1 => n60610, A2 => n61129, B1 => n9787, B2 => 
                           n60605, ZN => n13084);
   U10596 : OAI22_X1 port map( A1 => n60579, A2 => n61968, B1 => n4905, B2 => 
                           n60578, ZN => n12965);
   U10597 : OAI22_X1 port map( A1 => n60579, A2 => n61982, B1 => n4904, B2 => 
                           n60578, ZN => n12966);
   U10598 : OAI22_X1 port map( A1 => n60579, A2 => n61996, B1 => n4903, B2 => 
                           n60578, ZN => n12967);
   U10599 : OAI22_X1 port map( A1 => n60579, A2 => n62010, B1 => n4902, B2 => 
                           n60578, ZN => n12968);
   U10600 : OAI22_X1 port map( A1 => n60579, A2 => n62024, B1 => n4901, B2 => 
                           n60578, ZN => n12969);
   U10601 : OAI22_X1 port map( A1 => n60580, A2 => n62038, B1 => n4900, B2 => 
                           n60578, ZN => n12970);
   U10602 : OAI22_X1 port map( A1 => n60580, A2 => n62052, B1 => n4899, B2 => 
                           n60578, ZN => n12971);
   U10603 : OAI22_X1 port map( A1 => n60580, A2 => n62066, B1 => n4898, B2 => 
                           n60578, ZN => n12972);
   U10604 : OAI22_X1 port map( A1 => n60580, A2 => n62080, B1 => n4897, B2 => 
                           n60578, ZN => n12973);
   U10605 : OAI22_X1 port map( A1 => n60580, A2 => n62094, B1 => n4896, B2 => 
                           n60578, ZN => n12974);
   U10606 : OAI22_X1 port map( A1 => n60581, A2 => n62108, B1 => n4895, B2 => 
                           n60578, ZN => n12975);
   U10607 : OAI22_X1 port map( A1 => n60581, A2 => n60961, B1 => n4894, B2 => 
                           n60578, ZN => n12976);
   U10608 : OAI22_X1 port map( A1 => n60581, A2 => n60975, B1 => n4893, B2 => 
                           n15157, ZN => n12977);
   U10609 : OAI22_X1 port map( A1 => n60581, A2 => n60989, B1 => n4892, B2 => 
                           n15157, ZN => n12978);
   U10610 : OAI22_X1 port map( A1 => n60581, A2 => n61003, B1 => n4891, B2 => 
                           n15157, ZN => n12979);
   U10611 : OAI22_X1 port map( A1 => n60582, A2 => n61017, B1 => n4890, B2 => 
                           n15157, ZN => n12980);
   U10612 : OAI22_X1 port map( A1 => n60582, A2 => n61031, B1 => n4889, B2 => 
                           n15157, ZN => n12981);
   U10613 : OAI22_X1 port map( A1 => n60582, A2 => n61045, B1 => n4888, B2 => 
                           n15157, ZN => n12982);
   U10614 : OAI22_X1 port map( A1 => n60582, A2 => n61059, B1 => n4887, B2 => 
                           n15157, ZN => n12983);
   U10615 : OAI22_X1 port map( A1 => n60582, A2 => n61073, B1 => n4886, B2 => 
                           n60578, ZN => n12984);
   U10616 : OAI22_X1 port map( A1 => n60583, A2 => n61087, B1 => n4885, B2 => 
                           n60578, ZN => n12985);
   U10617 : OAI22_X1 port map( A1 => n60583, A2 => n61101, B1 => n4884, B2 => 
                           n60578, ZN => n12986);
   U10618 : OAI22_X1 port map( A1 => n60583, A2 => n61115, B1 => n4883, B2 => 
                           n60578, ZN => n12987);
   U10619 : OAI22_X1 port map( A1 => n60583, A2 => n61129, B1 => n4882, B2 => 
                           n60578, ZN => n12988);
   U10620 : OAI22_X1 port map( A1 => n60570, A2 => n61968, B1 => n4881, B2 => 
                           n60569, ZN => n12933);
   U10621 : OAI22_X1 port map( A1 => n60570, A2 => n61982, B1 => n4880, B2 => 
                           n60569, ZN => n12934);
   U10622 : OAI22_X1 port map( A1 => n60570, A2 => n61996, B1 => n4879, B2 => 
                           n60569, ZN => n12935);
   U10623 : OAI22_X1 port map( A1 => n60570, A2 => n62010, B1 => n4878, B2 => 
                           n60569, ZN => n12936);
   U10624 : OAI22_X1 port map( A1 => n60570, A2 => n62024, B1 => n4877, B2 => 
                           n60569, ZN => n12937);
   U10625 : OAI22_X1 port map( A1 => n60571, A2 => n62038, B1 => n4876, B2 => 
                           n60569, ZN => n12938);
   U10626 : OAI22_X1 port map( A1 => n60571, A2 => n62052, B1 => n4875, B2 => 
                           n60569, ZN => n12939);
   U10627 : OAI22_X1 port map( A1 => n60571, A2 => n62066, B1 => n4874, B2 => 
                           n60569, ZN => n12940);
   U10628 : OAI22_X1 port map( A1 => n60571, A2 => n62080, B1 => n4873, B2 => 
                           n60569, ZN => n12941);
   U10629 : OAI22_X1 port map( A1 => n60571, A2 => n62094, B1 => n4872, B2 => 
                           n60569, ZN => n12942);
   U10630 : OAI22_X1 port map( A1 => n60572, A2 => n62108, B1 => n4871, B2 => 
                           n60569, ZN => n12943);
   U10631 : OAI22_X1 port map( A1 => n60572, A2 => n60961, B1 => n4870, B2 => 
                           n60569, ZN => n12944);
   U10632 : OAI22_X1 port map( A1 => n60572, A2 => n60975, B1 => n4869, B2 => 
                           n15158, ZN => n12945);
   U10633 : OAI22_X1 port map( A1 => n60572, A2 => n60989, B1 => n4868, B2 => 
                           n15158, ZN => n12946);
   U10634 : OAI22_X1 port map( A1 => n60572, A2 => n61003, B1 => n4867, B2 => 
                           n15158, ZN => n12947);
   U10635 : OAI22_X1 port map( A1 => n60573, A2 => n61017, B1 => n4866, B2 => 
                           n15158, ZN => n12948);
   U10636 : OAI22_X1 port map( A1 => n60573, A2 => n61031, B1 => n4865, B2 => 
                           n15158, ZN => n12949);
   U10637 : OAI22_X1 port map( A1 => n60573, A2 => n61045, B1 => n4864, B2 => 
                           n15158, ZN => n12950);
   U10638 : OAI22_X1 port map( A1 => n60573, A2 => n61059, B1 => n4863, B2 => 
                           n15158, ZN => n12951);
   U10639 : OAI22_X1 port map( A1 => n60573, A2 => n61073, B1 => n4862, B2 => 
                           n60569, ZN => n12952);
   U10640 : OAI22_X1 port map( A1 => n60574, A2 => n61087, B1 => n4861, B2 => 
                           n60569, ZN => n12953);
   U10641 : OAI22_X1 port map( A1 => n60574, A2 => n61101, B1 => n4860, B2 => 
                           n60569, ZN => n12954);
   U10642 : OAI22_X1 port map( A1 => n60574, A2 => n61115, B1 => n4859, B2 => 
                           n60569, ZN => n12955);
   U10643 : OAI22_X1 port map( A1 => n60574, A2 => n61129, B1 => n4858, B2 => 
                           n60569, ZN => n12956);
   U10644 : OAI22_X1 port map( A1 => n60563, A2 => n62108, B1 => n53257, B2 => 
                           n60560, ZN => n12911);
   U10645 : OAI22_X1 port map( A1 => n60563, A2 => n60961, B1 => n53256, B2 => 
                           n60560, ZN => n12912);
   U10646 : OAI22_X1 port map( A1 => n60563, A2 => n60975, B1 => n53255, B2 => 
                           n15159, ZN => n12913);
   U10647 : OAI22_X1 port map( A1 => n60563, A2 => n60989, B1 => n53254, B2 => 
                           n15159, ZN => n12914);
   U10648 : OAI22_X1 port map( A1 => n60563, A2 => n61003, B1 => n53253, B2 => 
                           n15159, ZN => n12915);
   U10649 : OAI22_X1 port map( A1 => n60564, A2 => n61017, B1 => n53252, B2 => 
                           n15159, ZN => n12916);
   U10650 : OAI22_X1 port map( A1 => n60564, A2 => n61031, B1 => n53251, B2 => 
                           n15159, ZN => n12917);
   U10651 : OAI22_X1 port map( A1 => n60564, A2 => n61045, B1 => n53250, B2 => 
                           n15159, ZN => n12918);
   U10652 : OAI22_X1 port map( A1 => n60564, A2 => n61059, B1 => n53249, B2 => 
                           n15159, ZN => n12919);
   U10653 : OAI22_X1 port map( A1 => n60564, A2 => n61073, B1 => n53248, B2 => 
                           n60560, ZN => n12920);
   U10654 : OAI22_X1 port map( A1 => n60565, A2 => n61087, B1 => n53247, B2 => 
                           n60560, ZN => n12921);
   U10655 : OAI22_X1 port map( A1 => n60565, A2 => n61101, B1 => n53246, B2 => 
                           n60560, ZN => n12922);
   U10656 : OAI22_X1 port map( A1 => n60565, A2 => n61115, B1 => n53245, B2 => 
                           n60560, ZN => n12923);
   U10657 : OAI22_X1 port map( A1 => n60565, A2 => n61129, B1 => n53244, B2 => 
                           n60560, ZN => n12924);
   U10658 : OAI22_X1 port map( A1 => n60527, A2 => n62108, B1 => n53185, B2 => 
                           n60524, ZN => n12783);
   U10659 : OAI22_X1 port map( A1 => n60527, A2 => n60962, B1 => n53184, B2 => 
                           n60524, ZN => n12784);
   U10660 : OAI22_X1 port map( A1 => n60527, A2 => n60976, B1 => n53183, B2 => 
                           n15163, ZN => n12785);
   U10661 : OAI22_X1 port map( A1 => n60527, A2 => n60990, B1 => n53182, B2 => 
                           n15163, ZN => n12786);
   U10662 : OAI22_X1 port map( A1 => n60527, A2 => n61004, B1 => n53181, B2 => 
                           n15163, ZN => n12787);
   U10663 : OAI22_X1 port map( A1 => n60528, A2 => n61018, B1 => n53180, B2 => 
                           n15163, ZN => n12788);
   U10664 : OAI22_X1 port map( A1 => n60528, A2 => n61032, B1 => n53179, B2 => 
                           n15163, ZN => n12789);
   U10665 : OAI22_X1 port map( A1 => n60528, A2 => n61046, B1 => n53178, B2 => 
                           n15163, ZN => n12790);
   U10666 : OAI22_X1 port map( A1 => n60528, A2 => n61060, B1 => n53177, B2 => 
                           n15163, ZN => n12791);
   U10667 : OAI22_X1 port map( A1 => n60528, A2 => n61074, B1 => n53176, B2 => 
                           n60524, ZN => n12792);
   U10668 : OAI22_X1 port map( A1 => n60529, A2 => n61088, B1 => n53175, B2 => 
                           n60524, ZN => n12793);
   U10669 : OAI22_X1 port map( A1 => n60529, A2 => n61102, B1 => n53174, B2 => 
                           n60524, ZN => n12794);
   U10670 : OAI22_X1 port map( A1 => n60529, A2 => n61116, B1 => n53173, B2 => 
                           n60524, ZN => n12795);
   U10671 : OAI22_X1 port map( A1 => n60529, A2 => n61130, B1 => n53172, B2 => 
                           n60524, ZN => n12796);
   U10672 : OAI22_X1 port map( A1 => n60417, A2 => n61969, B1 => n53051, B2 => 
                           n60416, ZN => n12389);
   U10673 : OAI22_X1 port map( A1 => n60417, A2 => n61983, B1 => n53050, B2 => 
                           n60416, ZN => n12390);
   U10674 : OAI22_X1 port map( A1 => n60417, A2 => n61997, B1 => n53049, B2 => 
                           n60416, ZN => n12391);
   U10675 : OAI22_X1 port map( A1 => n60417, A2 => n62011, B1 => n53048, B2 => 
                           n60416, ZN => n12392);
   U10676 : OAI22_X1 port map( A1 => n60417, A2 => n62025, B1 => n53047, B2 => 
                           n60416, ZN => n12393);
   U10677 : OAI22_X1 port map( A1 => n60418, A2 => n62039, B1 => n53046, B2 => 
                           n60416, ZN => n12394);
   U10678 : OAI22_X1 port map( A1 => n60418, A2 => n62053, B1 => n53045, B2 => 
                           n60416, ZN => n12395);
   U10679 : OAI22_X1 port map( A1 => n60418, A2 => n62067, B1 => n53044, B2 => 
                           n60416, ZN => n12396);
   U10680 : OAI22_X1 port map( A1 => n60418, A2 => n62081, B1 => n53043, B2 => 
                           n60416, ZN => n12397);
   U10681 : OAI22_X1 port map( A1 => n60418, A2 => n62095, B1 => n53042, B2 => 
                           n60416, ZN => n12398);
   U10682 : OAI22_X1 port map( A1 => n60419, A2 => n62109, B1 => n53041, B2 => 
                           n60416, ZN => n12399);
   U10683 : OAI22_X1 port map( A1 => n60419, A2 => n60963, B1 => n53040, B2 => 
                           n60416, ZN => n12400);
   U10684 : OAI22_X1 port map( A1 => n60419, A2 => n60977, B1 => n53039, B2 => 
                           n15183, ZN => n12401);
   U10685 : OAI22_X1 port map( A1 => n60419, A2 => n60991, B1 => n53038, B2 => 
                           n15183, ZN => n12402);
   U10686 : OAI22_X1 port map( A1 => n60419, A2 => n61005, B1 => n53037, B2 => 
                           n15183, ZN => n12403);
   U10687 : OAI22_X1 port map( A1 => n60420, A2 => n61019, B1 => n53036, B2 => 
                           n15183, ZN => n12404);
   U10688 : OAI22_X1 port map( A1 => n60420, A2 => n61033, B1 => n53035, B2 => 
                           n15183, ZN => n12405);
   U10689 : OAI22_X1 port map( A1 => n60420, A2 => n61047, B1 => n53034, B2 => 
                           n15183, ZN => n12406);
   U10690 : OAI22_X1 port map( A1 => n60420, A2 => n61061, B1 => n53033, B2 => 
                           n15183, ZN => n12407);
   U10691 : OAI22_X1 port map( A1 => n60420, A2 => n61075, B1 => n53032, B2 => 
                           n60416, ZN => n12408);
   U10692 : OAI22_X1 port map( A1 => n60421, A2 => n61089, B1 => n53031, B2 => 
                           n60416, ZN => n12409);
   U10693 : OAI22_X1 port map( A1 => n60421, A2 => n61103, B1 => n53030, B2 => 
                           n60416, ZN => n12410);
   U10694 : OAI22_X1 port map( A1 => n60421, A2 => n61117, B1 => n53029, B2 => 
                           n60416, ZN => n12411);
   U10695 : OAI22_X1 port map( A1 => n60421, A2 => n61131, B1 => n53028, B2 => 
                           n60416, ZN => n12412);
   U10696 : OAI22_X1 port map( A1 => n60941, A2 => n61000, B1 => n53583, B2 => 
                           n15098, ZN => n14259);
   U10697 : OAI22_X1 port map( A1 => n60942, A2 => n61014, B1 => n53582, B2 => 
                           n15098, ZN => n14260);
   U10698 : OAI22_X1 port map( A1 => n60942, A2 => n61028, B1 => n53581, B2 => 
                           n15098, ZN => n14261);
   U10699 : OAI22_X1 port map( A1 => n60942, A2 => n61042, B1 => n53580, B2 => 
                           n15098, ZN => n14262);
   U10700 : OAI22_X1 port map( A1 => n60942, A2 => n61056, B1 => n53579, B2 => 
                           n60938, ZN => n14263);
   U10701 : OAI22_X1 port map( A1 => n60942, A2 => n61070, B1 => n53578, B2 => 
                           n60938, ZN => n14264);
   U10702 : OAI22_X1 port map( A1 => n60943, A2 => n61084, B1 => n53577, B2 => 
                           n60938, ZN => n14265);
   U10703 : OAI22_X1 port map( A1 => n60943, A2 => n61098, B1 => n53576, B2 => 
                           n60938, ZN => n14266);
   U10704 : OAI22_X1 port map( A1 => n60943, A2 => n61126, B1 => n53575, B2 => 
                           n60938, ZN => n14268);
   U10705 : OAI22_X1 port map( A1 => n60930, A2 => n61965, B1 => n53574, B2 => 
                           n60929, ZN => n14213);
   U10706 : OAI22_X1 port map( A1 => n60930, A2 => n61979, B1 => n53573, B2 => 
                           n60929, ZN => n14214);
   U10707 : OAI22_X1 port map( A1 => n60930, A2 => n61993, B1 => n53572, B2 => 
                           n60929, ZN => n14215);
   U10708 : OAI22_X1 port map( A1 => n60903, A2 => n61965, B1 => n53571, B2 => 
                           n60902, ZN => n14117);
   U10709 : OAI22_X1 port map( A1 => n60903, A2 => n61979, B1 => n53570, B2 => 
                           n60902, ZN => n14118);
   U10710 : OAI22_X1 port map( A1 => n60903, A2 => n61993, B1 => n53569, B2 => 
                           n60902, ZN => n14119);
   U10711 : OAI22_X1 port map( A1 => n60903, A2 => n62007, B1 => n53568, B2 => 
                           n60902, ZN => n14120);
   U10712 : OAI22_X1 port map( A1 => n60903, A2 => n62021, B1 => n53567, B2 => 
                           n60902, ZN => n14121);
   U10713 : OAI22_X1 port map( A1 => n60904, A2 => n62035, B1 => n53566, B2 => 
                           n60902, ZN => n14122);
   U10714 : OAI22_X1 port map( A1 => n60904, A2 => n62049, B1 => n53565, B2 => 
                           n60902, ZN => n14123);
   U10715 : OAI22_X1 port map( A1 => n60904, A2 => n62063, B1 => n53564, B2 => 
                           n60902, ZN => n14124);
   U10716 : OAI22_X1 port map( A1 => n60904, A2 => n62077, B1 => n53563, B2 => 
                           n60902, ZN => n14125);
   U10717 : OAI22_X1 port map( A1 => n60904, A2 => n62091, B1 => n53562, B2 => 
                           n60902, ZN => n14126);
   U10718 : OAI22_X1 port map( A1 => n60905, A2 => n62105, B1 => n53561, B2 => 
                           n60902, ZN => n14127);
   U10719 : OAI22_X1 port map( A1 => n60905, A2 => n60958, B1 => n53560, B2 => 
                           n60902, ZN => n14128);
   U10720 : OAI22_X1 port map( A1 => n60905, A2 => n60972, B1 => n53559, B2 => 
                           n15106, ZN => n14129);
   U10721 : OAI22_X1 port map( A1 => n60905, A2 => n60986, B1 => n53558, B2 => 
                           n15106, ZN => n14130);
   U10722 : OAI22_X1 port map( A1 => n60905, A2 => n61000, B1 => n53557, B2 => 
                           n15106, ZN => n14131);
   U10723 : OAI22_X1 port map( A1 => n60906, A2 => n61014, B1 => n53556, B2 => 
                           n15106, ZN => n14132);
   U10724 : OAI22_X1 port map( A1 => n60906, A2 => n61028, B1 => n53555, B2 => 
                           n15106, ZN => n14133);
   U10725 : OAI22_X1 port map( A1 => n60906, A2 => n61042, B1 => n53554, B2 => 
                           n15106, ZN => n14134);
   U10726 : OAI22_X1 port map( A1 => n60906, A2 => n61056, B1 => n53553, B2 => 
                           n15106, ZN => n14135);
   U10727 : OAI22_X1 port map( A1 => n60906, A2 => n61070, B1 => n53552, B2 => 
                           n60902, ZN => n14136);
   U10728 : OAI22_X1 port map( A1 => n60907, A2 => n61084, B1 => n53551, B2 => 
                           n60902, ZN => n14137);
   U10729 : OAI22_X1 port map( A1 => n60907, A2 => n61098, B1 => n53550, B2 => 
                           n60902, ZN => n14138);
   U10730 : OAI22_X1 port map( A1 => n60907, A2 => n61112, B1 => n53549, B2 => 
                           n60902, ZN => n14139);
   U10731 : OAI22_X1 port map( A1 => n60907, A2 => n61126, B1 => n53548, B2 => 
                           n60902, ZN => n14140);
   U10732 : OAI22_X1 port map( A1 => n60858, A2 => n61965, B1 => n935, B2 => 
                           n60857, ZN => n13957);
   U10733 : OAI22_X1 port map( A1 => n60858, A2 => n61979, B1 => n934, B2 => 
                           n60857, ZN => n13958);
   U10734 : OAI22_X1 port map( A1 => n60858, A2 => n61993, B1 => n933, B2 => 
                           n60857, ZN => n13959);
   U10735 : OAI22_X1 port map( A1 => n60858, A2 => n62007, B1 => n932, B2 => 
                           n60857, ZN => n13960);
   U10736 : OAI22_X1 port map( A1 => n60858, A2 => n62021, B1 => n931, B2 => 
                           n60857, ZN => n13961);
   U10737 : OAI22_X1 port map( A1 => n60859, A2 => n62035, B1 => n930, B2 => 
                           n60857, ZN => n13962);
   U10738 : OAI22_X1 port map( A1 => n60859, A2 => n62049, B1 => n929, B2 => 
                           n60857, ZN => n13963);
   U10739 : OAI22_X1 port map( A1 => n60859, A2 => n62063, B1 => n928, B2 => 
                           n60857, ZN => n13964);
   U10740 : OAI22_X1 port map( A1 => n60859, A2 => n62077, B1 => n927, B2 => 
                           n60857, ZN => n13965);
   U10741 : OAI22_X1 port map( A1 => n60859, A2 => n62091, B1 => n926, B2 => 
                           n60857, ZN => n13966);
   U10742 : OAI22_X1 port map( A1 => n60860, A2 => n62105, B1 => n925, B2 => 
                           n60857, ZN => n13967);
   U10743 : OAI22_X1 port map( A1 => n60860, A2 => n60958, B1 => n924, B2 => 
                           n60857, ZN => n13968);
   U10744 : OAI22_X1 port map( A1 => n60860, A2 => n60972, B1 => n923, B2 => 
                           n15116, ZN => n13969);
   U10745 : OAI22_X1 port map( A1 => n60860, A2 => n60986, B1 => n922, B2 => 
                           n15116, ZN => n13970);
   U10746 : OAI22_X1 port map( A1 => n60860, A2 => n61000, B1 => n921, B2 => 
                           n15116, ZN => n13971);
   U10747 : OAI22_X1 port map( A1 => n60861, A2 => n61014, B1 => n920, B2 => 
                           n15116, ZN => n13972);
   U10748 : OAI22_X1 port map( A1 => n60861, A2 => n61028, B1 => n919, B2 => 
                           n15116, ZN => n13973);
   U10749 : OAI22_X1 port map( A1 => n60861, A2 => n61042, B1 => n918, B2 => 
                           n15116, ZN => n13974);
   U10750 : OAI22_X1 port map( A1 => n60861, A2 => n61056, B1 => n917, B2 => 
                           n15116, ZN => n13975);
   U10751 : OAI22_X1 port map( A1 => n60861, A2 => n61070, B1 => n916, B2 => 
                           n60857, ZN => n13976);
   U10752 : OAI22_X1 port map( A1 => n60862, A2 => n61084, B1 => n915, B2 => 
                           n60857, ZN => n13977);
   U10753 : OAI22_X1 port map( A1 => n60862, A2 => n61098, B1 => n914, B2 => 
                           n60857, ZN => n13978);
   U10754 : OAI22_X1 port map( A1 => n60862, A2 => n61112, B1 => n913, B2 => 
                           n60857, ZN => n13979);
   U10755 : OAI22_X1 port map( A1 => n60862, A2 => n61126, B1 => n912, B2 => 
                           n60857, ZN => n13980);
   U10756 : OAI22_X1 port map( A1 => n60822, A2 => n61966, B1 => n887, B2 => 
                           n60821, ZN => n13829);
   U10757 : OAI22_X1 port map( A1 => n60822, A2 => n61980, B1 => n886, B2 => 
                           n60821, ZN => n13830);
   U10758 : OAI22_X1 port map( A1 => n60822, A2 => n61994, B1 => n885, B2 => 
                           n60821, ZN => n13831);
   U10759 : OAI22_X1 port map( A1 => n60822, A2 => n62008, B1 => n884, B2 => 
                           n60821, ZN => n13832);
   U10760 : OAI22_X1 port map( A1 => n60822, A2 => n62022, B1 => n883, B2 => 
                           n60821, ZN => n13833);
   U10761 : OAI22_X1 port map( A1 => n60823, A2 => n62036, B1 => n882, B2 => 
                           n60821, ZN => n13834);
   U10762 : OAI22_X1 port map( A1 => n60823, A2 => n62050, B1 => n881, B2 => 
                           n60821, ZN => n13835);
   U10763 : OAI22_X1 port map( A1 => n60823, A2 => n62064, B1 => n880, B2 => 
                           n60821, ZN => n13836);
   U10764 : OAI22_X1 port map( A1 => n60823, A2 => n62078, B1 => n879, B2 => 
                           n60821, ZN => n13837);
   U10765 : OAI22_X1 port map( A1 => n60823, A2 => n62092, B1 => n878, B2 => 
                           n60821, ZN => n13838);
   U10766 : OAI22_X1 port map( A1 => n60824, A2 => n62106, B1 => n877, B2 => 
                           n60821, ZN => n13839);
   U10767 : OAI22_X1 port map( A1 => n60824, A2 => n60959, B1 => n876, B2 => 
                           n60821, ZN => n13840);
   U10768 : OAI22_X1 port map( A1 => n60824, A2 => n60973, B1 => n875, B2 => 
                           n15124, ZN => n13841);
   U10769 : OAI22_X1 port map( A1 => n60824, A2 => n60987, B1 => n874, B2 => 
                           n15124, ZN => n13842);
   U10770 : OAI22_X1 port map( A1 => n60824, A2 => n61001, B1 => n873, B2 => 
                           n15124, ZN => n13843);
   U10771 : OAI22_X1 port map( A1 => n60825, A2 => n61015, B1 => n872, B2 => 
                           n15124, ZN => n13844);
   U10772 : OAI22_X1 port map( A1 => n60825, A2 => n61029, B1 => n871, B2 => 
                           n15124, ZN => n13845);
   U10773 : OAI22_X1 port map( A1 => n60825, A2 => n61043, B1 => n870, B2 => 
                           n15124, ZN => n13846);
   U10774 : OAI22_X1 port map( A1 => n60825, A2 => n61057, B1 => n869, B2 => 
                           n15124, ZN => n13847);
   U10775 : OAI22_X1 port map( A1 => n60825, A2 => n61071, B1 => n868, B2 => 
                           n60821, ZN => n13848);
   U10776 : OAI22_X1 port map( A1 => n60826, A2 => n61085, B1 => n867, B2 => 
                           n60821, ZN => n13849);
   U10777 : OAI22_X1 port map( A1 => n60826, A2 => n61099, B1 => n866, B2 => 
                           n60821, ZN => n13850);
   U10778 : OAI22_X1 port map( A1 => n60826, A2 => n61113, B1 => n865, B2 => 
                           n60821, ZN => n13851);
   U10779 : OAI22_X1 port map( A1 => n60826, A2 => n61127, B1 => n864, B2 => 
                           n60821, ZN => n13852);
   U10780 : OAI22_X1 port map( A1 => n60894, A2 => n61965, B1 => n53427, B2 => 
                           n60893, ZN => n14085);
   U10781 : OAI22_X1 port map( A1 => n60894, A2 => n61979, B1 => n53426, B2 => 
                           n60893, ZN => n14086);
   U10782 : OAI22_X1 port map( A1 => n60894, A2 => n61993, B1 => n53425, B2 => 
                           n60893, ZN => n14087);
   U10783 : OAI22_X1 port map( A1 => n60894, A2 => n62007, B1 => n53424, B2 => 
                           n60893, ZN => n14088);
   U10784 : OAI22_X1 port map( A1 => n60894, A2 => n62021, B1 => n53423, B2 => 
                           n60893, ZN => n14089);
   U10785 : OAI22_X1 port map( A1 => n60895, A2 => n62035, B1 => n53422, B2 => 
                           n60893, ZN => n14090);
   U10786 : OAI22_X1 port map( A1 => n60895, A2 => n62049, B1 => n53421, B2 => 
                           n60893, ZN => n14091);
   U10787 : OAI22_X1 port map( A1 => n60895, A2 => n62063, B1 => n53420, B2 => 
                           n60893, ZN => n14092);
   U10788 : OAI22_X1 port map( A1 => n60895, A2 => n62077, B1 => n53419, B2 => 
                           n60893, ZN => n14093);
   U10789 : OAI22_X1 port map( A1 => n60895, A2 => n62091, B1 => n53418, B2 => 
                           n60893, ZN => n14094);
   U10790 : OAI22_X1 port map( A1 => n60896, A2 => n62105, B1 => n53417, B2 => 
                           n60893, ZN => n14095);
   U10791 : OAI22_X1 port map( A1 => n60896, A2 => n60958, B1 => n53416, B2 => 
                           n60893, ZN => n14096);
   U10792 : OAI22_X1 port map( A1 => n60896, A2 => n60972, B1 => n53415, B2 => 
                           n15108, ZN => n14097);
   U10793 : OAI22_X1 port map( A1 => n60896, A2 => n60986, B1 => n53414, B2 => 
                           n15108, ZN => n14098);
   U10794 : OAI22_X1 port map( A1 => n60896, A2 => n61000, B1 => n53413, B2 => 
                           n15108, ZN => n14099);
   U10795 : OAI22_X1 port map( A1 => n60897, A2 => n61014, B1 => n53412, B2 => 
                           n15108, ZN => n14100);
   U10796 : OAI22_X1 port map( A1 => n60897, A2 => n61028, B1 => n53411, B2 => 
                           n15108, ZN => n14101);
   U10797 : OAI22_X1 port map( A1 => n60897, A2 => n61042, B1 => n53410, B2 => 
                           n15108, ZN => n14102);
   U10798 : OAI22_X1 port map( A1 => n60897, A2 => n61056, B1 => n53409, B2 => 
                           n15108, ZN => n14103);
   U10799 : OAI22_X1 port map( A1 => n60897, A2 => n61070, B1 => n53408, B2 => 
                           n60893, ZN => n14104);
   U10800 : OAI22_X1 port map( A1 => n60898, A2 => n61084, B1 => n53407, B2 => 
                           n60893, ZN => n14105);
   U10801 : OAI22_X1 port map( A1 => n60898, A2 => n61098, B1 => n53406, B2 => 
                           n60893, ZN => n14106);
   U10802 : OAI22_X1 port map( A1 => n60898, A2 => n61112, B1 => n53405, B2 => 
                           n60893, ZN => n14107);
   U10803 : OAI22_X1 port map( A1 => n60898, A2 => n61126, B1 => n53404, B2 => 
                           n60893, ZN => n14108);
   U10804 : OAI22_X1 port map( A1 => n60174, A2 => n61972, B1 => n4431, B2 => 
                           n60173, ZN => n11525);
   U10805 : OAI22_X1 port map( A1 => n60174, A2 => n61986, B1 => n4430, B2 => 
                           n60173, ZN => n11526);
   U10806 : OAI22_X1 port map( A1 => n60174, A2 => n62000, B1 => n4429, B2 => 
                           n60173, ZN => n11527);
   U10807 : OAI22_X1 port map( A1 => n60174, A2 => n62014, B1 => n4428, B2 => 
                           n60173, ZN => n11528);
   U10808 : OAI22_X1 port map( A1 => n60174, A2 => n62028, B1 => n4427, B2 => 
                           n60173, ZN => n11529);
   U10809 : OAI22_X1 port map( A1 => n60175, A2 => n62042, B1 => n4426, B2 => 
                           n60173, ZN => n11530);
   U10810 : OAI22_X1 port map( A1 => n60175, A2 => n62056, B1 => n4425, B2 => 
                           n60173, ZN => n11531);
   U10811 : OAI22_X1 port map( A1 => n60175, A2 => n62070, B1 => n4424, B2 => 
                           n60173, ZN => n11532);
   U10812 : OAI22_X1 port map( A1 => n60175, A2 => n62084, B1 => n4423, B2 => 
                           n60173, ZN => n11533);
   U10813 : OAI22_X1 port map( A1 => n60175, A2 => n62098, B1 => n4422, B2 => 
                           n60173, ZN => n11534);
   U10814 : OAI22_X1 port map( A1 => n60176, A2 => n62112, B1 => n4421, B2 => 
                           n60173, ZN => n11535);
   U10815 : OAI22_X1 port map( A1 => n60176, A2 => n60965, B1 => n4420, B2 => 
                           n60173, ZN => n11536);
   U10816 : OAI22_X1 port map( A1 => n60176, A2 => n60979, B1 => n4419, B2 => 
                           n15220, ZN => n11537);
   U10817 : OAI22_X1 port map( A1 => n60176, A2 => n60993, B1 => n4418, B2 => 
                           n15220, ZN => n11538);
   U10818 : OAI22_X1 port map( A1 => n60176, A2 => n61007, B1 => n4417, B2 => 
                           n15220, ZN => n11539);
   U10819 : OAI22_X1 port map( A1 => n60177, A2 => n61021, B1 => n4416, B2 => 
                           n15220, ZN => n11540);
   U10820 : OAI22_X1 port map( A1 => n60177, A2 => n61035, B1 => n4415, B2 => 
                           n15220, ZN => n11541);
   U10821 : OAI22_X1 port map( A1 => n60177, A2 => n61049, B1 => n4414, B2 => 
                           n15220, ZN => n11542);
   U10822 : OAI22_X1 port map( A1 => n60177, A2 => n61063, B1 => n4413, B2 => 
                           n15220, ZN => n11543);
   U10823 : OAI22_X1 port map( A1 => n60177, A2 => n61077, B1 => n4412, B2 => 
                           n60173, ZN => n11544);
   U10824 : OAI22_X1 port map( A1 => n60178, A2 => n61091, B1 => n4411, B2 => 
                           n60173, ZN => n11545);
   U10825 : OAI22_X1 port map( A1 => n60178, A2 => n61105, B1 => n4410, B2 => 
                           n60173, ZN => n11546);
   U10826 : OAI22_X1 port map( A1 => n60178, A2 => n61119, B1 => n4409, B2 => 
                           n60173, ZN => n11547);
   U10827 : OAI22_X1 port map( A1 => n60178, A2 => n61133, B1 => n4408, B2 => 
                           n60173, ZN => n11548);
   U10828 : OAI22_X1 port map( A1 => n60813, A2 => n61966, B1 => n591, B2 => 
                           n60812, ZN => n13797);
   U10829 : OAI22_X1 port map( A1 => n60813, A2 => n61980, B1 => n590, B2 => 
                           n60812, ZN => n13798);
   U10830 : OAI22_X1 port map( A1 => n60813, A2 => n61994, B1 => n589, B2 => 
                           n60812, ZN => n13799);
   U10831 : OAI22_X1 port map( A1 => n60813, A2 => n62008, B1 => n588, B2 => 
                           n60812, ZN => n13800);
   U10832 : OAI22_X1 port map( A1 => n60813, A2 => n62022, B1 => n587, B2 => 
                           n60812, ZN => n13801);
   U10833 : OAI22_X1 port map( A1 => n60814, A2 => n62036, B1 => n586, B2 => 
                           n60812, ZN => n13802);
   U10834 : OAI22_X1 port map( A1 => n60814, A2 => n62050, B1 => n585, B2 => 
                           n60812, ZN => n13803);
   U10835 : OAI22_X1 port map( A1 => n60814, A2 => n62064, B1 => n584, B2 => 
                           n60812, ZN => n13804);
   U10836 : OAI22_X1 port map( A1 => n60814, A2 => n62078, B1 => n583, B2 => 
                           n60812, ZN => n13805);
   U10837 : OAI22_X1 port map( A1 => n60814, A2 => n62092, B1 => n582, B2 => 
                           n60812, ZN => n13806);
   U10838 : OAI22_X1 port map( A1 => n60815, A2 => n62106, B1 => n581, B2 => 
                           n60812, ZN => n13807);
   U10839 : OAI22_X1 port map( A1 => n60815, A2 => n60959, B1 => n580, B2 => 
                           n60812, ZN => n13808);
   U10840 : OAI22_X1 port map( A1 => n60815, A2 => n60973, B1 => n579, B2 => 
                           n15128, ZN => n13809);
   U10841 : OAI22_X1 port map( A1 => n60815, A2 => n60987, B1 => n578, B2 => 
                           n15128, ZN => n13810);
   U10842 : OAI22_X1 port map( A1 => n60815, A2 => n61001, B1 => n577, B2 => 
                           n15128, ZN => n13811);
   U10843 : OAI22_X1 port map( A1 => n60816, A2 => n61015, B1 => n576, B2 => 
                           n15128, ZN => n13812);
   U10844 : OAI22_X1 port map( A1 => n60816, A2 => n61029, B1 => n575, B2 => 
                           n15128, ZN => n13813);
   U10845 : OAI22_X1 port map( A1 => n60816, A2 => n61043, B1 => n574, B2 => 
                           n15128, ZN => n13814);
   U10846 : OAI22_X1 port map( A1 => n60816, A2 => n61057, B1 => n573, B2 => 
                           n15128, ZN => n13815);
   U10847 : OAI22_X1 port map( A1 => n60816, A2 => n61071, B1 => n572, B2 => 
                           n60812, ZN => n13816);
   U10848 : OAI22_X1 port map( A1 => n60817, A2 => n61085, B1 => n571, B2 => 
                           n60812, ZN => n13817);
   U10849 : OAI22_X1 port map( A1 => n60817, A2 => n61099, B1 => n570, B2 => 
                           n60812, ZN => n13818);
   U10850 : OAI22_X1 port map( A1 => n60817, A2 => n61113, B1 => n569, B2 => 
                           n60812, ZN => n13819);
   U10851 : OAI22_X1 port map( A1 => n60817, A2 => n61127, B1 => n568, B2 => 
                           n60812, ZN => n13820);
   U10852 : OAI22_X1 port map( A1 => n60804, A2 => n61966, B1 => n53003, B2 => 
                           n60803, ZN => n13765);
   U10853 : OAI22_X1 port map( A1 => n60804, A2 => n61980, B1 => n53002, B2 => 
                           n60803, ZN => n13766);
   U10854 : OAI22_X1 port map( A1 => n60804, A2 => n61994, B1 => n53001, B2 => 
                           n60803, ZN => n13767);
   U10855 : OAI22_X1 port map( A1 => n60804, A2 => n62008, B1 => n53000, B2 => 
                           n60803, ZN => n13768);
   U10856 : OAI22_X1 port map( A1 => n60804, A2 => n62022, B1 => n52999, B2 => 
                           n60803, ZN => n13769);
   U10857 : OAI22_X1 port map( A1 => n60805, A2 => n62036, B1 => n52998, B2 => 
                           n60803, ZN => n13770);
   U10858 : OAI22_X1 port map( A1 => n60805, A2 => n62050, B1 => n52997, B2 => 
                           n60803, ZN => n13771);
   U10859 : OAI22_X1 port map( A1 => n60805, A2 => n62064, B1 => n52996, B2 => 
                           n60803, ZN => n13772);
   U10860 : OAI22_X1 port map( A1 => n60805, A2 => n62078, B1 => n52995, B2 => 
                           n60803, ZN => n13773);
   U10861 : OAI22_X1 port map( A1 => n60805, A2 => n62092, B1 => n52994, B2 => 
                           n60803, ZN => n13774);
   U10862 : OAI22_X1 port map( A1 => n60806, A2 => n62106, B1 => n52993, B2 => 
                           n60803, ZN => n13775);
   U10863 : OAI22_X1 port map( A1 => n60806, A2 => n60959, B1 => n52992, B2 => 
                           n60803, ZN => n13776);
   U10864 : OAI22_X1 port map( A1 => n60806, A2 => n60973, B1 => n52991, B2 => 
                           n15130, ZN => n13777);
   U10865 : OAI22_X1 port map( A1 => n60806, A2 => n60987, B1 => n52990, B2 => 
                           n15130, ZN => n13778);
   U10866 : OAI22_X1 port map( A1 => n60806, A2 => n61001, B1 => n52989, B2 => 
                           n15130, ZN => n13779);
   U10867 : OAI22_X1 port map( A1 => n60807, A2 => n61015, B1 => n52988, B2 => 
                           n15130, ZN => n13780);
   U10868 : OAI22_X1 port map( A1 => n60807, A2 => n61029, B1 => n52987, B2 => 
                           n15130, ZN => n13781);
   U10869 : OAI22_X1 port map( A1 => n60807, A2 => n61043, B1 => n52986, B2 => 
                           n15130, ZN => n13782);
   U10870 : OAI22_X1 port map( A1 => n60807, A2 => n61057, B1 => n52985, B2 => 
                           n15130, ZN => n13783);
   U10871 : OAI22_X1 port map( A1 => n60807, A2 => n61071, B1 => n52984, B2 => 
                           n60803, ZN => n13784);
   U10872 : OAI22_X1 port map( A1 => n60808, A2 => n61085, B1 => n52983, B2 => 
                           n60803, ZN => n13785);
   U10873 : OAI22_X1 port map( A1 => n60808, A2 => n61099, B1 => n52982, B2 => 
                           n60803, ZN => n13786);
   U10874 : OAI22_X1 port map( A1 => n60808, A2 => n61113, B1 => n52981, B2 => 
                           n60803, ZN => n13787);
   U10875 : OAI22_X1 port map( A1 => n60808, A2 => n61127, B1 => n52980, B2 => 
                           n60803, ZN => n13788);
   U10876 : OAI22_X1 port map( A1 => n60714, A2 => n61967, B1 => n52955, B2 => 
                           n15140, ZN => n13445);
   U10877 : OAI22_X1 port map( A1 => n60714, A2 => n61981, B1 => n52954, B2 => 
                           n15140, ZN => n13446);
   U10878 : OAI22_X1 port map( A1 => n60714, A2 => n61995, B1 => n52953, B2 => 
                           n15140, ZN => n13447);
   U10879 : OAI22_X1 port map( A1 => n60714, A2 => n62009, B1 => n52952, B2 => 
                           n15140, ZN => n13448);
   U10880 : OAI22_X1 port map( A1 => n60715, A2 => n62037, B1 => n51826, B2 => 
                           n15140, ZN => n13450);
   U10881 : OAI22_X1 port map( A1 => n60715, A2 => n62051, B1 => n51825, B2 => 
                           n15140, ZN => n13451);
   U10882 : OAI22_X1 port map( A1 => n60715, A2 => n62065, B1 => n51824, B2 => 
                           n15140, ZN => n13452);
   U10883 : OAI22_X1 port map( A1 => n60715, A2 => n62079, B1 => n51823, B2 => 
                           n60713, ZN => n13453);
   U10884 : OAI22_X1 port map( A1 => n60715, A2 => n62093, B1 => n51822, B2 => 
                           n60713, ZN => n13454);
   U10885 : OAI22_X1 port map( A1 => n60716, A2 => n62107, B1 => n51821, B2 => 
                           n60713, ZN => n13455);
   U10886 : OAI22_X1 port map( A1 => n60716, A2 => n60960, B1 => n51820, B2 => 
                           n60713, ZN => n13456);
   U10887 : OAI22_X1 port map( A1 => n60716, A2 => n60974, B1 => n51819, B2 => 
                           n60713, ZN => n13457);
   U10888 : OAI22_X1 port map( A1 => n60716, A2 => n60988, B1 => n51818, B2 => 
                           n60713, ZN => n13458);
   U10889 : OAI22_X1 port map( A1 => n60716, A2 => n61002, B1 => n51817, B2 => 
                           n60713, ZN => n13459);
   U10890 : OAI22_X1 port map( A1 => n60717, A2 => n61016, B1 => n51816, B2 => 
                           n60713, ZN => n13460);
   U10891 : OAI22_X1 port map( A1 => n60717, A2 => n61030, B1 => n51815, B2 => 
                           n60713, ZN => n13461);
   U10892 : OAI22_X1 port map( A1 => n60717, A2 => n61044, B1 => n51814, B2 => 
                           n60713, ZN => n13462);
   U10893 : OAI22_X1 port map( A1 => n60717, A2 => n61058, B1 => n51813, B2 => 
                           n60713, ZN => n13463);
   U10894 : OAI22_X1 port map( A1 => n60717, A2 => n61072, B1 => n51812, B2 => 
                           n60713, ZN => n13464);
   U10895 : OAI22_X1 port map( A1 => n60718, A2 => n61086, B1 => n51811, B2 => 
                           n60713, ZN => n13465);
   U10896 : OAI22_X1 port map( A1 => n60718, A2 => n61100, B1 => n51810, B2 => 
                           n60713, ZN => n13466);
   U10897 : OAI22_X1 port map( A1 => n60718, A2 => n61114, B1 => n51809, B2 => 
                           n60713, ZN => n13467);
   U10898 : OAI22_X1 port map( A1 => n60718, A2 => n61128, B1 => n51808, B2 => 
                           n60713, ZN => n13468);
   U10899 : OAI22_X1 port map( A1 => n60705, A2 => n61967, B1 => n52951, B2 => 
                           n60704, ZN => n13413);
   U10900 : OAI22_X1 port map( A1 => n60705, A2 => n61981, B1 => n52950, B2 => 
                           n60704, ZN => n13414);
   U10901 : OAI22_X1 port map( A1 => n60705, A2 => n61995, B1 => n52949, B2 => 
                           n60704, ZN => n13415);
   U10902 : OAI22_X1 port map( A1 => n60705, A2 => n62009, B1 => n52948, B2 => 
                           n60704, ZN => n13416);
   U10903 : OAI22_X1 port map( A1 => n60705, A2 => n62023, B1 => n52947, B2 => 
                           n60704, ZN => n13417);
   U10904 : OAI22_X1 port map( A1 => n60706, A2 => n62037, B1 => n52946, B2 => 
                           n60704, ZN => n13418);
   U10905 : OAI22_X1 port map( A1 => n60706, A2 => n62051, B1 => n52945, B2 => 
                           n60704, ZN => n13419);
   U10906 : OAI22_X1 port map( A1 => n60706, A2 => n62065, B1 => n52944, B2 => 
                           n60704, ZN => n13420);
   U10907 : OAI22_X1 port map( A1 => n60706, A2 => n62079, B1 => n52943, B2 => 
                           n60704, ZN => n13421);
   U10908 : OAI22_X1 port map( A1 => n60706, A2 => n62093, B1 => n52942, B2 => 
                           n60704, ZN => n13422);
   U10909 : OAI22_X1 port map( A1 => n60707, A2 => n62107, B1 => n52941, B2 => 
                           n60704, ZN => n13423);
   U10910 : OAI22_X1 port map( A1 => n60707, A2 => n60960, B1 => n52940, B2 => 
                           n60704, ZN => n13424);
   U10911 : OAI22_X1 port map( A1 => n60707, A2 => n60974, B1 => n52939, B2 => 
                           n15141, ZN => n13425);
   U10912 : OAI22_X1 port map( A1 => n60707, A2 => n60988, B1 => n52938, B2 => 
                           n15141, ZN => n13426);
   U10913 : OAI22_X1 port map( A1 => n60707, A2 => n61002, B1 => n52937, B2 => 
                           n15141, ZN => n13427);
   U10914 : OAI22_X1 port map( A1 => n60708, A2 => n61016, B1 => n52936, B2 => 
                           n15141, ZN => n13428);
   U10915 : OAI22_X1 port map( A1 => n60708, A2 => n61030, B1 => n52935, B2 => 
                           n15141, ZN => n13429);
   U10916 : OAI22_X1 port map( A1 => n60708, A2 => n61044, B1 => n52934, B2 => 
                           n15141, ZN => n13430);
   U10917 : OAI22_X1 port map( A1 => n60708, A2 => n61058, B1 => n52933, B2 => 
                           n15141, ZN => n13431);
   U10918 : OAI22_X1 port map( A1 => n60708, A2 => n61072, B1 => n52932, B2 => 
                           n60704, ZN => n13432);
   U10919 : OAI22_X1 port map( A1 => n60709, A2 => n61086, B1 => n52931, B2 => 
                           n60704, ZN => n13433);
   U10920 : OAI22_X1 port map( A1 => n60709, A2 => n61100, B1 => n52930, B2 => 
                           n60704, ZN => n13434);
   U10921 : OAI22_X1 port map( A1 => n60709, A2 => n61114, B1 => n52929, B2 => 
                           n60704, ZN => n13435);
   U10922 : OAI22_X1 port map( A1 => n60709, A2 => n61128, B1 => n52928, B2 => 
                           n60704, ZN => n13436);
   U10923 : OAI22_X1 port map( A1 => n60066, A2 => n61973, B1 => n3846, B2 => 
                           n60065, ZN => n11141);
   U10924 : OAI22_X1 port map( A1 => n60066, A2 => n61987, B1 => n3845, B2 => 
                           n60065, ZN => n11142);
   U10925 : OAI22_X1 port map( A1 => n60066, A2 => n62001, B1 => n3844, B2 => 
                           n60065, ZN => n11143);
   U10926 : OAI22_X1 port map( A1 => n60066, A2 => n62015, B1 => n3843, B2 => 
                           n60065, ZN => n11144);
   U10927 : OAI22_X1 port map( A1 => n60066, A2 => n62029, B1 => n3842, B2 => 
                           n60065, ZN => n11145);
   U10928 : OAI22_X1 port map( A1 => n60067, A2 => n62043, B1 => n3841, B2 => 
                           n60065, ZN => n11146);
   U10929 : OAI22_X1 port map( A1 => n60067, A2 => n62057, B1 => n3840, B2 => 
                           n60065, ZN => n11147);
   U10930 : OAI22_X1 port map( A1 => n60067, A2 => n62071, B1 => n3839, B2 => 
                           n60065, ZN => n11148);
   U10931 : OAI22_X1 port map( A1 => n60067, A2 => n62085, B1 => n3838, B2 => 
                           n60065, ZN => n11149);
   U10932 : OAI22_X1 port map( A1 => n60067, A2 => n62099, B1 => n3837, B2 => 
                           n60065, ZN => n11150);
   U10933 : OAI22_X1 port map( A1 => n60068, A2 => n62113, B1 => n3836, B2 => 
                           n60065, ZN => n11151);
   U10934 : OAI22_X1 port map( A1 => n60068, A2 => n60966, B1 => n3835, B2 => 
                           n60065, ZN => n11152);
   U10935 : OAI22_X1 port map( A1 => n60068, A2 => n60980, B1 => n3834, B2 => 
                           n15233, ZN => n11153);
   U10936 : OAI22_X1 port map( A1 => n60068, A2 => n60994, B1 => n3833, B2 => 
                           n15233, ZN => n11154);
   U10937 : OAI22_X1 port map( A1 => n60068, A2 => n61008, B1 => n3832, B2 => 
                           n15233, ZN => n11155);
   U10938 : OAI22_X1 port map( A1 => n60069, A2 => n61022, B1 => n3831, B2 => 
                           n15233, ZN => n11156);
   U10939 : OAI22_X1 port map( A1 => n60069, A2 => n61036, B1 => n3830, B2 => 
                           n15233, ZN => n11157);
   U10940 : OAI22_X1 port map( A1 => n60069, A2 => n61050, B1 => n3829, B2 => 
                           n15233, ZN => n11158);
   U10941 : OAI22_X1 port map( A1 => n60069, A2 => n61064, B1 => n3828, B2 => 
                           n15233, ZN => n11159);
   U10942 : OAI22_X1 port map( A1 => n60069, A2 => n61078, B1 => n3827, B2 => 
                           n60065, ZN => n11160);
   U10943 : OAI22_X1 port map( A1 => n60070, A2 => n61092, B1 => n3826, B2 => 
                           n60065, ZN => n11161);
   U10944 : OAI22_X1 port map( A1 => n60070, A2 => n61106, B1 => n3825, B2 => 
                           n60065, ZN => n11162);
   U10945 : OAI22_X1 port map( A1 => n60070, A2 => n61120, B1 => n3824, B2 => 
                           n60065, ZN => n11163);
   U10946 : OAI22_X1 port map( A1 => n60070, A2 => n61134, B1 => n3823, B2 => 
                           n60065, ZN => n11164);
   U10947 : OAI22_X1 port map( A1 => n60048, A2 => n61973, B1 => n3798, B2 => 
                           n60047, ZN => n11077);
   U10948 : OAI22_X1 port map( A1 => n60048, A2 => n61987, B1 => n3797, B2 => 
                           n60047, ZN => n11078);
   U10949 : OAI22_X1 port map( A1 => n60048, A2 => n62001, B1 => n3796, B2 => 
                           n60047, ZN => n11079);
   U10950 : OAI22_X1 port map( A1 => n60048, A2 => n62015, B1 => n3795, B2 => 
                           n60047, ZN => n11080);
   U10951 : OAI22_X1 port map( A1 => n60048, A2 => n62029, B1 => n3794, B2 => 
                           n60047, ZN => n11081);
   U10952 : OAI22_X1 port map( A1 => n60049, A2 => n62043, B1 => n3793, B2 => 
                           n60047, ZN => n11082);
   U10953 : OAI22_X1 port map( A1 => n60049, A2 => n62057, B1 => n3792, B2 => 
                           n60047, ZN => n11083);
   U10954 : OAI22_X1 port map( A1 => n60049, A2 => n62071, B1 => n3791, B2 => 
                           n60047, ZN => n11084);
   U10955 : OAI22_X1 port map( A1 => n60049, A2 => n62085, B1 => n3790, B2 => 
                           n60047, ZN => n11085);
   U10956 : OAI22_X1 port map( A1 => n60049, A2 => n62099, B1 => n3789, B2 => 
                           n60047, ZN => n11086);
   U10957 : OAI22_X1 port map( A1 => n60050, A2 => n62113, B1 => n3788, B2 => 
                           n60047, ZN => n11087);
   U10958 : OAI22_X1 port map( A1 => n60050, A2 => n60966, B1 => n3787, B2 => 
                           n60047, ZN => n11088);
   U10959 : OAI22_X1 port map( A1 => n60050, A2 => n60980, B1 => n3786, B2 => 
                           n15235, ZN => n11089);
   U10960 : OAI22_X1 port map( A1 => n60050, A2 => n60994, B1 => n3785, B2 => 
                           n15235, ZN => n11090);
   U10961 : OAI22_X1 port map( A1 => n60050, A2 => n61008, B1 => n3784, B2 => 
                           n15235, ZN => n11091);
   U10962 : OAI22_X1 port map( A1 => n60051, A2 => n61022, B1 => n3783, B2 => 
                           n15235, ZN => n11092);
   U10963 : OAI22_X1 port map( A1 => n60051, A2 => n61036, B1 => n3782, B2 => 
                           n15235, ZN => n11093);
   U10964 : OAI22_X1 port map( A1 => n60051, A2 => n61050, B1 => n3781, B2 => 
                           n15235, ZN => n11094);
   U10965 : OAI22_X1 port map( A1 => n60051, A2 => n61064, B1 => n3780, B2 => 
                           n15235, ZN => n11095);
   U10966 : OAI22_X1 port map( A1 => n60051, A2 => n61078, B1 => n3779, B2 => 
                           n60047, ZN => n11096);
   U10967 : OAI22_X1 port map( A1 => n60052, A2 => n61092, B1 => n3778, B2 => 
                           n60047, ZN => n11097);
   U10968 : OAI22_X1 port map( A1 => n60052, A2 => n61106, B1 => n3777, B2 => 
                           n60047, ZN => n11098);
   U10969 : OAI22_X1 port map( A1 => n60052, A2 => n61120, B1 => n3776, B2 => 
                           n60047, ZN => n11099);
   U10970 : OAI22_X1 port map( A1 => n60052, A2 => n61134, B1 => n3775, B2 => 
                           n60047, ZN => n11100);
   U10971 : OAI22_X1 port map( A1 => n60039, A2 => n61973, B1 => n3774, B2 => 
                           n60038, ZN => n11045);
   U10972 : OAI22_X1 port map( A1 => n60039, A2 => n61987, B1 => n3773, B2 => 
                           n60038, ZN => n11046);
   U10973 : OAI22_X1 port map( A1 => n60039, A2 => n62001, B1 => n3772, B2 => 
                           n60038, ZN => n11047);
   U10974 : OAI22_X1 port map( A1 => n60039, A2 => n62015, B1 => n3771, B2 => 
                           n60038, ZN => n11048);
   U10975 : OAI22_X1 port map( A1 => n60039, A2 => n62029, B1 => n3770, B2 => 
                           n60038, ZN => n11049);
   U10976 : OAI22_X1 port map( A1 => n60040, A2 => n62043, B1 => n3769, B2 => 
                           n60038, ZN => n11050);
   U10977 : OAI22_X1 port map( A1 => n60040, A2 => n62057, B1 => n3768, B2 => 
                           n60038, ZN => n11051);
   U10978 : OAI22_X1 port map( A1 => n60040, A2 => n62071, B1 => n3767, B2 => 
                           n60038, ZN => n11052);
   U10979 : OAI22_X1 port map( A1 => n60040, A2 => n62085, B1 => n3766, B2 => 
                           n60038, ZN => n11053);
   U10980 : OAI22_X1 port map( A1 => n60040, A2 => n62099, B1 => n3765, B2 => 
                           n60038, ZN => n11054);
   U10981 : OAI22_X1 port map( A1 => n60041, A2 => n62113, B1 => n3764, B2 => 
                           n60038, ZN => n11055);
   U10982 : OAI22_X1 port map( A1 => n60041, A2 => n60966, B1 => n3763, B2 => 
                           n60038, ZN => n11056);
   U10983 : OAI22_X1 port map( A1 => n60041, A2 => n60980, B1 => n3762, B2 => 
                           n15236, ZN => n11057);
   U10984 : OAI22_X1 port map( A1 => n60041, A2 => n60994, B1 => n3761, B2 => 
                           n15236, ZN => n11058);
   U10985 : OAI22_X1 port map( A1 => n60041, A2 => n61008, B1 => n3760, B2 => 
                           n15236, ZN => n11059);
   U10986 : OAI22_X1 port map( A1 => n60042, A2 => n61022, B1 => n3759, B2 => 
                           n15236, ZN => n11060);
   U10987 : OAI22_X1 port map( A1 => n60042, A2 => n61036, B1 => n3758, B2 => 
                           n15236, ZN => n11061);
   U10988 : OAI22_X1 port map( A1 => n60042, A2 => n61050, B1 => n3757, B2 => 
                           n15236, ZN => n11062);
   U10989 : OAI22_X1 port map( A1 => n60042, A2 => n61064, B1 => n3756, B2 => 
                           n15236, ZN => n11063);
   U10990 : OAI22_X1 port map( A1 => n60042, A2 => n61078, B1 => n3755, B2 => 
                           n60038, ZN => n11064);
   U10991 : OAI22_X1 port map( A1 => n60043, A2 => n61092, B1 => n3754, B2 => 
                           n60038, ZN => n11065);
   U10992 : OAI22_X1 port map( A1 => n60043, A2 => n61106, B1 => n3753, B2 => 
                           n60038, ZN => n11066);
   U10993 : OAI22_X1 port map( A1 => n60043, A2 => n61120, B1 => n3752, B2 => 
                           n60038, ZN => n11067);
   U10994 : OAI22_X1 port map( A1 => n60043, A2 => n61134, B1 => n3751, B2 => 
                           n60038, ZN => n11068);
   U10995 : OAI22_X1 port map( A1 => n60030, A2 => n61973, B1 => n3750, B2 => 
                           n60029, ZN => n11013);
   U10996 : OAI22_X1 port map( A1 => n60030, A2 => n61987, B1 => n3749, B2 => 
                           n60029, ZN => n11014);
   U10997 : OAI22_X1 port map( A1 => n60030, A2 => n62001, B1 => n3748, B2 => 
                           n60029, ZN => n11015);
   U10998 : OAI22_X1 port map( A1 => n60030, A2 => n62015, B1 => n3747, B2 => 
                           n60029, ZN => n11016);
   U10999 : OAI22_X1 port map( A1 => n60030, A2 => n62029, B1 => n3746, B2 => 
                           n60029, ZN => n11017);
   U11000 : OAI22_X1 port map( A1 => n60031, A2 => n62043, B1 => n3745, B2 => 
                           n60029, ZN => n11018);
   U11001 : OAI22_X1 port map( A1 => n60031, A2 => n62057, B1 => n3744, B2 => 
                           n60029, ZN => n11019);
   U11002 : OAI22_X1 port map( A1 => n60031, A2 => n62071, B1 => n3743, B2 => 
                           n60029, ZN => n11020);
   U11003 : OAI22_X1 port map( A1 => n60031, A2 => n62085, B1 => n3742, B2 => 
                           n60029, ZN => n11021);
   U11004 : OAI22_X1 port map( A1 => n60031, A2 => n62099, B1 => n3741, B2 => 
                           n60029, ZN => n11022);
   U11005 : OAI22_X1 port map( A1 => n60032, A2 => n62113, B1 => n3740, B2 => 
                           n60029, ZN => n11023);
   U11006 : OAI22_X1 port map( A1 => n60032, A2 => n60966, B1 => n3739, B2 => 
                           n60029, ZN => n11024);
   U11007 : OAI22_X1 port map( A1 => n60032, A2 => n60980, B1 => n3738, B2 => 
                           n15237, ZN => n11025);
   U11008 : OAI22_X1 port map( A1 => n60032, A2 => n60994, B1 => n3737, B2 => 
                           n15237, ZN => n11026);
   U11009 : OAI22_X1 port map( A1 => n60032, A2 => n61008, B1 => n3736, B2 => 
                           n15237, ZN => n11027);
   U11010 : OAI22_X1 port map( A1 => n60033, A2 => n61022, B1 => n3735, B2 => 
                           n15237, ZN => n11028);
   U11011 : OAI22_X1 port map( A1 => n60033, A2 => n61036, B1 => n3734, B2 => 
                           n15237, ZN => n11029);
   U11012 : OAI22_X1 port map( A1 => n60033, A2 => n61050, B1 => n3733, B2 => 
                           n15237, ZN => n11030);
   U11013 : OAI22_X1 port map( A1 => n60033, A2 => n61064, B1 => n3732, B2 => 
                           n15237, ZN => n11031);
   U11014 : OAI22_X1 port map( A1 => n60033, A2 => n61078, B1 => n3731, B2 => 
                           n60029, ZN => n11032);
   U11015 : OAI22_X1 port map( A1 => n60034, A2 => n61092, B1 => n3730, B2 => 
                           n60029, ZN => n11033);
   U11016 : OAI22_X1 port map( A1 => n60034, A2 => n61106, B1 => n3729, B2 => 
                           n60029, ZN => n11034);
   U11017 : OAI22_X1 port map( A1 => n60034, A2 => n61120, B1 => n3728, B2 => 
                           n60029, ZN => n11035);
   U11018 : OAI22_X1 port map( A1 => n60034, A2 => n61134, B1 => n3727, B2 => 
                           n60029, ZN => n11036);
   U11019 : OAI22_X1 port map( A1 => n60003, A2 => n61973, B1 => n3678, B2 => 
                           n60002, ZN => n10917);
   U11020 : OAI22_X1 port map( A1 => n60003, A2 => n61987, B1 => n3677, B2 => 
                           n60002, ZN => n10918);
   U11021 : OAI22_X1 port map( A1 => n60003, A2 => n62001, B1 => n3676, B2 => 
                           n60002, ZN => n10919);
   U11022 : OAI22_X1 port map( A1 => n60003, A2 => n62015, B1 => n3675, B2 => 
                           n60002, ZN => n10920);
   U11023 : OAI22_X1 port map( A1 => n60003, A2 => n62029, B1 => n3674, B2 => 
                           n60002, ZN => n10921);
   U11024 : OAI22_X1 port map( A1 => n60004, A2 => n62043, B1 => n3673, B2 => 
                           n60002, ZN => n10922);
   U11025 : OAI22_X1 port map( A1 => n60004, A2 => n62057, B1 => n3672, B2 => 
                           n60002, ZN => n10923);
   U11026 : OAI22_X1 port map( A1 => n60004, A2 => n62071, B1 => n3671, B2 => 
                           n60002, ZN => n10924);
   U11027 : OAI22_X1 port map( A1 => n60004, A2 => n62085, B1 => n3670, B2 => 
                           n60002, ZN => n10925);
   U11028 : OAI22_X1 port map( A1 => n60004, A2 => n62099, B1 => n3669, B2 => 
                           n60002, ZN => n10926);
   U11029 : OAI22_X1 port map( A1 => n60005, A2 => n62113, B1 => n3668, B2 => 
                           n60002, ZN => n10927);
   U11030 : OAI22_X1 port map( A1 => n60005, A2 => n60966, B1 => n3667, B2 => 
                           n60002, ZN => n10928);
   U11031 : OAI22_X1 port map( A1 => n60005, A2 => n60980, B1 => n3666, B2 => 
                           n15240, ZN => n10929);
   U11032 : OAI22_X1 port map( A1 => n60005, A2 => n60994, B1 => n3665, B2 => 
                           n15240, ZN => n10930);
   U11033 : OAI22_X1 port map( A1 => n60005, A2 => n61008, B1 => n3664, B2 => 
                           n15240, ZN => n10931);
   U11034 : OAI22_X1 port map( A1 => n60006, A2 => n61022, B1 => n3663, B2 => 
                           n15240, ZN => n10932);
   U11035 : OAI22_X1 port map( A1 => n60006, A2 => n61036, B1 => n3662, B2 => 
                           n15240, ZN => n10933);
   U11036 : OAI22_X1 port map( A1 => n60006, A2 => n61050, B1 => n3661, B2 => 
                           n15240, ZN => n10934);
   U11037 : OAI22_X1 port map( A1 => n60006, A2 => n61064, B1 => n3660, B2 => 
                           n15240, ZN => n10935);
   U11038 : OAI22_X1 port map( A1 => n60006, A2 => n61078, B1 => n3659, B2 => 
                           n60002, ZN => n10936);
   U11039 : OAI22_X1 port map( A1 => n60007, A2 => n61092, B1 => n3658, B2 => 
                           n60002, ZN => n10937);
   U11040 : OAI22_X1 port map( A1 => n60007, A2 => n61106, B1 => n3657, B2 => 
                           n60002, ZN => n10938);
   U11041 : OAI22_X1 port map( A1 => n60007, A2 => n61120, B1 => n3656, B2 => 
                           n60002, ZN => n10939);
   U11042 : OAI22_X1 port map( A1 => n60007, A2 => n61134, B1 => n3655, B2 => 
                           n60002, ZN => n10940);
   U11043 : OAI22_X1 port map( A1 => n59994, A2 => n61974, B1 => n3654, B2 => 
                           n59993, ZN => n10885);
   U11044 : OAI22_X1 port map( A1 => n59994, A2 => n61988, B1 => n3653, B2 => 
                           n59993, ZN => n10886);
   U11045 : OAI22_X1 port map( A1 => n59994, A2 => n62002, B1 => n3652, B2 => 
                           n59993, ZN => n10887);
   U11046 : OAI22_X1 port map( A1 => n59994, A2 => n62016, B1 => n3651, B2 => 
                           n59993, ZN => n10888);
   U11047 : OAI22_X1 port map( A1 => n59994, A2 => n62030, B1 => n3650, B2 => 
                           n59993, ZN => n10889);
   U11048 : OAI22_X1 port map( A1 => n59995, A2 => n62044, B1 => n3649, B2 => 
                           n59993, ZN => n10890);
   U11049 : OAI22_X1 port map( A1 => n59996, A2 => n60980, B1 => n3648, B2 => 
                           n15241, ZN => n10897);
   U11050 : OAI22_X1 port map( A1 => n59996, A2 => n60994, B1 => n3647, B2 => 
                           n15241, ZN => n10898);
   U11051 : OAI22_X1 port map( A1 => n59996, A2 => n61008, B1 => n3646, B2 => 
                           n15241, ZN => n10899);
   U11052 : OAI22_X1 port map( A1 => n59997, A2 => n61022, B1 => n3645, B2 => 
                           n59993, ZN => n10900);
   U11053 : OAI22_X1 port map( A1 => n59997, A2 => n61036, B1 => n3620, B2 => 
                           n59993, ZN => n10901);
   U11054 : OAI22_X1 port map( A1 => n59997, A2 => n61050, B1 => n3619, B2 => 
                           n59993, ZN => n10902);
   U11055 : OAI22_X1 port map( A1 => n59997, A2 => n61064, B1 => n3618, B2 => 
                           n59993, ZN => n10903);
   U11056 : OAI22_X1 port map( A1 => n59997, A2 => n61078, B1 => n3617, B2 => 
                           n59993, ZN => n10904);
   U11057 : OAI22_X1 port map( A1 => n59985, A2 => n61973, B1 => n3990, B2 => 
                           n59984, ZN => n10853);
   U11058 : OAI22_X1 port map( A1 => n59985, A2 => n61987, B1 => n3989, B2 => 
                           n59984, ZN => n10854);
   U11059 : OAI22_X1 port map( A1 => n59985, A2 => n62001, B1 => n3988, B2 => 
                           n59984, ZN => n10855);
   U11060 : OAI22_X1 port map( A1 => n59985, A2 => n62015, B1 => n3987, B2 => 
                           n59984, ZN => n10856);
   U11061 : OAI22_X1 port map( A1 => n59985, A2 => n62029, B1 => n3986, B2 => 
                           n59984, ZN => n10857);
   U11062 : OAI22_X1 port map( A1 => n59986, A2 => n62043, B1 => n3985, B2 => 
                           n59984, ZN => n10858);
   U11063 : OAI22_X1 port map( A1 => n59986, A2 => n62057, B1 => n3984, B2 => 
                           n59984, ZN => n10859);
   U11064 : OAI22_X1 port map( A1 => n59986, A2 => n62071, B1 => n3983, B2 => 
                           n59984, ZN => n10860);
   U11065 : OAI22_X1 port map( A1 => n59986, A2 => n62085, B1 => n3982, B2 => 
                           n59984, ZN => n10861);
   U11066 : OAI22_X1 port map( A1 => n59986, A2 => n62099, B1 => n3981, B2 => 
                           n59984, ZN => n10862);
   U11067 : OAI22_X1 port map( A1 => n59987, A2 => n62113, B1 => n3980, B2 => 
                           n59984, ZN => n10863);
   U11068 : OAI22_X1 port map( A1 => n59987, A2 => n60967, B1 => n3979, B2 => 
                           n59984, ZN => n10864);
   U11069 : OAI22_X1 port map( A1 => n59987, A2 => n60981, B1 => n3978, B2 => 
                           n15242, ZN => n10865);
   U11070 : OAI22_X1 port map( A1 => n59987, A2 => n60995, B1 => n3977, B2 => 
                           n15242, ZN => n10866);
   U11071 : OAI22_X1 port map( A1 => n59987, A2 => n61009, B1 => n3976, B2 => 
                           n15242, ZN => n10867);
   U11072 : OAI22_X1 port map( A1 => n59988, A2 => n61023, B1 => n3975, B2 => 
                           n15242, ZN => n10868);
   U11073 : OAI22_X1 port map( A1 => n59988, A2 => n61037, B1 => n3974, B2 => 
                           n15242, ZN => n10869);
   U11074 : OAI22_X1 port map( A1 => n59988, A2 => n61051, B1 => n3973, B2 => 
                           n15242, ZN => n10870);
   U11075 : OAI22_X1 port map( A1 => n59988, A2 => n61065, B1 => n3972, B2 => 
                           n15242, ZN => n10871);
   U11076 : OAI22_X1 port map( A1 => n59988, A2 => n61079, B1 => n3971, B2 => 
                           n59984, ZN => n10872);
   U11077 : OAI22_X1 port map( A1 => n59989, A2 => n61093, B1 => n3970, B2 => 
                           n59984, ZN => n10873);
   U11078 : OAI22_X1 port map( A1 => n59989, A2 => n61107, B1 => n3969, B2 => 
                           n59984, ZN => n10874);
   U11079 : OAI22_X1 port map( A1 => n59989, A2 => n61121, B1 => n3968, B2 => 
                           n59984, ZN => n10875);
   U11080 : OAI22_X1 port map( A1 => n59989, A2 => n61135, B1 => n3967, B2 => 
                           n59984, ZN => n10876);
   U11081 : OAI22_X1 port map( A1 => n59967, A2 => n62030, B1 => n3616, B2 => 
                           n59966, ZN => n10793);
   U11082 : OAI22_X1 port map( A1 => n59968, A2 => n62044, B1 => n3615, B2 => 
                           n59966, ZN => n10794);
   U11083 : OAI22_X1 port map( A1 => n59968, A2 => n62058, B1 => n3614, B2 => 
                           n59966, ZN => n10795);
   U11084 : OAI22_X1 port map( A1 => n59968, A2 => n62072, B1 => n3613, B2 => 
                           n59966, ZN => n10796);
   U11085 : OAI22_X1 port map( A1 => n59968, A2 => n62086, B1 => n3612, B2 => 
                           n59966, ZN => n10797);
   U11086 : OAI22_X1 port map( A1 => n59968, A2 => n62100, B1 => n3611, B2 => 
                           n59966, ZN => n10798);
   U11087 : OAI22_X1 port map( A1 => n59969, A2 => n62114, B1 => n3610, B2 => 
                           n59966, ZN => n10799);
   U11088 : OAI22_X1 port map( A1 => n59969, A2 => n60967, B1 => n3609, B2 => 
                           n59966, ZN => n10800);
   U11089 : OAI22_X1 port map( A1 => n59969, A2 => n60981, B1 => n3608, B2 => 
                           n15244, ZN => n10801);
   U11090 : OAI22_X1 port map( A1 => n59969, A2 => n60995, B1 => n3607, B2 => 
                           n15244, ZN => n10802);
   U11091 : OAI22_X1 port map( A1 => n59969, A2 => n61009, B1 => n3606, B2 => 
                           n15244, ZN => n10803);
   U11092 : OAI22_X1 port map( A1 => n59970, A2 => n61023, B1 => n3605, B2 => 
                           n15244, ZN => n10804);
   U11093 : OAI22_X1 port map( A1 => n59970, A2 => n61037, B1 => n3604, B2 => 
                           n15244, ZN => n10805);
   U11094 : OAI22_X1 port map( A1 => n59970, A2 => n61051, B1 => n3603, B2 => 
                           n15244, ZN => n10806);
   U11095 : OAI22_X1 port map( A1 => n59970, A2 => n61065, B1 => n3602, B2 => 
                           n15244, ZN => n10807);
   U11096 : OAI22_X1 port map( A1 => n59970, A2 => n61079, B1 => n3601, B2 => 
                           n59966, ZN => n10808);
   U11097 : OAI22_X1 port map( A1 => n59971, A2 => n61093, B1 => n3600, B2 => 
                           n59966, ZN => n10809);
   U11098 : OAI22_X1 port map( A1 => n59971, A2 => n61107, B1 => n3599, B2 => 
                           n59966, ZN => n10810);
   U11099 : OAI22_X1 port map( A1 => n59971, A2 => n61121, B1 => n3598, B2 => 
                           n59966, ZN => n10811);
   U11100 : OAI22_X1 port map( A1 => n59971, A2 => n61135, B1 => n3597, B2 => 
                           n59966, ZN => n10812);
   U11101 : OAI22_X1 port map( A1 => n59913, A2 => n61974, B1 => n3500, B2 => 
                           n59912, ZN => n10597);
   U11102 : OAI22_X1 port map( A1 => n59913, A2 => n61988, B1 => n3499, B2 => 
                           n59912, ZN => n10598);
   U11103 : OAI22_X1 port map( A1 => n59913, A2 => n62002, B1 => n3498, B2 => 
                           n59912, ZN => n10599);
   U11104 : OAI22_X1 port map( A1 => n59913, A2 => n62016, B1 => n3497, B2 => 
                           n59912, ZN => n10600);
   U11105 : OAI22_X1 port map( A1 => n59913, A2 => n62030, B1 => n3496, B2 => 
                           n59912, ZN => n10601);
   U11106 : OAI22_X1 port map( A1 => n59914, A2 => n62044, B1 => n3495, B2 => 
                           n59912, ZN => n10602);
   U11107 : OAI22_X1 port map( A1 => n59914, A2 => n62058, B1 => n3494, B2 => 
                           n59912, ZN => n10603);
   U11108 : OAI22_X1 port map( A1 => n59914, A2 => n62072, B1 => n3493, B2 => 
                           n59912, ZN => n10604);
   U11109 : OAI22_X1 port map( A1 => n59914, A2 => n62086, B1 => n3492, B2 => 
                           n59912, ZN => n10605);
   U11110 : OAI22_X1 port map( A1 => n59914, A2 => n62100, B1 => n3491, B2 => 
                           n59912, ZN => n10606);
   U11111 : OAI22_X1 port map( A1 => n59915, A2 => n62114, B1 => n3490, B2 => 
                           n59912, ZN => n10607);
   U11112 : OAI22_X1 port map( A1 => n59915, A2 => n60967, B1 => n3489, B2 => 
                           n59912, ZN => n10608);
   U11113 : OAI22_X1 port map( A1 => n59915, A2 => n60981, B1 => n3488, B2 => 
                           n15251, ZN => n10609);
   U11114 : OAI22_X1 port map( A1 => n59915, A2 => n60995, B1 => n3487, B2 => 
                           n15251, ZN => n10610);
   U11115 : OAI22_X1 port map( A1 => n59915, A2 => n61009, B1 => n3486, B2 => 
                           n15251, ZN => n10611);
   U11116 : OAI22_X1 port map( A1 => n59916, A2 => n61023, B1 => n3485, B2 => 
                           n15251, ZN => n10612);
   U11117 : OAI22_X1 port map( A1 => n59916, A2 => n61037, B1 => n3484, B2 => 
                           n15251, ZN => n10613);
   U11118 : OAI22_X1 port map( A1 => n59916, A2 => n61051, B1 => n3483, B2 => 
                           n15251, ZN => n10614);
   U11119 : OAI22_X1 port map( A1 => n59916, A2 => n61065, B1 => n3482, B2 => 
                           n15251, ZN => n10615);
   U11120 : OAI22_X1 port map( A1 => n59916, A2 => n61079, B1 => n3481, B2 => 
                           n59912, ZN => n10616);
   U11121 : OAI22_X1 port map( A1 => n59917, A2 => n61093, B1 => n3480, B2 => 
                           n59912, ZN => n10617);
   U11122 : OAI22_X1 port map( A1 => n59917, A2 => n61107, B1 => n3479, B2 => 
                           n59912, ZN => n10618);
   U11123 : OAI22_X1 port map( A1 => n59917, A2 => n61121, B1 => n3478, B2 => 
                           n59912, ZN => n10619);
   U11124 : OAI22_X1 port map( A1 => n59917, A2 => n61135, B1 => n3477, B2 => 
                           n59912, ZN => n10620);
   U11125 : OAI22_X1 port map( A1 => n59904, A2 => n61974, B1 => n3476, B2 => 
                           n59903, ZN => n10565);
   U11126 : OAI22_X1 port map( A1 => n59904, A2 => n61988, B1 => n3475, B2 => 
                           n59903, ZN => n10566);
   U11127 : OAI22_X1 port map( A1 => n59904, A2 => n62002, B1 => n3474, B2 => 
                           n59903, ZN => n10567);
   U11128 : OAI22_X1 port map( A1 => n59904, A2 => n62016, B1 => n3473, B2 => 
                           n59903, ZN => n10568);
   U11129 : OAI22_X1 port map( A1 => n59904, A2 => n62030, B1 => n3472, B2 => 
                           n59903, ZN => n10569);
   U11130 : OAI22_X1 port map( A1 => n59905, A2 => n62044, B1 => n3471, B2 => 
                           n59903, ZN => n10570);
   U11131 : OAI22_X1 port map( A1 => n59905, A2 => n62058, B1 => n3470, B2 => 
                           n59903, ZN => n10571);
   U11132 : OAI22_X1 port map( A1 => n59905, A2 => n62072, B1 => n3469, B2 => 
                           n59903, ZN => n10572);
   U11133 : OAI22_X1 port map( A1 => n59905, A2 => n62086, B1 => n3468, B2 => 
                           n59903, ZN => n10573);
   U11134 : OAI22_X1 port map( A1 => n59905, A2 => n62100, B1 => n3467, B2 => 
                           n59903, ZN => n10574);
   U11135 : OAI22_X1 port map( A1 => n59906, A2 => n62114, B1 => n3466, B2 => 
                           n59903, ZN => n10575);
   U11136 : OAI22_X1 port map( A1 => n59906, A2 => n60967, B1 => n3465, B2 => 
                           n59903, ZN => n10576);
   U11137 : OAI22_X1 port map( A1 => n59906, A2 => n60981, B1 => n3464, B2 => 
                           n15252, ZN => n10577);
   U11138 : OAI22_X1 port map( A1 => n59906, A2 => n60995, B1 => n3463, B2 => 
                           n15252, ZN => n10578);
   U11139 : OAI22_X1 port map( A1 => n59906, A2 => n61009, B1 => n3462, B2 => 
                           n15252, ZN => n10579);
   U11140 : OAI22_X1 port map( A1 => n59907, A2 => n61023, B1 => n3461, B2 => 
                           n15252, ZN => n10580);
   U11141 : OAI22_X1 port map( A1 => n59907, A2 => n61037, B1 => n3460, B2 => 
                           n15252, ZN => n10581);
   U11142 : OAI22_X1 port map( A1 => n59907, A2 => n61051, B1 => n3459, B2 => 
                           n15252, ZN => n10582);
   U11143 : OAI22_X1 port map( A1 => n59907, A2 => n61065, B1 => n3458, B2 => 
                           n15252, ZN => n10583);
   U11144 : OAI22_X1 port map( A1 => n59907, A2 => n61079, B1 => n3457, B2 => 
                           n59903, ZN => n10584);
   U11145 : OAI22_X1 port map( A1 => n59908, A2 => n61093, B1 => n3408, B2 => 
                           n59903, ZN => n10585);
   U11146 : OAI22_X1 port map( A1 => n59908, A2 => n61107, B1 => n3407, B2 => 
                           n59903, ZN => n10586);
   U11147 : OAI22_X1 port map( A1 => n59908, A2 => n61121, B1 => n3406, B2 => 
                           n59903, ZN => n10587);
   U11148 : OAI22_X1 port map( A1 => n59908, A2 => n61135, B1 => n3405, B2 => 
                           n59903, ZN => n10588);
   U11149 : OAI22_X1 port map( A1 => n59895, A2 => n61974, B1 => n3404, B2 => 
                           n59894, ZN => n10533);
   U11150 : OAI22_X1 port map( A1 => n59895, A2 => n61988, B1 => n3403, B2 => 
                           n59894, ZN => n10534);
   U11151 : OAI22_X1 port map( A1 => n59895, A2 => n62002, B1 => n3402, B2 => 
                           n59894, ZN => n10535);
   U11152 : OAI22_X1 port map( A1 => n59895, A2 => n62016, B1 => n3401, B2 => 
                           n59894, ZN => n10536);
   U11153 : OAI22_X1 port map( A1 => n59895, A2 => n62030, B1 => n3400, B2 => 
                           n59894, ZN => n10537);
   U11154 : OAI22_X1 port map( A1 => n59896, A2 => n62044, B1 => n3399, B2 => 
                           n59894, ZN => n10538);
   U11155 : OAI22_X1 port map( A1 => n59896, A2 => n62058, B1 => n3398, B2 => 
                           n59894, ZN => n10539);
   U11156 : OAI22_X1 port map( A1 => n59896, A2 => n62072, B1 => n3397, B2 => 
                           n59894, ZN => n10540);
   U11157 : OAI22_X1 port map( A1 => n59896, A2 => n62086, B1 => n3396, B2 => 
                           n59894, ZN => n10541);
   U11158 : OAI22_X1 port map( A1 => n59896, A2 => n62100, B1 => n3395, B2 => 
                           n59894, ZN => n10542);
   U11159 : OAI22_X1 port map( A1 => n59897, A2 => n62114, B1 => n3394, B2 => 
                           n59894, ZN => n10543);
   U11160 : OAI22_X1 port map( A1 => n59897, A2 => n60967, B1 => n3393, B2 => 
                           n59894, ZN => n10544);
   U11161 : OAI22_X1 port map( A1 => n59897, A2 => n60981, B1 => n3392, B2 => 
                           n15253, ZN => n10545);
   U11162 : OAI22_X1 port map( A1 => n59897, A2 => n60995, B1 => n3391, B2 => 
                           n15253, ZN => n10546);
   U11163 : OAI22_X1 port map( A1 => n59897, A2 => n61009, B1 => n3390, B2 => 
                           n15253, ZN => n10547);
   U11164 : OAI22_X1 port map( A1 => n59898, A2 => n61023, B1 => n3389, B2 => 
                           n15253, ZN => n10548);
   U11165 : OAI22_X1 port map( A1 => n59898, A2 => n61037, B1 => n3388, B2 => 
                           n15253, ZN => n10549);
   U11166 : OAI22_X1 port map( A1 => n59898, A2 => n61051, B1 => n3387, B2 => 
                           n15253, ZN => n10550);
   U11167 : OAI22_X1 port map( A1 => n59898, A2 => n61065, B1 => n3386, B2 => 
                           n15253, ZN => n10551);
   U11168 : OAI22_X1 port map( A1 => n59898, A2 => n61079, B1 => n3385, B2 => 
                           n59894, ZN => n10552);
   U11169 : OAI22_X1 port map( A1 => n59899, A2 => n61093, B1 => n3384, B2 => 
                           n59894, ZN => n10553);
   U11170 : OAI22_X1 port map( A1 => n59899, A2 => n61107, B1 => n3383, B2 => 
                           n59894, ZN => n10554);
   U11171 : OAI22_X1 port map( A1 => n59899, A2 => n61121, B1 => n3382, B2 => 
                           n59894, ZN => n10555);
   U11172 : OAI22_X1 port map( A1 => n59899, A2 => n61135, B1 => n3381, B2 => 
                           n59894, ZN => n10556);
   U11173 : OAI22_X1 port map( A1 => n59886, A2 => n61975, B1 => n2390, B2 => 
                           n59885, ZN => n10501);
   U11174 : OAI22_X1 port map( A1 => n59886, A2 => n61989, B1 => n2389, B2 => 
                           n59885, ZN => n10502);
   U11175 : OAI22_X1 port map( A1 => n59886, A2 => n62003, B1 => n2388, B2 => 
                           n59885, ZN => n10503);
   U11176 : OAI22_X1 port map( A1 => n59886, A2 => n62017, B1 => n2387, B2 => 
                           n59885, ZN => n10504);
   U11177 : OAI22_X1 port map( A1 => n59886, A2 => n62031, B1 => n2386, B2 => 
                           n59885, ZN => n10505);
   U11178 : OAI22_X1 port map( A1 => n59887, A2 => n62045, B1 => n2385, B2 => 
                           n59885, ZN => n10506);
   U11179 : OAI22_X1 port map( A1 => n59887, A2 => n62059, B1 => n2384, B2 => 
                           n59885, ZN => n10507);
   U11180 : OAI22_X1 port map( A1 => n59887, A2 => n62073, B1 => n2383, B2 => 
                           n59885, ZN => n10508);
   U11181 : OAI22_X1 port map( A1 => n59887, A2 => n62087, B1 => n2382, B2 => 
                           n59885, ZN => n10509);
   U11182 : OAI22_X1 port map( A1 => n59887, A2 => n62101, B1 => n2381, B2 => 
                           n59885, ZN => n10510);
   U11183 : OAI22_X1 port map( A1 => n59888, A2 => n62115, B1 => n2380, B2 => 
                           n59885, ZN => n10511);
   U11184 : OAI22_X1 port map( A1 => n59888, A2 => n60967, B1 => n2379, B2 => 
                           n59885, ZN => n10512);
   U11185 : OAI22_X1 port map( A1 => n59888, A2 => n60981, B1 => n2378, B2 => 
                           n15254, ZN => n10513);
   U11186 : OAI22_X1 port map( A1 => n59888, A2 => n60995, B1 => n2377, B2 => 
                           n15254, ZN => n10514);
   U11187 : OAI22_X1 port map( A1 => n59888, A2 => n61009, B1 => n2376, B2 => 
                           n15254, ZN => n10515);
   U11188 : OAI22_X1 port map( A1 => n59889, A2 => n61023, B1 => n2375, B2 => 
                           n15254, ZN => n10516);
   U11189 : OAI22_X1 port map( A1 => n59889, A2 => n61037, B1 => n2374, B2 => 
                           n15254, ZN => n10517);
   U11190 : OAI22_X1 port map( A1 => n59889, A2 => n61051, B1 => n2373, B2 => 
                           n15254, ZN => n10518);
   U11191 : OAI22_X1 port map( A1 => n59889, A2 => n61065, B1 => n2372, B2 => 
                           n15254, ZN => n10519);
   U11192 : OAI22_X1 port map( A1 => n59889, A2 => n61079, B1 => n2371, B2 => 
                           n59885, ZN => n10520);
   U11193 : OAI22_X1 port map( A1 => n59890, A2 => n61093, B1 => n2370, B2 => 
                           n59885, ZN => n10521);
   U11194 : OAI22_X1 port map( A1 => n59890, A2 => n61107, B1 => n2369, B2 => 
                           n59885, ZN => n10522);
   U11195 : OAI22_X1 port map( A1 => n59890, A2 => n61121, B1 => n2368, B2 => 
                           n59885, ZN => n10523);
   U11196 : OAI22_X1 port map( A1 => n59890, A2 => n61135, B1 => n2367, B2 => 
                           n59885, ZN => n10524);
   U11197 : OAI22_X1 port map( A1 => n59877, A2 => n61974, B1 => n2366, B2 => 
                           n59876, ZN => n10469);
   U11198 : OAI22_X1 port map( A1 => n59877, A2 => n61988, B1 => n2365, B2 => 
                           n59876, ZN => n10470);
   U11199 : OAI22_X1 port map( A1 => n59877, A2 => n62002, B1 => n2364, B2 => 
                           n59876, ZN => n10471);
   U11200 : OAI22_X1 port map( A1 => n59877, A2 => n62016, B1 => n2363, B2 => 
                           n59876, ZN => n10472);
   U11201 : OAI22_X1 port map( A1 => n59877, A2 => n62030, B1 => n2362, B2 => 
                           n59876, ZN => n10473);
   U11202 : OAI22_X1 port map( A1 => n59878, A2 => n62044, B1 => n2361, B2 => 
                           n59876, ZN => n10474);
   U11203 : OAI22_X1 port map( A1 => n59878, A2 => n62058, B1 => n2360, B2 => 
                           n59876, ZN => n10475);
   U11204 : OAI22_X1 port map( A1 => n59878, A2 => n62072, B1 => n2359, B2 => 
                           n59876, ZN => n10476);
   U11205 : OAI22_X1 port map( A1 => n59878, A2 => n62086, B1 => n2358, B2 => 
                           n59876, ZN => n10477);
   U11206 : OAI22_X1 port map( A1 => n59878, A2 => n62100, B1 => n2357, B2 => 
                           n59876, ZN => n10478);
   U11207 : OAI22_X1 port map( A1 => n59879, A2 => n62114, B1 => n2356, B2 => 
                           n59876, ZN => n10479);
   U11208 : OAI22_X1 port map( A1 => n59879, A2 => n60968, B1 => n2355, B2 => 
                           n59876, ZN => n10480);
   U11209 : OAI22_X1 port map( A1 => n59879, A2 => n60982, B1 => n2354, B2 => 
                           n15255, ZN => n10481);
   U11210 : OAI22_X1 port map( A1 => n59879, A2 => n60996, B1 => n2353, B2 => 
                           n15255, ZN => n10482);
   U11211 : OAI22_X1 port map( A1 => n59879, A2 => n61010, B1 => n2352, B2 => 
                           n15255, ZN => n10483);
   U11212 : OAI22_X1 port map( A1 => n59880, A2 => n61024, B1 => n2351, B2 => 
                           n15255, ZN => n10484);
   U11213 : OAI22_X1 port map( A1 => n59880, A2 => n61038, B1 => n2350, B2 => 
                           n15255, ZN => n10485);
   U11214 : OAI22_X1 port map( A1 => n59880, A2 => n61052, B1 => n2349, B2 => 
                           n15255, ZN => n10486);
   U11215 : OAI22_X1 port map( A1 => n59880, A2 => n61066, B1 => n2348, B2 => 
                           n15255, ZN => n10487);
   U11216 : OAI22_X1 port map( A1 => n59880, A2 => n61080, B1 => n2347, B2 => 
                           n59876, ZN => n10488);
   U11217 : OAI22_X1 port map( A1 => n59881, A2 => n61094, B1 => n2346, B2 => 
                           n59876, ZN => n10489);
   U11218 : OAI22_X1 port map( A1 => n59881, A2 => n61108, B1 => n2345, B2 => 
                           n59876, ZN => n10490);
   U11219 : OAI22_X1 port map( A1 => n59881, A2 => n61122, B1 => n2344, B2 => 
                           n59876, ZN => n10491);
   U11220 : OAI22_X1 port map( A1 => n59881, A2 => n61136, B1 => n2343, B2 => 
                           n59876, ZN => n10492);
   U11221 : OAI22_X1 port map( A1 => n59827, A2 => n61094, B1 => n3284, B2 => 
                           n59822, ZN => n10297);
   U11222 : OAI22_X1 port map( A1 => n59827, A2 => n61108, B1 => n3283, B2 => 
                           n59822, ZN => n10298);
   U11223 : OAI22_X1 port map( A1 => n59827, A2 => n61122, B1 => n3282, B2 => 
                           n59822, ZN => n10299);
   U11224 : OAI22_X1 port map( A1 => n59827, A2 => n61136, B1 => n3281, B2 => 
                           n59822, ZN => n10300);
   U11225 : OAI22_X1 port map( A1 => n59814, A2 => n61975, B1 => n3280, B2 => 
                           n59813, ZN => n10245);
   U11226 : OAI22_X1 port map( A1 => n59814, A2 => n61989, B1 => n3279, B2 => 
                           n59813, ZN => n10246);
   U11227 : OAI22_X1 port map( A1 => n59814, A2 => n62003, B1 => n3278, B2 => 
                           n59813, ZN => n10247);
   U11228 : OAI22_X1 port map( A1 => n59814, A2 => n62017, B1 => n3277, B2 => 
                           n59813, ZN => n10248);
   U11229 : OAI22_X1 port map( A1 => n59814, A2 => n62031, B1 => n3276, B2 => 
                           n59813, ZN => n10249);
   U11230 : OAI22_X1 port map( A1 => n59815, A2 => n62045, B1 => n3275, B2 => 
                           n59813, ZN => n10250);
   U11231 : OAI22_X1 port map( A1 => n59815, A2 => n62059, B1 => n3274, B2 => 
                           n59813, ZN => n10251);
   U11232 : OAI22_X1 port map( A1 => n59815, A2 => n62073, B1 => n3273, B2 => 
                           n59813, ZN => n10252);
   U11233 : OAI22_X1 port map( A1 => n59815, A2 => n62087, B1 => n3272, B2 => 
                           n59813, ZN => n10253);
   U11234 : OAI22_X1 port map( A1 => n59815, A2 => n62101, B1 => n3271, B2 => 
                           n59813, ZN => n10254);
   U11235 : OAI22_X1 port map( A1 => n59816, A2 => n62115, B1 => n3270, B2 => 
                           n59813, ZN => n10255);
   U11236 : OAI22_X1 port map( A1 => n59816, A2 => n60968, B1 => n3269, B2 => 
                           n59813, ZN => n10256);
   U11237 : OAI22_X1 port map( A1 => n59816, A2 => n60982, B1 => n3268, B2 => 
                           n15268, ZN => n10257);
   U11238 : OAI22_X1 port map( A1 => n59816, A2 => n60996, B1 => n3267, B2 => 
                           n15268, ZN => n10258);
   U11239 : OAI22_X1 port map( A1 => n59816, A2 => n61010, B1 => n3266, B2 => 
                           n15268, ZN => n10259);
   U11240 : OAI22_X1 port map( A1 => n59817, A2 => n61024, B1 => n3265, B2 => 
                           n15268, ZN => n10260);
   U11241 : OAI22_X1 port map( A1 => n59817, A2 => n61038, B1 => n3264, B2 => 
                           n15268, ZN => n10261);
   U11242 : OAI22_X1 port map( A1 => n59817, A2 => n61052, B1 => n3263, B2 => 
                           n15268, ZN => n10262);
   U11243 : OAI22_X1 port map( A1 => n59817, A2 => n61066, B1 => n3262, B2 => 
                           n15268, ZN => n10263);
   U11244 : OAI22_X1 port map( A1 => n59817, A2 => n61080, B1 => n3261, B2 => 
                           n59813, ZN => n10264);
   U11245 : OAI22_X1 port map( A1 => n59818, A2 => n61094, B1 => n3260, B2 => 
                           n59813, ZN => n10265);
   U11246 : OAI22_X1 port map( A1 => n59818, A2 => n61108, B1 => n3259, B2 => 
                           n59813, ZN => n10266);
   U11247 : OAI22_X1 port map( A1 => n59818, A2 => n61122, B1 => n3258, B2 => 
                           n59813, ZN => n10267);
   U11248 : OAI22_X1 port map( A1 => n59818, A2 => n61136, B1 => n3257, B2 => 
                           n59813, ZN => n10268);
   U11249 : OAI22_X1 port map( A1 => n60633, A2 => n61967, B1 => n2022, B2 => 
                           n60632, ZN => n13157);
   U11250 : OAI22_X1 port map( A1 => n60633, A2 => n61981, B1 => n2021, B2 => 
                           n60632, ZN => n13158);
   U11251 : OAI22_X1 port map( A1 => n60633, A2 => n61995, B1 => n2020, B2 => 
                           n60632, ZN => n13159);
   U11252 : OAI22_X1 port map( A1 => n60633, A2 => n62009, B1 => n2019, B2 => 
                           n60632, ZN => n13160);
   U11253 : OAI22_X1 port map( A1 => n60633, A2 => n62023, B1 => n2018, B2 => 
                           n60632, ZN => n13161);
   U11254 : OAI22_X1 port map( A1 => n60634, A2 => n62037, B1 => n2017, B2 => 
                           n60632, ZN => n13162);
   U11255 : OAI22_X1 port map( A1 => n60634, A2 => n62051, B1 => n2016, B2 => 
                           n60632, ZN => n13163);
   U11256 : OAI22_X1 port map( A1 => n60634, A2 => n62065, B1 => n2015, B2 => 
                           n60632, ZN => n13164);
   U11257 : OAI22_X1 port map( A1 => n60634, A2 => n62079, B1 => n2014, B2 => 
                           n60632, ZN => n13165);
   U11258 : OAI22_X1 port map( A1 => n60634, A2 => n62093, B1 => n2013, B2 => 
                           n60632, ZN => n13166);
   U11259 : OAI22_X1 port map( A1 => n60635, A2 => n62107, B1 => n2012, B2 => 
                           n60632, ZN => n13167);
   U11260 : OAI22_X1 port map( A1 => n60635, A2 => n60961, B1 => n2011, B2 => 
                           n60632, ZN => n13168);
   U11261 : OAI22_X1 port map( A1 => n60635, A2 => n60975, B1 => n2010, B2 => 
                           n15151, ZN => n13169);
   U11262 : OAI22_X1 port map( A1 => n60635, A2 => n60989, B1 => n2009, B2 => 
                           n15151, ZN => n13170);
   U11263 : OAI22_X1 port map( A1 => n60635, A2 => n61003, B1 => n2008, B2 => 
                           n15151, ZN => n13171);
   U11264 : OAI22_X1 port map( A1 => n60636, A2 => n61017, B1 => n2007, B2 => 
                           n15151, ZN => n13172);
   U11265 : OAI22_X1 port map( A1 => n60636, A2 => n61031, B1 => n2006, B2 => 
                           n15151, ZN => n13173);
   U11266 : OAI22_X1 port map( A1 => n60636, A2 => n61045, B1 => n2005, B2 => 
                           n15151, ZN => n13174);
   U11267 : OAI22_X1 port map( A1 => n60636, A2 => n61059, B1 => n2004, B2 => 
                           n15151, ZN => n13175);
   U11268 : OAI22_X1 port map( A1 => n60636, A2 => n61073, B1 => n2003, B2 => 
                           n60632, ZN => n13176);
   U11269 : OAI22_X1 port map( A1 => n60637, A2 => n61087, B1 => n2002, B2 => 
                           n60632, ZN => n13177);
   U11270 : OAI22_X1 port map( A1 => n60637, A2 => n61101, B1 => n2001, B2 => 
                           n60632, ZN => n13178);
   U11271 : OAI22_X1 port map( A1 => n60637, A2 => n61115, B1 => n2000, B2 => 
                           n60632, ZN => n13179);
   U11272 : OAI22_X1 port map( A1 => n60637, A2 => n61129, B1 => n1999, B2 => 
                           n60632, ZN => n13180);
   U11273 : OAI22_X1 port map( A1 => n60624, A2 => n61968, B1 => n3644, B2 => 
                           n60623, ZN => n13125);
   U11274 : OAI22_X1 port map( A1 => n60624, A2 => n61982, B1 => n3643, B2 => 
                           n60623, ZN => n13126);
   U11275 : OAI22_X1 port map( A1 => n60624, A2 => n61996, B1 => n3642, B2 => 
                           n60623, ZN => n13127);
   U11276 : OAI22_X1 port map( A1 => n60624, A2 => n62010, B1 => n3641, B2 => 
                           n60623, ZN => n13128);
   U11277 : OAI22_X1 port map( A1 => n60624, A2 => n62024, B1 => n3640, B2 => 
                           n60623, ZN => n13129);
   U11278 : OAI22_X1 port map( A1 => n60625, A2 => n62038, B1 => n3639, B2 => 
                           n60623, ZN => n13130);
   U11279 : OAI22_X1 port map( A1 => n60625, A2 => n62052, B1 => n3638, B2 => 
                           n60623, ZN => n13131);
   U11280 : OAI22_X1 port map( A1 => n60625, A2 => n62066, B1 => n3637, B2 => 
                           n60623, ZN => n13132);
   U11281 : OAI22_X1 port map( A1 => n60625, A2 => n62080, B1 => n3636, B2 => 
                           n60623, ZN => n13133);
   U11282 : OAI22_X1 port map( A1 => n60625, A2 => n62094, B1 => n3635, B2 => 
                           n60623, ZN => n13134);
   U11283 : OAI22_X1 port map( A1 => n60626, A2 => n62108, B1 => n3634, B2 => 
                           n60623, ZN => n13135);
   U11284 : OAI22_X1 port map( A1 => n60626, A2 => n60961, B1 => n3633, B2 => 
                           n60623, ZN => n13136);
   U11285 : OAI22_X1 port map( A1 => n60626, A2 => n60975, B1 => n3632, B2 => 
                           n15152, ZN => n13137);
   U11286 : OAI22_X1 port map( A1 => n60626, A2 => n60989, B1 => n3631, B2 => 
                           n15152, ZN => n13138);
   U11287 : OAI22_X1 port map( A1 => n60626, A2 => n61003, B1 => n3630, B2 => 
                           n15152, ZN => n13139);
   U11288 : OAI22_X1 port map( A1 => n60627, A2 => n61017, B1 => n3629, B2 => 
                           n15152, ZN => n13140);
   U11289 : OAI22_X1 port map( A1 => n60627, A2 => n61031, B1 => n3628, B2 => 
                           n15152, ZN => n13141);
   U11290 : OAI22_X1 port map( A1 => n60627, A2 => n61045, B1 => n3627, B2 => 
                           n15152, ZN => n13142);
   U11291 : OAI22_X1 port map( A1 => n60627, A2 => n61059, B1 => n3626, B2 => 
                           n15152, ZN => n13143);
   U11292 : OAI22_X1 port map( A1 => n60627, A2 => n61073, B1 => n3625, B2 => 
                           n60623, ZN => n13144);
   U11293 : OAI22_X1 port map( A1 => n60628, A2 => n61087, B1 => n3624, B2 => 
                           n60623, ZN => n13145);
   U11294 : OAI22_X1 port map( A1 => n60628, A2 => n61101, B1 => n3623, B2 => 
                           n60623, ZN => n13146);
   U11295 : OAI22_X1 port map( A1 => n60628, A2 => n61115, B1 => n3622, B2 => 
                           n60623, ZN => n13147);
   U11296 : OAI22_X1 port map( A1 => n60628, A2 => n61129, B1 => n3621, B2 => 
                           n60623, ZN => n13148);
   U11297 : OAI22_X1 port map( A1 => n60480, A2 => n61969, B1 => n3126, B2 => 
                           n60479, ZN => n12613);
   U11298 : OAI22_X1 port map( A1 => n60480, A2 => n61983, B1 => n3125, B2 => 
                           n60479, ZN => n12614);
   U11299 : OAI22_X1 port map( A1 => n60480, A2 => n61997, B1 => n3124, B2 => 
                           n60479, ZN => n12615);
   U11300 : OAI22_X1 port map( A1 => n60480, A2 => n62011, B1 => n3123, B2 => 
                           n60479, ZN => n12616);
   U11301 : OAI22_X1 port map( A1 => n60480, A2 => n62025, B1 => n3098, B2 => 
                           n60479, ZN => n12617);
   U11302 : OAI22_X1 port map( A1 => n60481, A2 => n62039, B1 => n3097, B2 => 
                           n60479, ZN => n12618);
   U11303 : OAI22_X1 port map( A1 => n60481, A2 => n62053, B1 => n3096, B2 => 
                           n60479, ZN => n12619);
   U11304 : OAI22_X1 port map( A1 => n60481, A2 => n62067, B1 => n3095, B2 => 
                           n60479, ZN => n12620);
   U11305 : OAI22_X1 port map( A1 => n60481, A2 => n62081, B1 => n3094, B2 => 
                           n60479, ZN => n12621);
   U11306 : OAI22_X1 port map( A1 => n60481, A2 => n62095, B1 => n3093, B2 => 
                           n60479, ZN => n12622);
   U11307 : OAI22_X1 port map( A1 => n60482, A2 => n62109, B1 => n3092, B2 => 
                           n60479, ZN => n12623);
   U11308 : OAI22_X1 port map( A1 => n60482, A2 => n60962, B1 => n3091, B2 => 
                           n60479, ZN => n12624);
   U11309 : OAI22_X1 port map( A1 => n60482, A2 => n60976, B1 => n3090, B2 => 
                           n15169, ZN => n12625);
   U11310 : OAI22_X1 port map( A1 => n60482, A2 => n60990, B1 => n3089, B2 => 
                           n15169, ZN => n12626);
   U11311 : OAI22_X1 port map( A1 => n60482, A2 => n61004, B1 => n3088, B2 => 
                           n15169, ZN => n12627);
   U11312 : OAI22_X1 port map( A1 => n60483, A2 => n61018, B1 => n3087, B2 => 
                           n15169, ZN => n12628);
   U11313 : OAI22_X1 port map( A1 => n60483, A2 => n61032, B1 => n3086, B2 => 
                           n15169, ZN => n12629);
   U11314 : OAI22_X1 port map( A1 => n60483, A2 => n61046, B1 => n3085, B2 => 
                           n15169, ZN => n12630);
   U11315 : OAI22_X1 port map( A1 => n60483, A2 => n61060, B1 => n3084, B2 => 
                           n15169, ZN => n12631);
   U11316 : OAI22_X1 port map( A1 => n60483, A2 => n61074, B1 => n3083, B2 => 
                           n60479, ZN => n12632);
   U11317 : OAI22_X1 port map( A1 => n60484, A2 => n61088, B1 => n3082, B2 => 
                           n60479, ZN => n12633);
   U11318 : OAI22_X1 port map( A1 => n60484, A2 => n61102, B1 => n3081, B2 => 
                           n60479, ZN => n12634);
   U11319 : OAI22_X1 port map( A1 => n60484, A2 => n61116, B1 => n3080, B2 => 
                           n60479, ZN => n12635);
   U11320 : OAI22_X1 port map( A1 => n60484, A2 => n61130, B1 => n3079, B2 => 
                           n60479, ZN => n12636);
   U11321 : OAI22_X1 port map( A1 => n60471, A2 => n61969, B1 => n3078, B2 => 
                           n60470, ZN => n12581);
   U11322 : OAI22_X1 port map( A1 => n60471, A2 => n61983, B1 => n3077, B2 => 
                           n60470, ZN => n12582);
   U11323 : OAI22_X1 port map( A1 => n60471, A2 => n61997, B1 => n3076, B2 => 
                           n60470, ZN => n12583);
   U11324 : OAI22_X1 port map( A1 => n60471, A2 => n62011, B1 => n3075, B2 => 
                           n60470, ZN => n12584);
   U11325 : OAI22_X1 port map( A1 => n60471, A2 => n62025, B1 => n3074, B2 => 
                           n60470, ZN => n12585);
   U11326 : OAI22_X1 port map( A1 => n60472, A2 => n62039, B1 => n3073, B2 => 
                           n60470, ZN => n12586);
   U11327 : OAI22_X1 port map( A1 => n60472, A2 => n62053, B1 => n3072, B2 => 
                           n60470, ZN => n12587);
   U11328 : OAI22_X1 port map( A1 => n60472, A2 => n62067, B1 => n3071, B2 => 
                           n60470, ZN => n12588);
   U11329 : OAI22_X1 port map( A1 => n60472, A2 => n62081, B1 => n3070, B2 => 
                           n60470, ZN => n12589);
   U11330 : OAI22_X1 port map( A1 => n60472, A2 => n62095, B1 => n3069, B2 => 
                           n60470, ZN => n12590);
   U11331 : OAI22_X1 port map( A1 => n60473, A2 => n62109, B1 => n3068, B2 => 
                           n60470, ZN => n12591);
   U11332 : OAI22_X1 port map( A1 => n60473, A2 => n60962, B1 => n3067, B2 => 
                           n60470, ZN => n12592);
   U11333 : OAI22_X1 port map( A1 => n60473, A2 => n60976, B1 => n3066, B2 => 
                           n15170, ZN => n12593);
   U11334 : OAI22_X1 port map( A1 => n60473, A2 => n60990, B1 => n3065, B2 => 
                           n15170, ZN => n12594);
   U11335 : OAI22_X1 port map( A1 => n60473, A2 => n61004, B1 => n3064, B2 => 
                           n15170, ZN => n12595);
   U11336 : OAI22_X1 port map( A1 => n60474, A2 => n61018, B1 => n3063, B2 => 
                           n15170, ZN => n12596);
   U11337 : OAI22_X1 port map( A1 => n60474, A2 => n61032, B1 => n3062, B2 => 
                           n15170, ZN => n12597);
   U11338 : OAI22_X1 port map( A1 => n60474, A2 => n61046, B1 => n3061, B2 => 
                           n15170, ZN => n12598);
   U11339 : OAI22_X1 port map( A1 => n60474, A2 => n61060, B1 => n3060, B2 => 
                           n15170, ZN => n12599);
   U11340 : OAI22_X1 port map( A1 => n60474, A2 => n61074, B1 => n3059, B2 => 
                           n60470, ZN => n12600);
   U11341 : OAI22_X1 port map( A1 => n60475, A2 => n61088, B1 => n3058, B2 => 
                           n60470, ZN => n12601);
   U11342 : OAI22_X1 port map( A1 => n60475, A2 => n61102, B1 => n3057, B2 => 
                           n60470, ZN => n12602);
   U11343 : OAI22_X1 port map( A1 => n60475, A2 => n61116, B1 => n3056, B2 => 
                           n60470, ZN => n12603);
   U11344 : OAI22_X1 port map( A1 => n60475, A2 => n61130, B1 => n3055, B2 => 
                           n60470, ZN => n12604);
   U11345 : OAI22_X1 port map( A1 => n60453, A2 => n61969, B1 => n3030, B2 => 
                           n60452, ZN => n12517);
   U11346 : OAI22_X1 port map( A1 => n60453, A2 => n61983, B1 => n3029, B2 => 
                           n60452, ZN => n12518);
   U11347 : OAI22_X1 port map( A1 => n60453, A2 => n61997, B1 => n3028, B2 => 
                           n60452, ZN => n12519);
   U11348 : OAI22_X1 port map( A1 => n60453, A2 => n62011, B1 => n3027, B2 => 
                           n60452, ZN => n12520);
   U11349 : OAI22_X1 port map( A1 => n60453, A2 => n62025, B1 => n2978, B2 => 
                           n60452, ZN => n12521);
   U11350 : OAI22_X1 port map( A1 => n60454, A2 => n62039, B1 => n2977, B2 => 
                           n60452, ZN => n12522);
   U11351 : OAI22_X1 port map( A1 => n60454, A2 => n62053, B1 => n2976, B2 => 
                           n60452, ZN => n12523);
   U11352 : OAI22_X1 port map( A1 => n60454, A2 => n62067, B1 => n2975, B2 => 
                           n60452, ZN => n12524);
   U11353 : OAI22_X1 port map( A1 => n60454, A2 => n62081, B1 => n2974, B2 => 
                           n60452, ZN => n12525);
   U11354 : OAI22_X1 port map( A1 => n60454, A2 => n62095, B1 => n2973, B2 => 
                           n60452, ZN => n12526);
   U11355 : OAI22_X1 port map( A1 => n60455, A2 => n62109, B1 => n2972, B2 => 
                           n60452, ZN => n12527);
   U11356 : OAI22_X1 port map( A1 => n60455, A2 => n60962, B1 => n2971, B2 => 
                           n60452, ZN => n12528);
   U11357 : OAI22_X1 port map( A1 => n60455, A2 => n60976, B1 => n2970, B2 => 
                           n15179, ZN => n12529);
   U11358 : OAI22_X1 port map( A1 => n60455, A2 => n60990, B1 => n2969, B2 => 
                           n15179, ZN => n12530);
   U11359 : OAI22_X1 port map( A1 => n60455, A2 => n61004, B1 => n2968, B2 => 
                           n15179, ZN => n12531);
   U11360 : OAI22_X1 port map( A1 => n60456, A2 => n61018, B1 => n2967, B2 => 
                           n15179, ZN => n12532);
   U11361 : OAI22_X1 port map( A1 => n60456, A2 => n61032, B1 => n2966, B2 => 
                           n15179, ZN => n12533);
   U11362 : OAI22_X1 port map( A1 => n60456, A2 => n61046, B1 => n2965, B2 => 
                           n15179, ZN => n12534);
   U11363 : OAI22_X1 port map( A1 => n60456, A2 => n61060, B1 => n2964, B2 => 
                           n15179, ZN => n12535);
   U11364 : OAI22_X1 port map( A1 => n60456, A2 => n61074, B1 => n2963, B2 => 
                           n60452, ZN => n12536);
   U11365 : OAI22_X1 port map( A1 => n60457, A2 => n61088, B1 => n2962, B2 => 
                           n60452, ZN => n12537);
   U11366 : OAI22_X1 port map( A1 => n60457, A2 => n61102, B1 => n2961, B2 => 
                           n60452, ZN => n12538);
   U11367 : OAI22_X1 port map( A1 => n60457, A2 => n61116, B1 => n2960, B2 => 
                           n60452, ZN => n12539);
   U11368 : OAI22_X1 port map( A1 => n60457, A2 => n61130, B1 => n2959, B2 => 
                           n60452, ZN => n12540);
   U11369 : OAI22_X1 port map( A1 => n60390, A2 => n61970, B1 => n1692, B2 => 
                           n60389, ZN => n12293);
   U11370 : OAI22_X1 port map( A1 => n60390, A2 => n61984, B1 => n1691, B2 => 
                           n60389, ZN => n12294);
   U11371 : OAI22_X1 port map( A1 => n60390, A2 => n61998, B1 => n1690, B2 => 
                           n60389, ZN => n12295);
   U11372 : OAI22_X1 port map( A1 => n60390, A2 => n62012, B1 => n1689, B2 => 
                           n60389, ZN => n12296);
   U11373 : OAI22_X1 port map( A1 => n60390, A2 => n62026, B1 => n1688, B2 => 
                           n60389, ZN => n12297);
   U11374 : OAI22_X1 port map( A1 => n60391, A2 => n62040, B1 => n1687, B2 => 
                           n60389, ZN => n12298);
   U11375 : OAI22_X1 port map( A1 => n60391, A2 => n62054, B1 => n1686, B2 => 
                           n60389, ZN => n12299);
   U11376 : OAI22_X1 port map( A1 => n60391, A2 => n62068, B1 => n1685, B2 => 
                           n60389, ZN => n12300);
   U11377 : OAI22_X1 port map( A1 => n60391, A2 => n62082, B1 => n1684, B2 => 
                           n60389, ZN => n12301);
   U11378 : OAI22_X1 port map( A1 => n60391, A2 => n62096, B1 => n1683, B2 => 
                           n60389, ZN => n12302);
   U11379 : OAI22_X1 port map( A1 => n60392, A2 => n62110, B1 => n1682, B2 => 
                           n60389, ZN => n12303);
   U11380 : OAI22_X1 port map( A1 => n60392, A2 => n60963, B1 => n1681, B2 => 
                           n60389, ZN => n12304);
   U11381 : OAI22_X1 port map( A1 => n60392, A2 => n60977, B1 => n1680, B2 => 
                           n15186, ZN => n12305);
   U11382 : OAI22_X1 port map( A1 => n60392, A2 => n60991, B1 => n1679, B2 => 
                           n15186, ZN => n12306);
   U11383 : OAI22_X1 port map( A1 => n60392, A2 => n61005, B1 => n1678, B2 => 
                           n15186, ZN => n12307);
   U11384 : OAI22_X1 port map( A1 => n60393, A2 => n61019, B1 => n1677, B2 => 
                           n15186, ZN => n12308);
   U11385 : OAI22_X1 port map( A1 => n60393, A2 => n61033, B1 => n1676, B2 => 
                           n15186, ZN => n12309);
   U11386 : OAI22_X1 port map( A1 => n60393, A2 => n61047, B1 => n1675, B2 => 
                           n15186, ZN => n12310);
   U11387 : OAI22_X1 port map( A1 => n60393, A2 => n61061, B1 => n1674, B2 => 
                           n15186, ZN => n12311);
   U11388 : OAI22_X1 port map( A1 => n60393, A2 => n61075, B1 => n1673, B2 => 
                           n60389, ZN => n12312);
   U11389 : OAI22_X1 port map( A1 => n60394, A2 => n61089, B1 => n1672, B2 => 
                           n60389, ZN => n12313);
   U11390 : OAI22_X1 port map( A1 => n60394, A2 => n61103, B1 => n1671, B2 => 
                           n60389, ZN => n12314);
   U11391 : OAI22_X1 port map( A1 => n60394, A2 => n61117, B1 => n1670, B2 => 
                           n60389, ZN => n12315);
   U11392 : OAI22_X1 port map( A1 => n60394, A2 => n61131, B1 => n1669, B2 => 
                           n60389, ZN => n12316);
   U11393 : OAI22_X1 port map( A1 => n61237, A2 => n61965, B1 => n2078, B2 => 
                           n61236, ZN => n14309);
   U11394 : OAI22_X1 port map( A1 => n61237, A2 => n61979, B1 => n2270, B2 => 
                           n61236, ZN => n14310);
   U11395 : OAI22_X1 port map( A1 => n61237, A2 => n61993, B1 => n2269, B2 => 
                           n61236, ZN => n14311);
   U11396 : OAI22_X1 port map( A1 => n61237, A2 => n62007, B1 => n2268, B2 => 
                           n61236, ZN => n14312);
   U11397 : OAI22_X1 port map( A1 => n61237, A2 => n62021, B1 => n2267, B2 => 
                           n61236, ZN => n14313);
   U11398 : OAI22_X1 port map( A1 => n61238, A2 => n62035, B1 => n2266, B2 => 
                           n61236, ZN => n14314);
   U11399 : OAI22_X1 port map( A1 => n61238, A2 => n62049, B1 => n2265, B2 => 
                           n61236, ZN => n14315);
   U11400 : OAI22_X1 port map( A1 => n61238, A2 => n62063, B1 => n2264, B2 => 
                           n61236, ZN => n14316);
   U11401 : OAI22_X1 port map( A1 => n61238, A2 => n62077, B1 => n2263, B2 => 
                           n61236, ZN => n14317);
   U11402 : OAI22_X1 port map( A1 => n61238, A2 => n62091, B1 => n2262, B2 => 
                           n61236, ZN => n14318);
   U11403 : OAI22_X1 port map( A1 => n61239, A2 => n62105, B1 => n2261, B2 => 
                           n61236, ZN => n14319);
   U11404 : OAI22_X1 port map( A1 => n61239, A2 => n60958, B1 => n2077, B2 => 
                           n61236, ZN => n14320);
   U11405 : OAI22_X1 port map( A1 => n61239, A2 => n60972, B1 => n2260, B2 => 
                           n15073, ZN => n14321);
   U11406 : OAI22_X1 port map( A1 => n61239, A2 => n60986, B1 => n2259, B2 => 
                           n15073, ZN => n14322);
   U11407 : OAI22_X1 port map( A1 => n61239, A2 => n61000, B1 => n2258, B2 => 
                           n15073, ZN => n14323);
   U11408 : OAI22_X1 port map( A1 => n61240, A2 => n61014, B1 => n2257, B2 => 
                           n15073, ZN => n14324);
   U11409 : OAI22_X1 port map( A1 => n61240, A2 => n61028, B1 => n2256, B2 => 
                           n15073, ZN => n14325);
   U11410 : OAI22_X1 port map( A1 => n61240, A2 => n61042, B1 => n2255, B2 => 
                           n15073, ZN => n14326);
   U11411 : OAI22_X1 port map( A1 => n61240, A2 => n61056, B1 => n2254, B2 => 
                           n15073, ZN => n14327);
   U11412 : OAI22_X1 port map( A1 => n61240, A2 => n61070, B1 => n2253, B2 => 
                           n61236, ZN => n14328);
   U11413 : OAI22_X1 port map( A1 => n61241, A2 => n61084, B1 => n2252, B2 => 
                           n61236, ZN => n14329);
   U11414 : OAI22_X1 port map( A1 => n61241, A2 => n61098, B1 => n2251, B2 => 
                           n61236, ZN => n14330);
   U11415 : OAI22_X1 port map( A1 => n61241, A2 => n61112, B1 => n2250, B2 => 
                           n61236, ZN => n14331);
   U11416 : OAI22_X1 port map( A1 => n61241, A2 => n61126, B1 => n2249, B2 => 
                           n61236, ZN => n14332);
   U11417 : OAI22_X1 port map( A1 => n60867, A2 => n61965, B1 => n2748, B2 => 
                           n60866, ZN => n13989);
   U11418 : OAI22_X1 port map( A1 => n60867, A2 => n61979, B1 => n2747, B2 => 
                           n60866, ZN => n13990);
   U11419 : OAI22_X1 port map( A1 => n60867, A2 => n61993, B1 => n2746, B2 => 
                           n60866, ZN => n13991);
   U11420 : OAI22_X1 port map( A1 => n60867, A2 => n62007, B1 => n2745, B2 => 
                           n60866, ZN => n13992);
   U11421 : OAI22_X1 port map( A1 => n60867, A2 => n62021, B1 => n2744, B2 => 
                           n60866, ZN => n13993);
   U11422 : OAI22_X1 port map( A1 => n60868, A2 => n62035, B1 => n2743, B2 => 
                           n60866, ZN => n13994);
   U11423 : OAI22_X1 port map( A1 => n60868, A2 => n62049, B1 => n2742, B2 => 
                           n60866, ZN => n13995);
   U11424 : OAI22_X1 port map( A1 => n60868, A2 => n62063, B1 => n2741, B2 => 
                           n60866, ZN => n13996);
   U11425 : OAI22_X1 port map( A1 => n60868, A2 => n62077, B1 => n2740, B2 => 
                           n60866, ZN => n13997);
   U11426 : OAI22_X1 port map( A1 => n60868, A2 => n62091, B1 => n2739, B2 => 
                           n60866, ZN => n13998);
   U11427 : OAI22_X1 port map( A1 => n60869, A2 => n62105, B1 => n2738, B2 => 
                           n60866, ZN => n13999);
   U11428 : OAI22_X1 port map( A1 => n60869, A2 => n60958, B1 => n2737, B2 => 
                           n60866, ZN => n14000);
   U11429 : OAI22_X1 port map( A1 => n60869, A2 => n60972, B1 => n2736, B2 => 
                           n15114, ZN => n14001);
   U11430 : OAI22_X1 port map( A1 => n60869, A2 => n60986, B1 => n2735, B2 => 
                           n15114, ZN => n14002);
   U11431 : OAI22_X1 port map( A1 => n60869, A2 => n61000, B1 => n2734, B2 => 
                           n15114, ZN => n14003);
   U11432 : OAI22_X1 port map( A1 => n60870, A2 => n61014, B1 => n2733, B2 => 
                           n15114, ZN => n14004);
   U11433 : OAI22_X1 port map( A1 => n60870, A2 => n61028, B1 => n2732, B2 => 
                           n15114, ZN => n14005);
   U11434 : OAI22_X1 port map( A1 => n60870, A2 => n61042, B1 => n2731, B2 => 
                           n15114, ZN => n14006);
   U11435 : OAI22_X1 port map( A1 => n60870, A2 => n61056, B1 => n2730, B2 => 
                           n15114, ZN => n14007);
   U11436 : OAI22_X1 port map( A1 => n60870, A2 => n61070, B1 => n2729, B2 => 
                           n60866, ZN => n14008);
   U11437 : OAI22_X1 port map( A1 => n60871, A2 => n61084, B1 => n2728, B2 => 
                           n60866, ZN => n14009);
   U11438 : OAI22_X1 port map( A1 => n60871, A2 => n61098, B1 => n2727, B2 => 
                           n60866, ZN => n14010);
   U11439 : OAI22_X1 port map( A1 => n60871, A2 => n61112, B1 => n2726, B2 => 
                           n60866, ZN => n14011);
   U11440 : OAI22_X1 port map( A1 => n60871, A2 => n61126, B1 => n2725, B2 => 
                           n60866, ZN => n14012);
   U11441 : OAI22_X1 port map( A1 => n60381, A2 => n61970, B1 => n452, B2 => 
                           n60380, ZN => n12261);
   U11442 : OAI22_X1 port map( A1 => n60381, A2 => n61984, B1 => n435, B2 => 
                           n60380, ZN => n12262);
   U11443 : OAI22_X1 port map( A1 => n60381, A2 => n61998, B1 => n434, B2 => 
                           n60380, ZN => n12263);
   U11444 : OAI22_X1 port map( A1 => n60381, A2 => n62012, B1 => n433, B2 => 
                           n60380, ZN => n12264);
   U11445 : OAI22_X1 port map( A1 => n60381, A2 => n62026, B1 => n432, B2 => 
                           n60380, ZN => n12265);
   U11446 : OAI22_X1 port map( A1 => n60382, A2 => n62040, B1 => n431, B2 => 
                           n60380, ZN => n12266);
   U11447 : OAI22_X1 port map( A1 => n60382, A2 => n62054, B1 => n430, B2 => 
                           n60380, ZN => n12267);
   U11448 : OAI22_X1 port map( A1 => n60382, A2 => n62068, B1 => n429, B2 => 
                           n60380, ZN => n12268);
   U11449 : OAI22_X1 port map( A1 => n60382, A2 => n62082, B1 => n428, B2 => 
                           n60380, ZN => n12269);
   U11450 : OAI22_X1 port map( A1 => n60382, A2 => n62096, B1 => n427, B2 => 
                           n60380, ZN => n12270);
   U11451 : OAI22_X1 port map( A1 => n60383, A2 => n62110, B1 => n426, B2 => 
                           n60380, ZN => n12271);
   U11452 : OAI22_X1 port map( A1 => n60383, A2 => n60963, B1 => n425, B2 => 
                           n60380, ZN => n12272);
   U11453 : OAI22_X1 port map( A1 => n60383, A2 => n60977, B1 => n424, B2 => 
                           n15187, ZN => n12273);
   U11454 : OAI22_X1 port map( A1 => n60383, A2 => n60991, B1 => n423, B2 => 
                           n15187, ZN => n12274);
   U11455 : OAI22_X1 port map( A1 => n60383, A2 => n61005, B1 => n422, B2 => 
                           n15187, ZN => n12275);
   U11456 : OAI22_X1 port map( A1 => n60384, A2 => n61019, B1 => n421, B2 => 
                           n15187, ZN => n12276);
   U11457 : OAI22_X1 port map( A1 => n60384, A2 => n61033, B1 => n420, B2 => 
                           n15187, ZN => n12277);
   U11458 : OAI22_X1 port map( A1 => n60384, A2 => n61047, B1 => n419, B2 => 
                           n15187, ZN => n12278);
   U11459 : OAI22_X1 port map( A1 => n60384, A2 => n61061, B1 => n418, B2 => 
                           n15187, ZN => n12279);
   U11460 : OAI22_X1 port map( A1 => n60384, A2 => n61075, B1 => n417, B2 => 
                           n60380, ZN => n12280);
   U11461 : OAI22_X1 port map( A1 => n60385, A2 => n61089, B1 => n416, B2 => 
                           n60380, ZN => n12281);
   U11462 : OAI22_X1 port map( A1 => n60385, A2 => n61103, B1 => n415, B2 => 
                           n60380, ZN => n12282);
   U11463 : OAI22_X1 port map( A1 => n60385, A2 => n61117, B1 => n414, B2 => 
                           n60380, ZN => n12283);
   U11464 : OAI22_X1 port map( A1 => n60385, A2 => n61131, B1 => n413, B2 => 
                           n60380, ZN => n12284);
   U11465 : OAI22_X1 port map( A1 => n60354, A2 => n61970, B1 => n2676, B2 => 
                           n60353, ZN => n12165);
   U11466 : OAI22_X1 port map( A1 => n60354, A2 => n61984, B1 => n2675, B2 => 
                           n60353, ZN => n12166);
   U11467 : OAI22_X1 port map( A1 => n60354, A2 => n61998, B1 => n2674, B2 => 
                           n60353, ZN => n12167);
   U11468 : OAI22_X1 port map( A1 => n60354, A2 => n62012, B1 => n2673, B2 => 
                           n60353, ZN => n12168);
   U11469 : OAI22_X1 port map( A1 => n60354, A2 => n62026, B1 => n2672, B2 => 
                           n60353, ZN => n12169);
   U11470 : OAI22_X1 port map( A1 => n60355, A2 => n62040, B1 => n2671, B2 => 
                           n60353, ZN => n12170);
   U11471 : OAI22_X1 port map( A1 => n60355, A2 => n62054, B1 => n2670, B2 => 
                           n60353, ZN => n12171);
   U11472 : OAI22_X1 port map( A1 => n60355, A2 => n62068, B1 => n2669, B2 => 
                           n60353, ZN => n12172);
   U11473 : OAI22_X1 port map( A1 => n60355, A2 => n62082, B1 => n2668, B2 => 
                           n60353, ZN => n12173);
   U11474 : OAI22_X1 port map( A1 => n60355, A2 => n62096, B1 => n2667, B2 => 
                           n60353, ZN => n12174);
   U11475 : OAI22_X1 port map( A1 => n60356, A2 => n62110, B1 => n2666, B2 => 
                           n60353, ZN => n12175);
   U11476 : OAI22_X1 port map( A1 => n60356, A2 => n60963, B1 => n2665, B2 => 
                           n60353, ZN => n12176);
   U11477 : OAI22_X1 port map( A1 => n60356, A2 => n60977, B1 => n2664, B2 => 
                           n15191, ZN => n12177);
   U11478 : OAI22_X1 port map( A1 => n60356, A2 => n60991, B1 => n2663, B2 => 
                           n15191, ZN => n12178);
   U11479 : OAI22_X1 port map( A1 => n60356, A2 => n61005, B1 => n2662, B2 => 
                           n15191, ZN => n12179);
   U11480 : OAI22_X1 port map( A1 => n60357, A2 => n61019, B1 => n2661, B2 => 
                           n15191, ZN => n12180);
   U11481 : OAI22_X1 port map( A1 => n60357, A2 => n61033, B1 => n2660, B2 => 
                           n15191, ZN => n12181);
   U11482 : OAI22_X1 port map( A1 => n60357, A2 => n61047, B1 => n2659, B2 => 
                           n15191, ZN => n12182);
   U11483 : OAI22_X1 port map( A1 => n60357, A2 => n61061, B1 => n2658, B2 => 
                           n15191, ZN => n12183);
   U11484 : OAI22_X1 port map( A1 => n60357, A2 => n61075, B1 => n2657, B2 => 
                           n60353, ZN => n12184);
   U11485 : OAI22_X1 port map( A1 => n60358, A2 => n61089, B1 => n2656, B2 => 
                           n60353, ZN => n12185);
   U11486 : OAI22_X1 port map( A1 => n60358, A2 => n61103, B1 => n2655, B2 => 
                           n60353, ZN => n12186);
   U11487 : OAI22_X1 port map( A1 => n60358, A2 => n61117, B1 => n2654, B2 => 
                           n60353, ZN => n12187);
   U11488 : OAI22_X1 port map( A1 => n60358, A2 => n61131, B1 => n2653, B2 => 
                           n60353, ZN => n12188);
   U11489 : OAI22_X1 port map( A1 => n60327, A2 => n61970, B1 => n2597, B2 => 
                           n60326, ZN => n12069);
   U11490 : OAI22_X1 port map( A1 => n60327, A2 => n61984, B1 => n2596, B2 => 
                           n60326, ZN => n12070);
   U11491 : OAI22_X1 port map( A1 => n60327, A2 => n61998, B1 => n2595, B2 => 
                           n60326, ZN => n12071);
   U11492 : OAI22_X1 port map( A1 => n60327, A2 => n62012, B1 => n2594, B2 => 
                           n60326, ZN => n12072);
   U11493 : OAI22_X1 port map( A1 => n60327, A2 => n62026, B1 => n2593, B2 => 
                           n60326, ZN => n12073);
   U11494 : OAI22_X1 port map( A1 => n60328, A2 => n62040, B1 => n2592, B2 => 
                           n60326, ZN => n12074);
   U11495 : OAI22_X1 port map( A1 => n60328, A2 => n62054, B1 => n2591, B2 => 
                           n60326, ZN => n12075);
   U11496 : OAI22_X1 port map( A1 => n60328, A2 => n62068, B1 => n2590, B2 => 
                           n60326, ZN => n12076);
   U11497 : OAI22_X1 port map( A1 => n60328, A2 => n62082, B1 => n2589, B2 => 
                           n60326, ZN => n12077);
   U11498 : OAI22_X1 port map( A1 => n60328, A2 => n62096, B1 => n2588, B2 => 
                           n60326, ZN => n12078);
   U11499 : OAI22_X1 port map( A1 => n60329, A2 => n62110, B1 => n2587, B2 => 
                           n60326, ZN => n12079);
   U11500 : OAI22_X1 port map( A1 => n60329, A2 => n60963, B1 => n2586, B2 => 
                           n60326, ZN => n12080);
   U11501 : OAI22_X1 port map( A1 => n60329, A2 => n60977, B1 => n2585, B2 => 
                           n15194, ZN => n12081);
   U11502 : OAI22_X1 port map( A1 => n60329, A2 => n60991, B1 => n2584, B2 => 
                           n15194, ZN => n12082);
   U11503 : OAI22_X1 port map( A1 => n60329, A2 => n61005, B1 => n2583, B2 => 
                           n15194, ZN => n12083);
   U11504 : OAI22_X1 port map( A1 => n60330, A2 => n61019, B1 => n2582, B2 => 
                           n15194, ZN => n12084);
   U11505 : OAI22_X1 port map( A1 => n60330, A2 => n61033, B1 => n2581, B2 => 
                           n15194, ZN => n12085);
   U11506 : OAI22_X1 port map( A1 => n60330, A2 => n61047, B1 => n2580, B2 => 
                           n15194, ZN => n12086);
   U11507 : OAI22_X1 port map( A1 => n60330, A2 => n61061, B1 => n2579, B2 => 
                           n15194, ZN => n12087);
   U11508 : OAI22_X1 port map( A1 => n60330, A2 => n61075, B1 => n2578, B2 => 
                           n60326, ZN => n12088);
   U11509 : OAI22_X1 port map( A1 => n60331, A2 => n61089, B1 => n2577, B2 => 
                           n60326, ZN => n12089);
   U11510 : OAI22_X1 port map( A1 => n60331, A2 => n61103, B1 => n2576, B2 => 
                           n60326, ZN => n12090);
   U11511 : OAI22_X1 port map( A1 => n60331, A2 => n61117, B1 => n2575, B2 => 
                           n60326, ZN => n12091);
   U11512 : OAI22_X1 port map( A1 => n60331, A2 => n61131, B1 => n2574, B2 => 
                           n60326, ZN => n12092);
   U11513 : OAI22_X1 port map( A1 => n60318, A2 => n61970, B1 => n2573, B2 => 
                           n60317, ZN => n12037);
   U11514 : OAI22_X1 port map( A1 => n60318, A2 => n61984, B1 => n2572, B2 => 
                           n60317, ZN => n12038);
   U11515 : OAI22_X1 port map( A1 => n60318, A2 => n61998, B1 => n2571, B2 => 
                           n60317, ZN => n12039);
   U11516 : OAI22_X1 port map( A1 => n60318, A2 => n62012, B1 => n2570, B2 => 
                           n60317, ZN => n12040);
   U11517 : OAI22_X1 port map( A1 => n60318, A2 => n62026, B1 => n2569, B2 => 
                           n60317, ZN => n12041);
   U11518 : OAI22_X1 port map( A1 => n60319, A2 => n62040, B1 => n2568, B2 => 
                           n60317, ZN => n12042);
   U11519 : OAI22_X1 port map( A1 => n60319, A2 => n62054, B1 => n2567, B2 => 
                           n60317, ZN => n12043);
   U11520 : OAI22_X1 port map( A1 => n60319, A2 => n62068, B1 => n2566, B2 => 
                           n60317, ZN => n12044);
   U11521 : OAI22_X1 port map( A1 => n60319, A2 => n62082, B1 => n2565, B2 => 
                           n60317, ZN => n12045);
   U11522 : OAI22_X1 port map( A1 => n60319, A2 => n62096, B1 => n2564, B2 => 
                           n60317, ZN => n12046);
   U11523 : OAI22_X1 port map( A1 => n60320, A2 => n62110, B1 => n2563, B2 => 
                           n60317, ZN => n12047);
   U11524 : OAI22_X1 port map( A1 => n60320, A2 => n60963, B1 => n2562, B2 => 
                           n60317, ZN => n12048);
   U11525 : OAI22_X1 port map( A1 => n60320, A2 => n60977, B1 => n2561, B2 => 
                           n15195, ZN => n12049);
   U11526 : OAI22_X1 port map( A1 => n60320, A2 => n60991, B1 => n2560, B2 => 
                           n15195, ZN => n12050);
   U11527 : OAI22_X1 port map( A1 => n60320, A2 => n61005, B1 => n2559, B2 => 
                           n15195, ZN => n12051);
   U11528 : OAI22_X1 port map( A1 => n60321, A2 => n61019, B1 => n2558, B2 => 
                           n15195, ZN => n12052);
   U11529 : OAI22_X1 port map( A1 => n60321, A2 => n61033, B1 => n2557, B2 => 
                           n15195, ZN => n12053);
   U11530 : OAI22_X1 port map( A1 => n60321, A2 => n61047, B1 => n2556, B2 => 
                           n15195, ZN => n12054);
   U11531 : OAI22_X1 port map( A1 => n60321, A2 => n61061, B1 => n2555, B2 => 
                           n15195, ZN => n12055);
   U11532 : OAI22_X1 port map( A1 => n60321, A2 => n61075, B1 => n2554, B2 => 
                           n60317, ZN => n12056);
   U11533 : OAI22_X1 port map( A1 => n60322, A2 => n61089, B1 => n2553, B2 => 
                           n60317, ZN => n12057);
   U11534 : OAI22_X1 port map( A1 => n60322, A2 => n61103, B1 => n2552, B2 => 
                           n60317, ZN => n12058);
   U11535 : OAI22_X1 port map( A1 => n60322, A2 => n61117, B1 => n2551, B2 => 
                           n60317, ZN => n12059);
   U11536 : OAI22_X1 port map( A1 => n60322, A2 => n61131, B1 => n2550, B2 => 
                           n60317, ZN => n12060);
   U11537 : OAI22_X1 port map( A1 => n60291, A2 => n61971, B1 => n2473, B2 => 
                           n60290, ZN => n11941);
   U11538 : OAI22_X1 port map( A1 => n60291, A2 => n61985, B1 => n2472, B2 => 
                           n60290, ZN => n11942);
   U11539 : OAI22_X1 port map( A1 => n60291, A2 => n61999, B1 => n2471, B2 => 
                           n60290, ZN => n11943);
   U11540 : OAI22_X1 port map( A1 => n60291, A2 => n62013, B1 => n2470, B2 => 
                           n60290, ZN => n11944);
   U11541 : OAI22_X1 port map( A1 => n60291, A2 => n62027, B1 => n2469, B2 => 
                           n60290, ZN => n11945);
   U11542 : OAI22_X1 port map( A1 => n60292, A2 => n62041, B1 => n2468, B2 => 
                           n60290, ZN => n11946);
   U11543 : OAI22_X1 port map( A1 => n60292, A2 => n62055, B1 => n2467, B2 => 
                           n60290, ZN => n11947);
   U11544 : OAI22_X1 port map( A1 => n60292, A2 => n62069, B1 => n2466, B2 => 
                           n60290, ZN => n11948);
   U11545 : OAI22_X1 port map( A1 => n60292, A2 => n62083, B1 => n2465, B2 => 
                           n60290, ZN => n11949);
   U11546 : OAI22_X1 port map( A1 => n60292, A2 => n62097, B1 => n2464, B2 => 
                           n60290, ZN => n11950);
   U11547 : OAI22_X1 port map( A1 => n60293, A2 => n62111, B1 => n2463, B2 => 
                           n60290, ZN => n11951);
   U11548 : OAI22_X1 port map( A1 => n60293, A2 => n60964, B1 => n2438, B2 => 
                           n60290, ZN => n11952);
   U11549 : OAI22_X1 port map( A1 => n60293, A2 => n60978, B1 => n2437, B2 => 
                           n15198, ZN => n11953);
   U11550 : OAI22_X1 port map( A1 => n60293, A2 => n60992, B1 => n2436, B2 => 
                           n15198, ZN => n11954);
   U11551 : OAI22_X1 port map( A1 => n60293, A2 => n61006, B1 => n2435, B2 => 
                           n15198, ZN => n11955);
   U11552 : OAI22_X1 port map( A1 => n60294, A2 => n61020, B1 => n2434, B2 => 
                           n15198, ZN => n11956);
   U11553 : OAI22_X1 port map( A1 => n60294, A2 => n61034, B1 => n2433, B2 => 
                           n15198, ZN => n11957);
   U11554 : OAI22_X1 port map( A1 => n60294, A2 => n61048, B1 => n2432, B2 => 
                           n15198, ZN => n11958);
   U11555 : OAI22_X1 port map( A1 => n60294, A2 => n61062, B1 => n2431, B2 => 
                           n15198, ZN => n11959);
   U11556 : OAI22_X1 port map( A1 => n60294, A2 => n61076, B1 => n2430, B2 => 
                           n60290, ZN => n11960);
   U11557 : OAI22_X1 port map( A1 => n60295, A2 => n61090, B1 => n2429, B2 => 
                           n60290, ZN => n11961);
   U11558 : OAI22_X1 port map( A1 => n60295, A2 => n61104, B1 => n2428, B2 => 
                           n60290, ZN => n11962);
   U11559 : OAI22_X1 port map( A1 => n60295, A2 => n61118, B1 => n2427, B2 => 
                           n60290, ZN => n11963);
   U11560 : OAI22_X1 port map( A1 => n60295, A2 => n61132, B1 => n2426, B2 => 
                           n60290, ZN => n11964);
   U11561 : OAI22_X1 port map( A1 => n60282, A2 => n61971, B1 => n2425, B2 => 
                           n60281, ZN => n11909);
   U11562 : OAI22_X1 port map( A1 => n60282, A2 => n61985, B1 => n2424, B2 => 
                           n60281, ZN => n11910);
   U11563 : OAI22_X1 port map( A1 => n60282, A2 => n61999, B1 => n2423, B2 => 
                           n60281, ZN => n11911);
   U11564 : OAI22_X1 port map( A1 => n60282, A2 => n62013, B1 => n2422, B2 => 
                           n60281, ZN => n11912);
   U11565 : OAI22_X1 port map( A1 => n60282, A2 => n62027, B1 => n2421, B2 => 
                           n60281, ZN => n11913);
   U11566 : OAI22_X1 port map( A1 => n60283, A2 => n62041, B1 => n2420, B2 => 
                           n60281, ZN => n11914);
   U11567 : OAI22_X1 port map( A1 => n60283, A2 => n62055, B1 => n2419, B2 => 
                           n60281, ZN => n11915);
   U11568 : OAI22_X1 port map( A1 => n60283, A2 => n62069, B1 => n2418, B2 => 
                           n60281, ZN => n11916);
   U11569 : OAI22_X1 port map( A1 => n60283, A2 => n62083, B1 => n2417, B2 => 
                           n60281, ZN => n11917);
   U11570 : OAI22_X1 port map( A1 => n60283, A2 => n62097, B1 => n2416, B2 => 
                           n60281, ZN => n11918);
   U11571 : OAI22_X1 port map( A1 => n60284, A2 => n62111, B1 => n2415, B2 => 
                           n60281, ZN => n11919);
   U11572 : OAI22_X1 port map( A1 => n60284, A2 => n60964, B1 => n2414, B2 => 
                           n60281, ZN => n11920);
   U11573 : OAI22_X1 port map( A1 => n60284, A2 => n60978, B1 => n2413, B2 => 
                           n15199, ZN => n11921);
   U11574 : OAI22_X1 port map( A1 => n60284, A2 => n60992, B1 => n2412, B2 => 
                           n15199, ZN => n11922);
   U11575 : OAI22_X1 port map( A1 => n60284, A2 => n61006, B1 => n2411, B2 => 
                           n15199, ZN => n11923);
   U11576 : OAI22_X1 port map( A1 => n60285, A2 => n61020, B1 => n2410, B2 => 
                           n15199, ZN => n11924);
   U11577 : OAI22_X1 port map( A1 => n60285, A2 => n61034, B1 => n2409, B2 => 
                           n15199, ZN => n11925);
   U11578 : OAI22_X1 port map( A1 => n60285, A2 => n61048, B1 => n2408, B2 => 
                           n15199, ZN => n11926);
   U11579 : OAI22_X1 port map( A1 => n60285, A2 => n61062, B1 => n2407, B2 => 
                           n15199, ZN => n11927);
   U11580 : OAI22_X1 port map( A1 => n60285, A2 => n61076, B1 => n2406, B2 => 
                           n60281, ZN => n11928);
   U11581 : OAI22_X1 port map( A1 => n60286, A2 => n61090, B1 => n2405, B2 => 
                           n60281, ZN => n11929);
   U11582 : OAI22_X1 port map( A1 => n60286, A2 => n61104, B1 => n2404, B2 => 
                           n60281, ZN => n11930);
   U11583 : OAI22_X1 port map( A1 => n60286, A2 => n61118, B1 => n2403, B2 => 
                           n60281, ZN => n11931);
   U11584 : OAI22_X1 port map( A1 => n60286, A2 => n61132, B1 => n2402, B2 => 
                           n60281, ZN => n11932);
   U11585 : OAI22_X1 port map( A1 => n60255, A2 => n61971, B1 => n2225, B2 => 
                           n60254, ZN => n11813);
   U11586 : OAI22_X1 port map( A1 => n60255, A2 => n61985, B1 => n2224, B2 => 
                           n60254, ZN => n11814);
   U11587 : OAI22_X1 port map( A1 => n60255, A2 => n61999, B1 => n2223, B2 => 
                           n60254, ZN => n11815);
   U11588 : OAI22_X1 port map( A1 => n60255, A2 => n62013, B1 => n2222, B2 => 
                           n60254, ZN => n11816);
   U11589 : OAI22_X1 port map( A1 => n60255, A2 => n62027, B1 => n2221, B2 => 
                           n60254, ZN => n11817);
   U11590 : OAI22_X1 port map( A1 => n60256, A2 => n62041, B1 => n2212, B2 => 
                           n60254, ZN => n11818);
   U11591 : OAI22_X1 port map( A1 => n60256, A2 => n62055, B1 => n2211, B2 => 
                           n60254, ZN => n11819);
   U11592 : OAI22_X1 port map( A1 => n60256, A2 => n62069, B1 => n2210, B2 => 
                           n60254, ZN => n11820);
   U11593 : OAI22_X1 port map( A1 => n60256, A2 => n62083, B1 => n2209, B2 => 
                           n60254, ZN => n11821);
   U11594 : OAI22_X1 port map( A1 => n60256, A2 => n62097, B1 => n2208, B2 => 
                           n60254, ZN => n11822);
   U11595 : OAI22_X1 port map( A1 => n60257, A2 => n62111, B1 => n2207, B2 => 
                           n60254, ZN => n11823);
   U11596 : OAI22_X1 port map( A1 => n60257, A2 => n60964, B1 => n2206, B2 => 
                           n60254, ZN => n11824);
   U11597 : OAI22_X1 port map( A1 => n60257, A2 => n60978, B1 => n2205, B2 => 
                           n15202, ZN => n11825);
   U11598 : OAI22_X1 port map( A1 => n60257, A2 => n60992, B1 => n2204, B2 => 
                           n15202, ZN => n11826);
   U11599 : OAI22_X1 port map( A1 => n60257, A2 => n61006, B1 => n2203, B2 => 
                           n15202, ZN => n11827);
   U11600 : OAI22_X1 port map( A1 => n60258, A2 => n61020, B1 => n2202, B2 => 
                           n15202, ZN => n11828);
   U11601 : OAI22_X1 port map( A1 => n60258, A2 => n61034, B1 => n2201, B2 => 
                           n15202, ZN => n11829);
   U11602 : OAI22_X1 port map( A1 => n60258, A2 => n61048, B1 => n2200, B2 => 
                           n15202, ZN => n11830);
   U11603 : OAI22_X1 port map( A1 => n60258, A2 => n61062, B1 => n2199, B2 => 
                           n15202, ZN => n11831);
   U11604 : OAI22_X1 port map( A1 => n60258, A2 => n61076, B1 => n2198, B2 => 
                           n60254, ZN => n11832);
   U11605 : OAI22_X1 port map( A1 => n60259, A2 => n61090, B1 => n2197, B2 => 
                           n60254, ZN => n11833);
   U11606 : OAI22_X1 port map( A1 => n60259, A2 => n61104, B1 => n2196, B2 => 
                           n60254, ZN => n11834);
   U11607 : OAI22_X1 port map( A1 => n60259, A2 => n61118, B1 => n2195, B2 => 
                           n60254, ZN => n11835);
   U11608 : OAI22_X1 port map( A1 => n60259, A2 => n61132, B1 => n2194, B2 => 
                           n60254, ZN => n11836);
   U11609 : OAI22_X1 port map( A1 => n60246, A2 => n61971, B1 => n2193, B2 => 
                           n60245, ZN => n11781);
   U11610 : OAI22_X1 port map( A1 => n60246, A2 => n61985, B1 => n2192, B2 => 
                           n60245, ZN => n11782);
   U11611 : OAI22_X1 port map( A1 => n60246, A2 => n61999, B1 => n2191, B2 => 
                           n60245, ZN => n11783);
   U11612 : OAI22_X1 port map( A1 => n60246, A2 => n62013, B1 => n2190, B2 => 
                           n60245, ZN => n11784);
   U11613 : OAI22_X1 port map( A1 => n60246, A2 => n62027, B1 => n2189, B2 => 
                           n60245, ZN => n11785);
   U11614 : OAI22_X1 port map( A1 => n60247, A2 => n62041, B1 => n2188, B2 => 
                           n60245, ZN => n11786);
   U11615 : OAI22_X1 port map( A1 => n60247, A2 => n62055, B1 => n2187, B2 => 
                           n60245, ZN => n11787);
   U11616 : OAI22_X1 port map( A1 => n60247, A2 => n62069, B1 => n2186, B2 => 
                           n60245, ZN => n11788);
   U11617 : OAI22_X1 port map( A1 => n60247, A2 => n62083, B1 => n2185, B2 => 
                           n60245, ZN => n11789);
   U11618 : OAI22_X1 port map( A1 => n60247, A2 => n62097, B1 => n2184, B2 => 
                           n60245, ZN => n11790);
   U11619 : OAI22_X1 port map( A1 => n60248, A2 => n62111, B1 => n2183, B2 => 
                           n60245, ZN => n11791);
   U11620 : OAI22_X1 port map( A1 => n60248, A2 => n60964, B1 => n2182, B2 => 
                           n60245, ZN => n11792);
   U11621 : OAI22_X1 port map( A1 => n60248, A2 => n60978, B1 => n2181, B2 => 
                           n15211, ZN => n11793);
   U11622 : OAI22_X1 port map( A1 => n60248, A2 => n60992, B1 => n2180, B2 => 
                           n15211, ZN => n11794);
   U11623 : OAI22_X1 port map( A1 => n60248, A2 => n61006, B1 => n2179, B2 => 
                           n15211, ZN => n11795);
   U11624 : OAI22_X1 port map( A1 => n60249, A2 => n61020, B1 => n2178, B2 => 
                           n15211, ZN => n11796);
   U11625 : OAI22_X1 port map( A1 => n60249, A2 => n61034, B1 => n2177, B2 => 
                           n15211, ZN => n11797);
   U11626 : OAI22_X1 port map( A1 => n60249, A2 => n61048, B1 => n2176, B2 => 
                           n15211, ZN => n11798);
   U11627 : OAI22_X1 port map( A1 => n60249, A2 => n61062, B1 => n2175, B2 => 
                           n15211, ZN => n11799);
   U11628 : OAI22_X1 port map( A1 => n60249, A2 => n61076, B1 => n2174, B2 => 
                           n60245, ZN => n11800);
   U11629 : OAI22_X1 port map( A1 => n60250, A2 => n61090, B1 => n2173, B2 => 
                           n60245, ZN => n11801);
   U11630 : OAI22_X1 port map( A1 => n60250, A2 => n61104, B1 => n2172, B2 => 
                           n60245, ZN => n11802);
   U11631 : OAI22_X1 port map( A1 => n60250, A2 => n61118, B1 => n2171, B2 => 
                           n60245, ZN => n11803);
   U11632 : OAI22_X1 port map( A1 => n60250, A2 => n61132, B1 => n2170, B2 => 
                           n60245, ZN => n11804);
   U11633 : OAI22_X1 port map( A1 => n60219, A2 => n61971, B1 => n2121, B2 => 
                           n60218, ZN => n11685);
   U11634 : OAI22_X1 port map( A1 => n60219, A2 => n61985, B1 => n2120, B2 => 
                           n60218, ZN => n11686);
   U11635 : OAI22_X1 port map( A1 => n60219, A2 => n61999, B1 => n2119, B2 => 
                           n60218, ZN => n11687);
   U11636 : OAI22_X1 port map( A1 => n60219, A2 => n62013, B1 => n2118, B2 => 
                           n60218, ZN => n11688);
   U11637 : OAI22_X1 port map( A1 => n60219, A2 => n62027, B1 => n2117, B2 => 
                           n60218, ZN => n11689);
   U11638 : OAI22_X1 port map( A1 => n60220, A2 => n62041, B1 => n2116, B2 => 
                           n60218, ZN => n11690);
   U11639 : OAI22_X1 port map( A1 => n60220, A2 => n62055, B1 => n2115, B2 => 
                           n60218, ZN => n11691);
   U11640 : OAI22_X1 port map( A1 => n60220, A2 => n62069, B1 => n2114, B2 => 
                           n60218, ZN => n11692);
   U11641 : OAI22_X1 port map( A1 => n60220, A2 => n62083, B1 => n2113, B2 => 
                           n60218, ZN => n11693);
   U11642 : OAI22_X1 port map( A1 => n60220, A2 => n62097, B1 => n2112, B2 => 
                           n60218, ZN => n11694);
   U11643 : OAI22_X1 port map( A1 => n60221, A2 => n62111, B1 => n2111, B2 => 
                           n60218, ZN => n11695);
   U11644 : OAI22_X1 port map( A1 => n60221, A2 => n60964, B1 => n2110, B2 => 
                           n60218, ZN => n11696);
   U11645 : OAI22_X1 port map( A1 => n60221, A2 => n60978, B1 => n2109, B2 => 
                           n15215, ZN => n11697);
   U11646 : OAI22_X1 port map( A1 => n60221, A2 => n60992, B1 => n2108, B2 => 
                           n15215, ZN => n11698);
   U11647 : OAI22_X1 port map( A1 => n60221, A2 => n61006, B1 => n2107, B2 => 
                           n15215, ZN => n11699);
   U11648 : OAI22_X1 port map( A1 => n60222, A2 => n61020, B1 => n2106, B2 => 
                           n15215, ZN => n11700);
   U11649 : OAI22_X1 port map( A1 => n60222, A2 => n61034, B1 => n2105, B2 => 
                           n15215, ZN => n11701);
   U11650 : OAI22_X1 port map( A1 => n60222, A2 => n61048, B1 => n2104, B2 => 
                           n15215, ZN => n11702);
   U11651 : OAI22_X1 port map( A1 => n60222, A2 => n61062, B1 => n2103, B2 => 
                           n15215, ZN => n11703);
   U11652 : OAI22_X1 port map( A1 => n60222, A2 => n61076, B1 => n2102, B2 => 
                           n60218, ZN => n11704);
   U11653 : OAI22_X1 port map( A1 => n60223, A2 => n61090, B1 => n2101, B2 => 
                           n60218, ZN => n11705);
   U11654 : OAI22_X1 port map( A1 => n60223, A2 => n61104, B1 => n2100, B2 => 
                           n60218, ZN => n11706);
   U11655 : OAI22_X1 port map( A1 => n60223, A2 => n61118, B1 => n2099, B2 => 
                           n60218, ZN => n11707);
   U11656 : OAI22_X1 port map( A1 => n60223, A2 => n61132, B1 => n2098, B2 => 
                           n60218, ZN => n11708);
   U11657 : OAI22_X1 port map( A1 => n60201, A2 => n61972, B1 => n2069, B2 => 
                           n60200, ZN => n11621);
   U11658 : OAI22_X1 port map( A1 => n60201, A2 => n61986, B1 => n2068, B2 => 
                           n60200, ZN => n11622);
   U11659 : OAI22_X1 port map( A1 => n60201, A2 => n62000, B1 => n2067, B2 => 
                           n60200, ZN => n11623);
   U11660 : OAI22_X1 port map( A1 => n60201, A2 => n62014, B1 => n2066, B2 => 
                           n60200, ZN => n11624);
   U11661 : OAI22_X1 port map( A1 => n60201, A2 => n62028, B1 => n2065, B2 => 
                           n60200, ZN => n11625);
   U11662 : OAI22_X1 port map( A1 => n60202, A2 => n62042, B1 => n2064, B2 => 
                           n60200, ZN => n11626);
   U11663 : OAI22_X1 port map( A1 => n60202, A2 => n62056, B1 => n2063, B2 => 
                           n60200, ZN => n11627);
   U11664 : OAI22_X1 port map( A1 => n60202, A2 => n62070, B1 => n2062, B2 => 
                           n60200, ZN => n11628);
   U11665 : OAI22_X1 port map( A1 => n60202, A2 => n62084, B1 => n2061, B2 => 
                           n60200, ZN => n11629);
   U11666 : OAI22_X1 port map( A1 => n60202, A2 => n62098, B1 => n2060, B2 => 
                           n60200, ZN => n11630);
   U11667 : OAI22_X1 port map( A1 => n60203, A2 => n62112, B1 => n2059, B2 => 
                           n60200, ZN => n11631);
   U11668 : OAI22_X1 port map( A1 => n60203, A2 => n60965, B1 => n2058, B2 => 
                           n60200, ZN => n11632);
   U11669 : OAI22_X1 port map( A1 => n60203, A2 => n60979, B1 => n2057, B2 => 
                           n15217, ZN => n11633);
   U11670 : OAI22_X1 port map( A1 => n60203, A2 => n60993, B1 => n2056, B2 => 
                           n15217, ZN => n11634);
   U11671 : OAI22_X1 port map( A1 => n60203, A2 => n61007, B1 => n2055, B2 => 
                           n15217, ZN => n11635);
   U11672 : OAI22_X1 port map( A1 => n60204, A2 => n61021, B1 => n2054, B2 => 
                           n15217, ZN => n11636);
   U11673 : OAI22_X1 port map( A1 => n60204, A2 => n61035, B1 => n2053, B2 => 
                           n15217, ZN => n11637);
   U11674 : OAI22_X1 port map( A1 => n60204, A2 => n61049, B1 => n2052, B2 => 
                           n15217, ZN => n11638);
   U11675 : OAI22_X1 port map( A1 => n60204, A2 => n61063, B1 => n2051, B2 => 
                           n15217, ZN => n11639);
   U11676 : OAI22_X1 port map( A1 => n60204, A2 => n61077, B1 => n2050, B2 => 
                           n60200, ZN => n11640);
   U11677 : OAI22_X1 port map( A1 => n60205, A2 => n61091, B1 => n2049, B2 => 
                           n60200, ZN => n11641);
   U11678 : OAI22_X1 port map( A1 => n60205, A2 => n61105, B1 => n2048, B2 => 
                           n60200, ZN => n11642);
   U11679 : OAI22_X1 port map( A1 => n60205, A2 => n61119, B1 => n2047, B2 => 
                           n60200, ZN => n11643);
   U11680 : OAI22_X1 port map( A1 => n60205, A2 => n61133, B1 => n2046, B2 => 
                           n60200, ZN => n11644);
   U11681 : OAI22_X1 port map( A1 => n60165, A2 => n61972, B1 => n1973, B2 => 
                           n60164, ZN => n11493);
   U11682 : OAI22_X1 port map( A1 => n60165, A2 => n61986, B1 => n1972, B2 => 
                           n60164, ZN => n11494);
   U11683 : OAI22_X1 port map( A1 => n60165, A2 => n62000, B1 => n1971, B2 => 
                           n60164, ZN => n11495);
   U11684 : OAI22_X1 port map( A1 => n60165, A2 => n62014, B1 => n1970, B2 => 
                           n60164, ZN => n11496);
   U11685 : OAI22_X1 port map( A1 => n60165, A2 => n62028, B1 => n1969, B2 => 
                           n60164, ZN => n11497);
   U11686 : OAI22_X1 port map( A1 => n60166, A2 => n62042, B1 => n1968, B2 => 
                           n60164, ZN => n11498);
   U11687 : OAI22_X1 port map( A1 => n60166, A2 => n62056, B1 => n1967, B2 => 
                           n60164, ZN => n11499);
   U11688 : OAI22_X1 port map( A1 => n60166, A2 => n62070, B1 => n1966, B2 => 
                           n60164, ZN => n11500);
   U11689 : OAI22_X1 port map( A1 => n60166, A2 => n62084, B1 => n1965, B2 => 
                           n60164, ZN => n11501);
   U11690 : OAI22_X1 port map( A1 => n60166, A2 => n62098, B1 => n1964, B2 => 
                           n60164, ZN => n11502);
   U11691 : OAI22_X1 port map( A1 => n60167, A2 => n62112, B1 => n1963, B2 => 
                           n60164, ZN => n11503);
   U11692 : OAI22_X1 port map( A1 => n60167, A2 => n60965, B1 => n1962, B2 => 
                           n60164, ZN => n11504);
   U11693 : OAI22_X1 port map( A1 => n60167, A2 => n60979, B1 => n1961, B2 => 
                           n15221, ZN => n11505);
   U11694 : OAI22_X1 port map( A1 => n60167, A2 => n60993, B1 => n1960, B2 => 
                           n15221, ZN => n11506);
   U11695 : OAI22_X1 port map( A1 => n60167, A2 => n61007, B1 => n1959, B2 => 
                           n15221, ZN => n11507);
   U11696 : OAI22_X1 port map( A1 => n60168, A2 => n61021, B1 => n1958, B2 => 
                           n15221, ZN => n11508);
   U11697 : OAI22_X1 port map( A1 => n60168, A2 => n61035, B1 => n1957, B2 => 
                           n15221, ZN => n11509);
   U11698 : OAI22_X1 port map( A1 => n60168, A2 => n61049, B1 => n1956, B2 => 
                           n15221, ZN => n11510);
   U11699 : OAI22_X1 port map( A1 => n60168, A2 => n61063, B1 => n1955, B2 => 
                           n15221, ZN => n11511);
   U11700 : OAI22_X1 port map( A1 => n60168, A2 => n61077, B1 => n1954, B2 => 
                           n60164, ZN => n11512);
   U11701 : OAI22_X1 port map( A1 => n60169, A2 => n61091, B1 => n1953, B2 => 
                           n60164, ZN => n11513);
   U11702 : OAI22_X1 port map( A1 => n60169, A2 => n61105, B1 => n1952, B2 => 
                           n60164, ZN => n11514);
   U11703 : OAI22_X1 port map( A1 => n60169, A2 => n61119, B1 => n1951, B2 => 
                           n60164, ZN => n11515);
   U11704 : OAI22_X1 port map( A1 => n60169, A2 => n61133, B1 => n1950, B2 => 
                           n60164, ZN => n11516);
   U11705 : OAI22_X1 port map( A1 => n60138, A2 => n61972, B1 => n212, B2 => 
                           n60137, ZN => n11397);
   U11706 : OAI22_X1 port map( A1 => n60138, A2 => n61986, B1 => n211, B2 => 
                           n60137, ZN => n11398);
   U11707 : OAI22_X1 port map( A1 => n60138, A2 => n62000, B1 => n210, B2 => 
                           n60137, ZN => n11399);
   U11708 : OAI22_X1 port map( A1 => n60138, A2 => n62014, B1 => n209, B2 => 
                           n60137, ZN => n11400);
   U11709 : OAI22_X1 port map( A1 => n60138, A2 => n62028, B1 => n208, B2 => 
                           n60137, ZN => n11401);
   U11710 : OAI22_X1 port map( A1 => n60139, A2 => n62042, B1 => n207, B2 => 
                           n60137, ZN => n11402);
   U11711 : OAI22_X1 port map( A1 => n60139, A2 => n62056, B1 => n206, B2 => 
                           n60137, ZN => n11403);
   U11712 : OAI22_X1 port map( A1 => n60139, A2 => n62070, B1 => n205, B2 => 
                           n60137, ZN => n11404);
   U11713 : OAI22_X1 port map( A1 => n60139, A2 => n62084, B1 => n204, B2 => 
                           n60137, ZN => n11405);
   U11714 : OAI22_X1 port map( A1 => n60139, A2 => n62098, B1 => n203, B2 => 
                           n60137, ZN => n11406);
   U11715 : OAI22_X1 port map( A1 => n60140, A2 => n62112, B1 => n202, B2 => 
                           n60137, ZN => n11407);
   U11716 : OAI22_X1 port map( A1 => n60140, A2 => n60965, B1 => n201, B2 => 
                           n60137, ZN => n11408);
   U11717 : OAI22_X1 port map( A1 => n60140, A2 => n60979, B1 => n200, B2 => 
                           n15224, ZN => n11409);
   U11718 : OAI22_X1 port map( A1 => n60140, A2 => n60993, B1 => n199, B2 => 
                           n15224, ZN => n11410);
   U11719 : OAI22_X1 port map( A1 => n60140, A2 => n61007, B1 => n198, B2 => 
                           n15224, ZN => n11411);
   U11720 : OAI22_X1 port map( A1 => n60141, A2 => n61021, B1 => n197, B2 => 
                           n15224, ZN => n11412);
   U11721 : OAI22_X1 port map( A1 => n60141, A2 => n61035, B1 => n196, B2 => 
                           n15224, ZN => n11413);
   U11722 : OAI22_X1 port map( A1 => n60141, A2 => n61049, B1 => n195, B2 => 
                           n15224, ZN => n11414);
   U11723 : OAI22_X1 port map( A1 => n60141, A2 => n61063, B1 => n194, B2 => 
                           n15224, ZN => n11415);
   U11724 : OAI22_X1 port map( A1 => n60141, A2 => n61077, B1 => n193, B2 => 
                           n60137, ZN => n11416);
   U11725 : OAI22_X1 port map( A1 => n60142, A2 => n61091, B1 => n192, B2 => 
                           n60137, ZN => n11417);
   U11726 : OAI22_X1 port map( A1 => n60142, A2 => n61105, B1 => n191, B2 => 
                           n60137, ZN => n11418);
   U11727 : OAI22_X1 port map( A1 => n60142, A2 => n61119, B1 => n190, B2 => 
                           n60137, ZN => n11419);
   U11728 : OAI22_X1 port map( A1 => n60142, A2 => n61133, B1 => n189, B2 => 
                           n60137, ZN => n11420);
   U11729 : OAI22_X1 port map( A1 => n60114, A2 => n61049, B1 => n2651, B2 => 
                           n15227, ZN => n11318);
   U11730 : OAI22_X1 port map( A1 => n60114, A2 => n61063, B1 => n2650, B2 => 
                           n15227, ZN => n11319);
   U11731 : OAI22_X1 port map( A1 => n60114, A2 => n61077, B1 => n2649, B2 => 
                           n60110, ZN => n11320);
   U11732 : OAI22_X1 port map( A1 => n60115, A2 => n61091, B1 => n2648, B2 => 
                           n60110, ZN => n11321);
   U11733 : OAI22_X1 port map( A1 => n60115, A2 => n61105, B1 => n2647, B2 => 
                           n60110, ZN => n11322);
   U11734 : OAI22_X1 port map( A1 => n60115, A2 => n61119, B1 => n2646, B2 => 
                           n60110, ZN => n11323);
   U11735 : OAI22_X1 port map( A1 => n60115, A2 => n61133, B1 => n2645, B2 => 
                           n60110, ZN => n11324);
   U11736 : OAI22_X1 port map( A1 => n60786, A2 => n61966, B1 => n3456, B2 => 
                           n60785, ZN => n13701);
   U11737 : OAI22_X1 port map( A1 => n60786, A2 => n61980, B1 => n3455, B2 => 
                           n60785, ZN => n13702);
   U11738 : OAI22_X1 port map( A1 => n60786, A2 => n61994, B1 => n3454, B2 => 
                           n60785, ZN => n13703);
   U11739 : OAI22_X1 port map( A1 => n60786, A2 => n62008, B1 => n3453, B2 => 
                           n60785, ZN => n13704);
   U11740 : OAI22_X1 port map( A1 => n60786, A2 => n62022, B1 => n3452, B2 => 
                           n60785, ZN => n13705);
   U11741 : OAI22_X1 port map( A1 => n60787, A2 => n62036, B1 => n3451, B2 => 
                           n60785, ZN => n13706);
   U11742 : OAI22_X1 port map( A1 => n60787, A2 => n62050, B1 => n3450, B2 => 
                           n60785, ZN => n13707);
   U11743 : OAI22_X1 port map( A1 => n60787, A2 => n62064, B1 => n3449, B2 => 
                           n60785, ZN => n13708);
   U11744 : OAI22_X1 port map( A1 => n60787, A2 => n62078, B1 => n3448, B2 => 
                           n60785, ZN => n13709);
   U11745 : OAI22_X1 port map( A1 => n60787, A2 => n62092, B1 => n3447, B2 => 
                           n60785, ZN => n13710);
   U11746 : OAI22_X1 port map( A1 => n60788, A2 => n62106, B1 => n3446, B2 => 
                           n60785, ZN => n13711);
   U11747 : OAI22_X1 port map( A1 => n60788, A2 => n60959, B1 => n3445, B2 => 
                           n60785, ZN => n13712);
   U11748 : OAI22_X1 port map( A1 => n60788, A2 => n60973, B1 => n3444, B2 => 
                           n15132, ZN => n13713);
   U11749 : OAI22_X1 port map( A1 => n60788, A2 => n60987, B1 => n3443, B2 => 
                           n15132, ZN => n13714);
   U11750 : OAI22_X1 port map( A1 => n60788, A2 => n61001, B1 => n3442, B2 => 
                           n15132, ZN => n13715);
   U11751 : OAI22_X1 port map( A1 => n60789, A2 => n61015, B1 => n3441, B2 => 
                           n15132, ZN => n13716);
   U11752 : OAI22_X1 port map( A1 => n60789, A2 => n61029, B1 => n3440, B2 => 
                           n15132, ZN => n13717);
   U11753 : OAI22_X1 port map( A1 => n60789, A2 => n61043, B1 => n3439, B2 => 
                           n15132, ZN => n13718);
   U11754 : OAI22_X1 port map( A1 => n60789, A2 => n61057, B1 => n3438, B2 => 
                           n15132, ZN => n13719);
   U11755 : OAI22_X1 port map( A1 => n60789, A2 => n61071, B1 => n3437, B2 => 
                           n60785, ZN => n13720);
   U11756 : OAI22_X1 port map( A1 => n60790, A2 => n61085, B1 => n3436, B2 => 
                           n60785, ZN => n13721);
   U11757 : OAI22_X1 port map( A1 => n60790, A2 => n61099, B1 => n3435, B2 => 
                           n60785, ZN => n13722);
   U11758 : OAI22_X1 port map( A1 => n60790, A2 => n61113, B1 => n3434, B2 => 
                           n60785, ZN => n13723);
   U11759 : OAI22_X1 port map( A1 => n60790, A2 => n61127, B1 => n3433, B2 => 
                           n60785, ZN => n13724);
   U11760 : OAI22_X1 port map( A1 => n60768, A2 => n61966, B1 => n1588, B2 => 
                           n60767, ZN => n13637);
   U11761 : OAI22_X1 port map( A1 => n60768, A2 => n61980, B1 => n1587, B2 => 
                           n60767, ZN => n13638);
   U11762 : OAI22_X1 port map( A1 => n60768, A2 => n61994, B1 => n1586, B2 => 
                           n60767, ZN => n13639);
   U11763 : OAI22_X1 port map( A1 => n60768, A2 => n62008, B1 => n1585, B2 => 
                           n60767, ZN => n13640);
   U11764 : OAI22_X1 port map( A1 => n60768, A2 => n62022, B1 => n1584, B2 => 
                           n60767, ZN => n13641);
   U11765 : OAI22_X1 port map( A1 => n60769, A2 => n62036, B1 => n1583, B2 => 
                           n60767, ZN => n13642);
   U11766 : OAI22_X1 port map( A1 => n60769, A2 => n62050, B1 => n1582, B2 => 
                           n60767, ZN => n13643);
   U11767 : OAI22_X1 port map( A1 => n60769, A2 => n62064, B1 => n1581, B2 => 
                           n60767, ZN => n13644);
   U11768 : OAI22_X1 port map( A1 => n60769, A2 => n62078, B1 => n1580, B2 => 
                           n60767, ZN => n13645);
   U11769 : OAI22_X1 port map( A1 => n60769, A2 => n62092, B1 => n1579, B2 => 
                           n60767, ZN => n13646);
   U11770 : OAI22_X1 port map( A1 => n60770, A2 => n62106, B1 => n1578, B2 => 
                           n60767, ZN => n13647);
   U11771 : OAI22_X1 port map( A1 => n60770, A2 => n60959, B1 => n1577, B2 => 
                           n60767, ZN => n13648);
   U11772 : OAI22_X1 port map( A1 => n60770, A2 => n60973, B1 => n1576, B2 => 
                           n60767, ZN => n13649);
   U11773 : OAI22_X1 port map( A1 => n60770, A2 => n60987, B1 => n1575, B2 => 
                           n60767, ZN => n13650);
   U11774 : OAI22_X1 port map( A1 => n60750, A2 => n61966, B1 => n1704, B2 => 
                           n60749, ZN => n13573);
   U11775 : OAI22_X1 port map( A1 => n60750, A2 => n61980, B1 => n1703, B2 => 
                           n60749, ZN => n13574);
   U11776 : OAI22_X1 port map( A1 => n60750, A2 => n61994, B1 => n1702, B2 => 
                           n60749, ZN => n13575);
   U11777 : OAI22_X1 port map( A1 => n60750, A2 => n62008, B1 => n1701, B2 => 
                           n60749, ZN => n13576);
   U11778 : OAI22_X1 port map( A1 => n60750, A2 => n62022, B1 => n1700, B2 => 
                           n60749, ZN => n13577);
   U11779 : OAI22_X1 port map( A1 => n60751, A2 => n62036, B1 => n1699, B2 => 
                           n60749, ZN => n13578);
   U11780 : OAI22_X1 port map( A1 => n60751, A2 => n62050, B1 => n1698, B2 => 
                           n60749, ZN => n13579);
   U11781 : OAI22_X1 port map( A1 => n60751, A2 => n62064, B1 => n1697, B2 => 
                           n60749, ZN => n13580);
   U11782 : OAI22_X1 port map( A1 => n60751, A2 => n62078, B1 => n1696, B2 => 
                           n60749, ZN => n13581);
   U11783 : OAI22_X1 port map( A1 => n60751, A2 => n62092, B1 => n1695, B2 => 
                           n60749, ZN => n13582);
   U11784 : OAI22_X1 port map( A1 => n60752, A2 => n62106, B1 => n1694, B2 => 
                           n60749, ZN => n13583);
   U11785 : OAI22_X1 port map( A1 => n60752, A2 => n60959, B1 => n1693, B2 => 
                           n60749, ZN => n13584);
   U11786 : OAI22_X1 port map( A1 => n60752, A2 => n60973, B1 => n1668, B2 => 
                           n15136, ZN => n13585);
   U11787 : OAI22_X1 port map( A1 => n60752, A2 => n60987, B1 => n1667, B2 => 
                           n15136, ZN => n13586);
   U11788 : OAI22_X1 port map( A1 => n60752, A2 => n61001, B1 => n1666, B2 => 
                           n15136, ZN => n13587);
   U11789 : OAI22_X1 port map( A1 => n60753, A2 => n61015, B1 => n1665, B2 => 
                           n15136, ZN => n13588);
   U11790 : OAI22_X1 port map( A1 => n60753, A2 => n61029, B1 => n1664, B2 => 
                           n15136, ZN => n13589);
   U11791 : OAI22_X1 port map( A1 => n60753, A2 => n61043, B1 => n1663, B2 => 
                           n15136, ZN => n13590);
   U11792 : OAI22_X1 port map( A1 => n60753, A2 => n61057, B1 => n1662, B2 => 
                           n15136, ZN => n13591);
   U11793 : OAI22_X1 port map( A1 => n60753, A2 => n61071, B1 => n1661, B2 => 
                           n60749, ZN => n13592);
   U11794 : OAI22_X1 port map( A1 => n60754, A2 => n61085, B1 => n1660, B2 => 
                           n60749, ZN => n13593);
   U11795 : OAI22_X1 port map( A1 => n60754, A2 => n61099, B1 => n1659, B2 => 
                           n60749, ZN => n13594);
   U11796 : OAI22_X1 port map( A1 => n60754, A2 => n61113, B1 => n1658, B2 => 
                           n60749, ZN => n13595);
   U11797 : OAI22_X1 port map( A1 => n60754, A2 => n61127, B1 => n1657, B2 => 
                           n60749, ZN => n13596);
   U11798 : OAI22_X1 port map( A1 => n60741, A2 => n61967, B1 => n1656, B2 => 
                           n60740, ZN => n13541);
   U11799 : OAI22_X1 port map( A1 => n60741, A2 => n61981, B1 => n1655, B2 => 
                           n60740, ZN => n13542);
   U11800 : OAI22_X1 port map( A1 => n60741, A2 => n61995, B1 => n1654, B2 => 
                           n60740, ZN => n13543);
   U11801 : OAI22_X1 port map( A1 => n60741, A2 => n62009, B1 => n1653, B2 => 
                           n60740, ZN => n13544);
   U11802 : OAI22_X1 port map( A1 => n60741, A2 => n62023, B1 => n1652, B2 => 
                           n60740, ZN => n13545);
   U11803 : OAI22_X1 port map( A1 => n60742, A2 => n62037, B1 => n1651, B2 => 
                           n60740, ZN => n13546);
   U11804 : OAI22_X1 port map( A1 => n60742, A2 => n62051, B1 => n1650, B2 => 
                           n60740, ZN => n13547);
   U11805 : OAI22_X1 port map( A1 => n60742, A2 => n62065, B1 => n1649, B2 => 
                           n60740, ZN => n13548);
   U11806 : OAI22_X1 port map( A1 => n60742, A2 => n62079, B1 => n1648, B2 => 
                           n60740, ZN => n13549);
   U11807 : OAI22_X1 port map( A1 => n60742, A2 => n62093, B1 => n1647, B2 => 
                           n60740, ZN => n13550);
   U11808 : OAI22_X1 port map( A1 => n60743, A2 => n62107, B1 => n1630, B2 => 
                           n60740, ZN => n13551);
   U11809 : OAI22_X1 port map( A1 => n60743, A2 => n60960, B1 => n1629, B2 => 
                           n60740, ZN => n13552);
   U11810 : OAI22_X1 port map( A1 => n60743, A2 => n60974, B1 => n1628, B2 => 
                           n15137, ZN => n13553);
   U11811 : OAI22_X1 port map( A1 => n60743, A2 => n60988, B1 => n1627, B2 => 
                           n15137, ZN => n13554);
   U11812 : OAI22_X1 port map( A1 => n60743, A2 => n61002, B1 => n1626, B2 => 
                           n15137, ZN => n13555);
   U11813 : OAI22_X1 port map( A1 => n60744, A2 => n61016, B1 => n1625, B2 => 
                           n15137, ZN => n13556);
   U11814 : OAI22_X1 port map( A1 => n60744, A2 => n61030, B1 => n1624, B2 => 
                           n15137, ZN => n13557);
   U11815 : OAI22_X1 port map( A1 => n60744, A2 => n61044, B1 => n1623, B2 => 
                           n15137, ZN => n13558);
   U11816 : OAI22_X1 port map( A1 => n60744, A2 => n61058, B1 => n1622, B2 => 
                           n15137, ZN => n13559);
   U11817 : OAI22_X1 port map( A1 => n60744, A2 => n61072, B1 => n1621, B2 => 
                           n60740, ZN => n13560);
   U11818 : OAI22_X1 port map( A1 => n60745, A2 => n61086, B1 => n1620, B2 => 
                           n60740, ZN => n13561);
   U11819 : OAI22_X1 port map( A1 => n60745, A2 => n61100, B1 => n1619, B2 => 
                           n60740, ZN => n13562);
   U11820 : OAI22_X1 port map( A1 => n60745, A2 => n61114, B1 => n1618, B2 => 
                           n60740, ZN => n13563);
   U11821 : OAI22_X1 port map( A1 => n60745, A2 => n61128, B1 => n1617, B2 => 
                           n60740, ZN => n13564);
   U11822 : OAI22_X1 port map( A1 => n60714, A2 => n62023, B1 => n1507, B2 => 
                           n60713, ZN => n13449);
   U11823 : OAI22_X1 port map( A1 => n60678, A2 => n61967, B1 => n1458, B2 => 
                           n60677, ZN => n13317);
   U11824 : OAI22_X1 port map( A1 => n60678, A2 => n61981, B1 => n1457, B2 => 
                           n60677, ZN => n13318);
   U11825 : OAI22_X1 port map( A1 => n60678, A2 => n61995, B1 => n1456, B2 => 
                           n60677, ZN => n13319);
   U11826 : OAI22_X1 port map( A1 => n60678, A2 => n62009, B1 => n1455, B2 => 
                           n60677, ZN => n13320);
   U11827 : OAI22_X1 port map( A1 => n60678, A2 => n62023, B1 => n1454, B2 => 
                           n60677, ZN => n13321);
   U11828 : OAI22_X1 port map( A1 => n60679, A2 => n62037, B1 => n1453, B2 => 
                           n60677, ZN => n13322);
   U11829 : OAI22_X1 port map( A1 => n60679, A2 => n62051, B1 => n1452, B2 => 
                           n60677, ZN => n13323);
   U11830 : OAI22_X1 port map( A1 => n60679, A2 => n62065, B1 => n1451, B2 => 
                           n60677, ZN => n13324);
   U11831 : OAI22_X1 port map( A1 => n60679, A2 => n62079, B1 => n1450, B2 => 
                           n60677, ZN => n13325);
   U11832 : OAI22_X1 port map( A1 => n60679, A2 => n62093, B1 => n1449, B2 => 
                           n60677, ZN => n13326);
   U11833 : OAI22_X1 port map( A1 => n60680, A2 => n62107, B1 => n1448, B2 => 
                           n60677, ZN => n13327);
   U11834 : OAI22_X1 port map( A1 => n60680, A2 => n60960, B1 => n1447, B2 => 
                           n60677, ZN => n13328);
   U11835 : OAI22_X1 port map( A1 => n60680, A2 => n60974, B1 => n1446, B2 => 
                           n15144, ZN => n13329);
   U11836 : OAI22_X1 port map( A1 => n60680, A2 => n60988, B1 => n1445, B2 => 
                           n15144, ZN => n13330);
   U11837 : OAI22_X1 port map( A1 => n60680, A2 => n61002, B1 => n1444, B2 => 
                           n15144, ZN => n13331);
   U11838 : OAI22_X1 port map( A1 => n60681, A2 => n61016, B1 => n1443, B2 => 
                           n15144, ZN => n13332);
   U11839 : OAI22_X1 port map( A1 => n60681, A2 => n61030, B1 => n1442, B2 => 
                           n15144, ZN => n13333);
   U11840 : OAI22_X1 port map( A1 => n60681, A2 => n61044, B1 => n1441, B2 => 
                           n15144, ZN => n13334);
   U11841 : OAI22_X1 port map( A1 => n60681, A2 => n61058, B1 => n1440, B2 => 
                           n15144, ZN => n13335);
   U11842 : OAI22_X1 port map( A1 => n60681, A2 => n61072, B1 => n1439, B2 => 
                           n60677, ZN => n13336);
   U11843 : OAI22_X1 port map( A1 => n60682, A2 => n61086, B1 => n1438, B2 => 
                           n60677, ZN => n13337);
   U11844 : OAI22_X1 port map( A1 => n60682, A2 => n61100, B1 => n1437, B2 => 
                           n60677, ZN => n13338);
   U11845 : OAI22_X1 port map( A1 => n60682, A2 => n61114, B1 => n1436, B2 => 
                           n60677, ZN => n13339);
   U11846 : OAI22_X1 port map( A1 => n60682, A2 => n61128, B1 => n1435, B2 => 
                           n60677, ZN => n13340);
   U11847 : OAI22_X1 port map( A1 => n59805, A2 => n61975, B1 => n1434, B2 => 
                           n59804, ZN => n10213);
   U11848 : OAI22_X1 port map( A1 => n59805, A2 => n61989, B1 => n1433, B2 => 
                           n59804, ZN => n10214);
   U11849 : OAI22_X1 port map( A1 => n59805, A2 => n62003, B1 => n1432, B2 => 
                           n59804, ZN => n10215);
   U11850 : OAI22_X1 port map( A1 => n59805, A2 => n62017, B1 => n1431, B2 => 
                           n59804, ZN => n10216);
   U11851 : OAI22_X1 port map( A1 => n59805, A2 => n62031, B1 => n1430, B2 => 
                           n59804, ZN => n10217);
   U11852 : OAI22_X1 port map( A1 => n59806, A2 => n62045, B1 => n1429, B2 => 
                           n59804, ZN => n10218);
   U11853 : OAI22_X1 port map( A1 => n59806, A2 => n62059, B1 => n1428, B2 => 
                           n59804, ZN => n10219);
   U11854 : OAI22_X1 port map( A1 => n59806, A2 => n62073, B1 => n1427, B2 => 
                           n59804, ZN => n10220);
   U11855 : OAI22_X1 port map( A1 => n59806, A2 => n62087, B1 => n1426, B2 => 
                           n59804, ZN => n10221);
   U11856 : OAI22_X1 port map( A1 => n59806, A2 => n62101, B1 => n1425, B2 => 
                           n59804, ZN => n10222);
   U11857 : OAI22_X1 port map( A1 => n59807, A2 => n62115, B1 => n1424, B2 => 
                           n59804, ZN => n10223);
   U11858 : OAI22_X1 port map( A1 => n59807, A2 => n60968, B1 => n1423, B2 => 
                           n59804, ZN => n10224);
   U11859 : OAI22_X1 port map( A1 => n59807, A2 => n60982, B1 => n1422, B2 => 
                           n15269, ZN => n10225);
   U11860 : OAI22_X1 port map( A1 => n59807, A2 => n60996, B1 => n1421, B2 => 
                           n15269, ZN => n10226);
   U11861 : OAI22_X1 port map( A1 => n59807, A2 => n61010, B1 => n1420, B2 => 
                           n15269, ZN => n10227);
   U11862 : OAI22_X1 port map( A1 => n59808, A2 => n61024, B1 => n1419, B2 => 
                           n15269, ZN => n10228);
   U11863 : OAI22_X1 port map( A1 => n59808, A2 => n61038, B1 => n1418, B2 => 
                           n15269, ZN => n10229);
   U11864 : OAI22_X1 port map( A1 => n59808, A2 => n61052, B1 => n1417, B2 => 
                           n15269, ZN => n10230);
   U11865 : OAI22_X1 port map( A1 => n59808, A2 => n61066, B1 => n1416, B2 => 
                           n15269, ZN => n10231);
   U11866 : OAI22_X1 port map( A1 => n59808, A2 => n61080, B1 => n1415, B2 => 
                           n59804, ZN => n10232);
   U11867 : OAI22_X1 port map( A1 => n59809, A2 => n61094, B1 => n1414, B2 => 
                           n59804, ZN => n10233);
   U11868 : OAI22_X1 port map( A1 => n59809, A2 => n61108, B1 => n1413, B2 => 
                           n59804, ZN => n10234);
   U11869 : OAI22_X1 port map( A1 => n59809, A2 => n61122, B1 => n1412, B2 => 
                           n59804, ZN => n10235);
   U11870 : OAI22_X1 port map( A1 => n59809, A2 => n61136, B1 => n1411, B2 => 
                           n59804, ZN => n10236);
   U11871 : OAI22_X1 port map( A1 => n59760, A2 => n61976, B1 => n1314, B2 => 
                           n59759, ZN => n10053);
   U11872 : OAI22_X1 port map( A1 => n59760, A2 => n61990, B1 => n1313, B2 => 
                           n59759, ZN => n10054);
   U11873 : OAI22_X1 port map( A1 => n59760, A2 => n62004, B1 => n1312, B2 => 
                           n59759, ZN => n10055);
   U11874 : OAI22_X1 port map( A1 => n59760, A2 => n62018, B1 => n1311, B2 => 
                           n59759, ZN => n10056);
   U11875 : OAI22_X1 port map( A1 => n59760, A2 => n62032, B1 => n1310, B2 => 
                           n59759, ZN => n10057);
   U11876 : OAI22_X1 port map( A1 => n59761, A2 => n62046, B1 => n1309, B2 => 
                           n59759, ZN => n10058);
   U11877 : OAI22_X1 port map( A1 => n59761, A2 => n62060, B1 => n1308, B2 => 
                           n59759, ZN => n10059);
   U11878 : OAI22_X1 port map( A1 => n59761, A2 => n62074, B1 => n1307, B2 => 
                           n59759, ZN => n10060);
   U11879 : OAI22_X1 port map( A1 => n59761, A2 => n62088, B1 => n1306, B2 => 
                           n59759, ZN => n10061);
   U11880 : OAI22_X1 port map( A1 => n59761, A2 => n62102, B1 => n1305, B2 => 
                           n59759, ZN => n10062);
   U11881 : OAI22_X1 port map( A1 => n59762, A2 => n62116, B1 => n1304, B2 => 
                           n59759, ZN => n10063);
   U11882 : OAI22_X1 port map( A1 => n59762, A2 => n60969, B1 => n1303, B2 => 
                           n59759, ZN => n10064);
   U11883 : OAI22_X1 port map( A1 => n59762, A2 => n60983, B1 => n1302, B2 => 
                           n15285, ZN => n10065);
   U11884 : OAI22_X1 port map( A1 => n59762, A2 => n60997, B1 => n1301, B2 => 
                           n15285, ZN => n10066);
   U11885 : OAI22_X1 port map( A1 => n59762, A2 => n61011, B1 => n1300, B2 => 
                           n15285, ZN => n10067);
   U11886 : OAI22_X1 port map( A1 => n59763, A2 => n61025, B1 => n1299, B2 => 
                           n15285, ZN => n10068);
   U11887 : OAI22_X1 port map( A1 => n59763, A2 => n61039, B1 => n1298, B2 => 
                           n15285, ZN => n10069);
   U11888 : OAI22_X1 port map( A1 => n59763, A2 => n61053, B1 => n1297, B2 => 
                           n15285, ZN => n10070);
   U11889 : OAI22_X1 port map( A1 => n59763, A2 => n61067, B1 => n1296, B2 => 
                           n15285, ZN => n10071);
   U11890 : OAI22_X1 port map( A1 => n59763, A2 => n61081, B1 => n1295, B2 => 
                           n59759, ZN => n10072);
   U11891 : OAI22_X1 port map( A1 => n59764, A2 => n61095, B1 => n1294, B2 => 
                           n59759, ZN => n10073);
   U11892 : OAI22_X1 port map( A1 => n59764, A2 => n61109, B1 => n1293, B2 => 
                           n59759, ZN => n10074);
   U11893 : OAI22_X1 port map( A1 => n59764, A2 => n61123, B1 => n1292, B2 => 
                           n59759, ZN => n10075);
   U11894 : OAI22_X1 port map( A1 => n59764, A2 => n61137, B1 => n1291, B2 => 
                           n59759, ZN => n10076);
   U11895 : OAI22_X1 port map( A1 => n59752, A2 => n60983, B1 => n54451, B2 => 
                           n59748, ZN => n10033);
   U11896 : OAI22_X1 port map( A1 => n59752, A2 => n60997, B1 => n54450, B2 => 
                           n59748, ZN => n10034);
   U11897 : OAI22_X1 port map( A1 => n59752, A2 => n61011, B1 => n54449, B2 => 
                           n59748, ZN => n10035);
   U11898 : OAI22_X1 port map( A1 => n59752, A2 => n61025, B1 => n54448, B2 => 
                           n59748, ZN => n10036);
   U11899 : OAI22_X1 port map( A1 => n59753, A2 => n61039, B1 => n54447, B2 => 
                           n59748, ZN => n10037);
   U11900 : OAI22_X1 port map( A1 => n59753, A2 => n61053, B1 => n54446, B2 => 
                           n59748, ZN => n10038);
   U11901 : OAI22_X1 port map( A1 => n59753, A2 => n61067, B1 => n54445, B2 => 
                           n59748, ZN => n10039);
   U11902 : OAI22_X1 port map( A1 => n59751, A2 => n60969, B1 => n54444, B2 => 
                           n15286, ZN => n10032);
   U11903 : OAI22_X1 port map( A1 => n59753, A2 => n61081, B1 => n3934, B2 => 
                           n59748, ZN => n10040);
   U11904 : OAI22_X1 port map( A1 => n59754, A2 => n61095, B1 => n3933, B2 => 
                           n59748, ZN => n10041);
   U11905 : OAI22_X1 port map( A1 => n59754, A2 => n61109, B1 => n3932, B2 => 
                           n59748, ZN => n10042);
   U11906 : OAI22_X1 port map( A1 => n59754, A2 => n61123, B1 => n3931, B2 => 
                           n59748, ZN => n10043);
   U11907 : OAI22_X1 port map( A1 => n59754, A2 => n61137, B1 => n3930, B2 => 
                           n59748, ZN => n10044);
   U11908 : AND4_X1 port map( A1 => WR, A2 => EN, A3 => n5280, A4 => n5277, ZN 
                           => n15126);
   U11909 : AND4_X1 port map( A1 => ADDR_WR(4), A2 => WR, A3 => EN, A4 => n5277
                           , ZN => n15145);
   U11910 : OAI21_X1 port map( B1 => n9306, B2 => n61959, A => n7236, ZN => 
                           n9965);
   U11911 : OAI21_X1 port map( B1 => n7237, B2 => n7238, A => n61960, ZN => 
                           n7236);
   U11912 : NAND4_X1 port map( A1 => n7275, A2 => n7276, A3 => n7277, A4 => 
                           n7278, ZN => n7237);
   U11913 : NAND4_X1 port map( A1 => n7239, A2 => n7240, A3 => n7241, A4 => 
                           n7242, ZN => n7238);
   U11914 : OAI21_X1 port map( B1 => n9314, B2 => n61959, A => n7836, ZN => 
                           n9957);
   U11915 : OAI21_X1 port map( B1 => n7837, B2 => n7838, A => n61962, ZN => 
                           n7836);
   U11916 : NAND4_X1 port map( A1 => n7900, A2 => n7901, A3 => n7902, A4 => 
                           n7903, ZN => n7837);
   U11917 : NAND4_X1 port map( A1 => n7839, A2 => n7840, A3 => n7841, A4 => 
                           n7842, ZN => n7838);
   U11918 : OAI21_X1 port map( B1 => n9313, B2 => n61959, A => n7761, ZN => 
                           n9958);
   U11919 : OAI21_X1 port map( B1 => n7762, B2 => n7763, A => n61962, ZN => 
                           n7761);
   U11920 : NAND4_X1 port map( A1 => n7800, A2 => n7801, A3 => n7802, A4 => 
                           n7803, ZN => n7762);
   U11921 : NAND4_X1 port map( A1 => n7764, A2 => n7765, A3 => n7766, A4 => 
                           n7767, ZN => n7763);
   U11922 : OAI21_X1 port map( B1 => n9312, B2 => n61959, A => n7686, ZN => 
                           n9959);
   U11923 : OAI21_X1 port map( B1 => n7687, B2 => n7688, A => n61961, ZN => 
                           n7686);
   U11924 : NAND4_X1 port map( A1 => n7725, A2 => n7726, A3 => n7727, A4 => 
                           n7728, ZN => n7687);
   U11925 : NAND4_X1 port map( A1 => n7689, A2 => n7690, A3 => n7691, A4 => 
                           n7692, ZN => n7688);
   U11926 : OAI21_X1 port map( B1 => n9311, B2 => n61959, A => n7611, ZN => 
                           n9960);
   U11927 : OAI21_X1 port map( B1 => n7612, B2 => n7613, A => n61961, ZN => 
                           n7611);
   U11928 : NAND4_X1 port map( A1 => n7650, A2 => n7651, A3 => n7652, A4 => 
                           n7653, ZN => n7612);
   U11929 : NAND4_X1 port map( A1 => n7614, A2 => n7615, A3 => n7616, A4 => 
                           n7617, ZN => n7613);
   U11930 : OAI21_X1 port map( B1 => n9310, B2 => n61959, A => n7536, ZN => 
                           n9961);
   U11931 : OAI21_X1 port map( B1 => n7537, B2 => n7538, A => n61961, ZN => 
                           n7536);
   U11932 : NAND4_X1 port map( A1 => n7575, A2 => n7576, A3 => n7577, A4 => 
                           n7578, ZN => n7537);
   U11933 : NAND4_X1 port map( A1 => n7539, A2 => n7540, A3 => n7541, A4 => 
                           n7542, ZN => n7538);
   U11934 : OAI21_X1 port map( B1 => n9309, B2 => n61959, A => n7461, ZN => 
                           n9962);
   U11935 : OAI21_X1 port map( B1 => n7462, B2 => n7463, A => n61960, ZN => 
                           n7461);
   U11936 : NAND4_X1 port map( A1 => n7500, A2 => n7501, A3 => n7502, A4 => 
                           n7503, ZN => n7462);
   U11937 : NAND4_X1 port map( A1 => n7464, A2 => n7465, A3 => n7466, A4 => 
                           n7467, ZN => n7463);
   U11938 : OAI21_X1 port map( B1 => n9308, B2 => n61959, A => n7386, ZN => 
                           n9963);
   U11939 : OAI21_X1 port map( B1 => n7387, B2 => n7388, A => n61961, ZN => 
                           n7386);
   U11940 : NAND4_X1 port map( A1 => n7425, A2 => n7426, A3 => n7427, A4 => 
                           n7428, ZN => n7387);
   U11941 : NAND4_X1 port map( A1 => n7389, A2 => n7390, A3 => n7391, A4 => 
                           n7392, ZN => n7388);
   U11942 : OAI21_X1 port map( B1 => n9338, B2 => n61669, A => n14365, ZN => 
                           n9933);
   U11943 : OAI21_X1 port map( B1 => n14366, B2 => n14367, A => n61670, ZN => 
                           n14365);
   U11944 : NAND4_X1 port map( A1 => n14404, A2 => n14405, A3 => n14406, A4 => 
                           n14407, ZN => n14366);
   U11945 : NAND4_X1 port map( A1 => n14368, A2 => n14369, A3 => n14370, A4 => 
                           n14371, ZN => n14367);
   U11946 : OAI21_X1 port map( B1 => n9346, B2 => n61669, A => n14965, ZN => 
                           n9925);
   U11947 : OAI21_X1 port map( B1 => n14966, B2 => n14967, A => n61672, ZN => 
                           n14965);
   U11948 : NAND4_X1 port map( A1 => n15027, A2 => n15028, A3 => n15029, A4 => 
                           n15030, ZN => n14966);
   U11949 : NAND4_X1 port map( A1 => n14968, A2 => n14969, A3 => n14970, A4 => 
                           n14971, ZN => n14967);
   U11950 : OAI21_X1 port map( B1 => n9345, B2 => n61669, A => n14890, ZN => 
                           n9926);
   U11951 : OAI21_X1 port map( B1 => n14891, B2 => n14892, A => n61672, ZN => 
                           n14890);
   U11952 : NAND4_X1 port map( A1 => n14929, A2 => n14930, A3 => n14931, A4 => 
                           n14932, ZN => n14891);
   U11953 : NAND4_X1 port map( A1 => n14893, A2 => n14894, A3 => n14895, A4 => 
                           n14896, ZN => n14892);
   U11954 : OAI21_X1 port map( B1 => n9344, B2 => n61669, A => n14815, ZN => 
                           n9927);
   U11955 : OAI21_X1 port map( B1 => n14816, B2 => n14817, A => n61671, ZN => 
                           n14815);
   U11956 : NAND4_X1 port map( A1 => n14854, A2 => n14855, A3 => n14856, A4 => 
                           n14857, ZN => n14816);
   U11957 : NAND4_X1 port map( A1 => n14818, A2 => n14819, A3 => n14820, A4 => 
                           n14821, ZN => n14817);
   U11958 : OAI21_X1 port map( B1 => n9343, B2 => n61669, A => n14740, ZN => 
                           n9928);
   U11959 : OAI21_X1 port map( B1 => n14741, B2 => n14742, A => n61671, ZN => 
                           n14740);
   U11960 : NAND4_X1 port map( A1 => n14779, A2 => n14780, A3 => n14781, A4 => 
                           n14782, ZN => n14741);
   U11961 : NAND4_X1 port map( A1 => n14743, A2 => n14744, A3 => n14745, A4 => 
                           n14746, ZN => n14742);
   U11962 : OAI21_X1 port map( B1 => n9342, B2 => n61669, A => n14665, ZN => 
                           n9929);
   U11963 : OAI21_X1 port map( B1 => n14666, B2 => n14667, A => n61671, ZN => 
                           n14665);
   U11964 : NAND4_X1 port map( A1 => n14704, A2 => n14705, A3 => n14706, A4 => 
                           n14707, ZN => n14666);
   U11965 : NAND4_X1 port map( A1 => n14668, A2 => n14669, A3 => n14670, A4 => 
                           n14671, ZN => n14667);
   U11966 : OAI21_X1 port map( B1 => n9341, B2 => n61669, A => n14590, ZN => 
                           n9930);
   U11967 : OAI21_X1 port map( B1 => n14591, B2 => n14592, A => n61670, ZN => 
                           n14590);
   U11968 : NAND4_X1 port map( A1 => n14629, A2 => n14630, A3 => n14631, A4 => 
                           n14632, ZN => n14591);
   U11969 : NAND4_X1 port map( A1 => n14593, A2 => n14594, A3 => n14595, A4 => 
                           n14596, ZN => n14592);
   U11970 : OAI21_X1 port map( B1 => n9340, B2 => n61669, A => n14515, ZN => 
                           n9931);
   U11971 : OAI21_X1 port map( B1 => n14516, B2 => n14517, A => n61671, ZN => 
                           n14515);
   U11972 : NAND4_X1 port map( A1 => n14554, A2 => n14555, A3 => n14556, A4 => 
                           n14557, ZN => n14516);
   U11973 : NAND4_X1 port map( A1 => n14518, A2 => n14519, A3 => n14520, A4 => 
                           n14521, ZN => n14517);
   U11974 : OAI21_X1 port map( B1 => n9299, B2 => n61958, A => n6711, ZN => 
                           n9972);
   U11975 : OAI21_X1 port map( B1 => n6712, B2 => n6713, A => n61960, ZN => 
                           n6711);
   U11976 : NAND4_X1 port map( A1 => n6750, A2 => n6751, A3 => n6752, A4 => 
                           n6753, ZN => n6712);
   U11977 : NAND4_X1 port map( A1 => n6714, A2 => n6715, A3 => n6716, A4 => 
                           n6717, ZN => n6713);
   U11978 : OAI21_X1 port map( B1 => n9298, B2 => n61958, A => n6636, ZN => 
                           n9973);
   U11979 : OAI21_X1 port map( B1 => n6637, B2 => n6638, A => n61960, ZN => 
                           n6636);
   U11980 : NAND4_X1 port map( A1 => n6675, A2 => n6676, A3 => n6677, A4 => 
                           n6678, ZN => n6637);
   U11981 : NAND4_X1 port map( A1 => n6639, A2 => n6640, A3 => n6641, A4 => 
                           n6642, ZN => n6638);
   U11982 : OAI21_X1 port map( B1 => n9297, B2 => n61958, A => n6561, ZN => 
                           n9974);
   U11983 : OAI21_X1 port map( B1 => n6562, B2 => n6563, A => n61960, ZN => 
                           n6561);
   U11984 : NAND4_X1 port map( A1 => n6600, A2 => n6601, A3 => n6602, A4 => 
                           n6603, ZN => n6562);
   U11985 : NAND4_X1 port map( A1 => n6564, A2 => n6565, A3 => n6566, A4 => 
                           n6567, ZN => n6563);
   U11986 : OAI21_X1 port map( B1 => n9296, B2 => n61958, A => n6486, ZN => 
                           n9975);
   U11987 : OAI21_X1 port map( B1 => n6487, B2 => n6488, A => n61960, ZN => 
                           n6486);
   U11988 : NAND4_X1 port map( A1 => n6525, A2 => n6526, A3 => n6527, A4 => 
                           n6528, ZN => n6487);
   U11989 : NAND4_X1 port map( A1 => n6489, A2 => n6490, A3 => n6491, A4 => 
                           n6492, ZN => n6488);
   U11990 : OAI21_X1 port map( B1 => n9295, B2 => n61957, A => n6411, ZN => 
                           n9976);
   U11991 : OAI21_X1 port map( B1 => n6412, B2 => n6413, A => n61960, ZN => 
                           n6411);
   U11992 : NAND4_X1 port map( A1 => n6450, A2 => n6451, A3 => n6452, A4 => 
                           n6453, ZN => n6412);
   U11993 : NAND4_X1 port map( A1 => n6414, A2 => n6415, A3 => n6416, A4 => 
                           n6417, ZN => n6413);
   U11994 : OAI21_X1 port map( B1 => n9294, B2 => n61957, A => n6336, ZN => 
                           n9977);
   U11995 : OAI21_X1 port map( B1 => n6337, B2 => n6338, A => n61960, ZN => 
                           n6336);
   U11996 : NAND4_X1 port map( A1 => n6375, A2 => n6376, A3 => n6377, A4 => 
                           n6378, ZN => n6337);
   U11997 : NAND4_X1 port map( A1 => n6339, A2 => n6340, A3 => n6341, A4 => 
                           n6342, ZN => n6338);
   U11998 : OAI21_X1 port map( B1 => n9293, B2 => n61957, A => n6261, ZN => 
                           n9978);
   U11999 : OAI21_X1 port map( B1 => n6262, B2 => n6263, A => n61961, ZN => 
                           n6261);
   U12000 : NAND4_X1 port map( A1 => n6300, A2 => n6301, A3 => n6302, A4 => 
                           n6303, ZN => n6262);
   U12001 : NAND4_X1 port map( A1 => n6264, A2 => n6265, A3 => n6266, A4 => 
                           n6267, ZN => n6263);
   U12002 : OAI21_X1 port map( B1 => n9292, B2 => n61957, A => n6186, ZN => 
                           n9979);
   U12003 : OAI21_X1 port map( B1 => n6187, B2 => n6188, A => n61960, ZN => 
                           n6186);
   U12004 : NAND4_X1 port map( A1 => n6225, A2 => n6226, A3 => n6227, A4 => 
                           n6228, ZN => n6187);
   U12005 : NAND4_X1 port map( A1 => n6189, A2 => n6190, A3 => n6191, A4 => 
                           n6192, ZN => n6188);
   U12006 : OAI21_X1 port map( B1 => n9291, B2 => n61957, A => n6111, ZN => 
                           n9980);
   U12007 : OAI21_X1 port map( B1 => n6112, B2 => n6113, A => n61961, ZN => 
                           n6111);
   U12008 : NAND4_X1 port map( A1 => n6150, A2 => n6151, A3 => n6152, A4 => 
                           n6153, ZN => n6112);
   U12009 : NAND4_X1 port map( A1 => n6114, A2 => n6115, A3 => n6116, A4 => 
                           n6117, ZN => n6113);
   U12010 : OAI21_X1 port map( B1 => n9304, B2 => n61958, A => n7086, ZN => 
                           n9967);
   U12011 : OAI21_X1 port map( B1 => n7087, B2 => n7088, A => n61959, ZN => 
                           n7086);
   U12012 : NAND4_X1 port map( A1 => n7125, A2 => n7126, A3 => n7127, A4 => 
                           n7128, ZN => n7087);
   U12013 : NAND4_X1 port map( A1 => n7089, A2 => n7090, A3 => n7091, A4 => 
                           n7092, ZN => n7088);
   U12014 : OAI21_X1 port map( B1 => n9303, B2 => n61958, A => n7011, ZN => 
                           n9968);
   U12015 : OAI21_X1 port map( B1 => n7012, B2 => n7013, A => n61959, ZN => 
                           n7011);
   U12016 : NAND4_X1 port map( A1 => n7050, A2 => n7051, A3 => n7052, A4 => 
                           n7053, ZN => n7012);
   U12017 : NAND4_X1 port map( A1 => n7014, A2 => n7015, A3 => n7016, A4 => 
                           n7017, ZN => n7013);
   U12018 : OAI21_X1 port map( B1 => n9301, B2 => n61958, A => n6861, ZN => 
                           n9970);
   U12019 : OAI21_X1 port map( B1 => n6862, B2 => n6863, A => n61959, ZN => 
                           n6861);
   U12020 : NAND4_X1 port map( A1 => n6900, A2 => n6901, A3 => n6902, A4 => 
                           n6903, ZN => n6862);
   U12021 : NAND4_X1 port map( A1 => n6864, A2 => n6865, A3 => n6866, A4 => 
                           n6867, ZN => n6863);
   U12022 : OAI21_X1 port map( B1 => n9300, B2 => n61958, A => n6786, ZN => 
                           n9971);
   U12023 : OAI21_X1 port map( B1 => n6787, B2 => n6788, A => n61959, ZN => 
                           n6786);
   U12024 : NAND4_X1 port map( A1 => n6825, A2 => n6826, A3 => n6827, A4 => 
                           n6828, ZN => n6787);
   U12025 : NAND4_X1 port map( A1 => n6789, A2 => n6790, A3 => n6791, A4 => 
                           n6792, ZN => n6788);
   U12026 : OAI21_X1 port map( B1 => n9307, B2 => n61958, A => n7311, ZN => 
                           n9964);
   U12027 : OAI21_X1 port map( B1 => n7312, B2 => n7313, A => n61960, ZN => 
                           n7311);
   U12028 : NAND4_X1 port map( A1 => n7350, A2 => n7351, A3 => n7352, A4 => 
                           n7353, ZN => n7312);
   U12029 : NAND4_X1 port map( A1 => n7314, A2 => n7315, A3 => n7316, A4 => 
                           n7317, ZN => n7313);
   U12030 : OAI21_X1 port map( B1 => n9305, B2 => n61958, A => n7161, ZN => 
                           n9966);
   U12031 : OAI21_X1 port map( B1 => n7162, B2 => n7163, A => n61960, ZN => 
                           n7161);
   U12032 : NAND4_X1 port map( A1 => n7200, A2 => n7201, A3 => n7202, A4 => 
                           n7203, ZN => n7162);
   U12033 : NAND4_X1 port map( A1 => n7164, A2 => n7165, A3 => n7166, A4 => 
                           n7167, ZN => n7163);
   U12034 : OAI21_X1 port map( B1 => n9302, B2 => n61958, A => n6936, ZN => 
                           n9969);
   U12035 : OAI21_X1 port map( B1 => n6937, B2 => n6938, A => n61960, ZN => 
                           n6936);
   U12036 : NAND4_X1 port map( A1 => n6975, A2 => n6976, A3 => n6977, A4 => 
                           n6978, ZN => n6937);
   U12037 : NAND4_X1 port map( A1 => n6939, A2 => n6940, A3 => n6941, A4 => 
                           n6942, ZN => n6938);
   U12038 : OAI21_X1 port map( B1 => n9290, B2 => n61957, A => n6005, ZN => 
                           n9981);
   U12039 : OAI21_X1 port map( B1 => n6006, B2 => n6007, A => n61961, ZN => 
                           n6005);
   U12040 : NAND4_X1 port map( A1 => n6063, A2 => n6064, A3 => n6065, A4 => 
                           n6066, ZN => n6006);
   U12041 : NAND4_X1 port map( A1 => n6008, A2 => n6009, A3 => n6010, A4 => 
                           n6011, ZN => n6007);
   U12042 : OAI21_X1 port map( B1 => n9289, B2 => n61957, A => n5930, ZN => 
                           n9982);
   U12043 : OAI21_X1 port map( B1 => n5931, B2 => n5932, A => n61961, ZN => 
                           n5930);
   U12044 : NAND4_X1 port map( A1 => n5969, A2 => n5970, A3 => n5971, A4 => 
                           n5972, ZN => n5931);
   U12045 : NAND4_X1 port map( A1 => n5933, A2 => n5934, A3 => n5935, A4 => 
                           n5936, ZN => n5932);
   U12046 : OAI21_X1 port map( B1 => n9288, B2 => n61957, A => n5855, ZN => 
                           n9983);
   U12047 : OAI21_X1 port map( B1 => n5856, B2 => n5857, A => n61961, ZN => 
                           n5855);
   U12048 : NAND4_X1 port map( A1 => n5894, A2 => n5895, A3 => n5896, A4 => 
                           n5897, ZN => n5856);
   U12049 : NAND4_X1 port map( A1 => n5858, A2 => n5859, A3 => n5860, A4 => 
                           n5861, ZN => n5857);
   U12050 : OAI21_X1 port map( B1 => n9287, B2 => n61957, A => n5780, ZN => 
                           n9984);
   U12051 : OAI21_X1 port map( B1 => n5781, B2 => n5782, A => n61961, ZN => 
                           n5780);
   U12052 : NAND4_X1 port map( A1 => n5819, A2 => n5820, A3 => n5821, A4 => 
                           n5822, ZN => n5781);
   U12053 : NAND4_X1 port map( A1 => n5783, A2 => n5784, A3 => n5785, A4 => 
                           n5786, ZN => n5782);
   U12054 : OAI21_X1 port map( B1 => n9286, B2 => n61957, A => n5705, ZN => 
                           n9985);
   U12055 : OAI21_X1 port map( B1 => n5706, B2 => n5707, A => n61961, ZN => 
                           n5705);
   U12056 : NAND4_X1 port map( A1 => n5744, A2 => n5745, A3 => n5746, A4 => 
                           n5747, ZN => n5706);
   U12057 : NAND4_X1 port map( A1 => n5708, A2 => n5709, A3 => n5710, A4 => 
                           n5711, ZN => n5707);
   U12058 : OAI21_X1 port map( B1 => n9285, B2 => n61957, A => n5630, ZN => 
                           n9986);
   U12059 : OAI21_X1 port map( B1 => n5631, B2 => n5632, A => n61961, ZN => 
                           n5630);
   U12060 : NAND4_X1 port map( A1 => n5669, A2 => n5670, A3 => n5671, A4 => 
                           n5672, ZN => n5631);
   U12061 : NAND4_X1 port map( A1 => n5633, A2 => n5634, A3 => n5635, A4 => 
                           n5636, ZN => n5632);
   U12062 : OAI21_X1 port map( B1 => n9284, B2 => n61957, A => n5555, ZN => 
                           n9987);
   U12063 : OAI21_X1 port map( B1 => n5556, B2 => n5557, A => n61962, ZN => 
                           n5555);
   U12064 : NAND4_X1 port map( A1 => n5594, A2 => n5595, A3 => n5596, A4 => 
                           n5597, ZN => n5556);
   U12065 : NAND4_X1 port map( A1 => n5558, A2 => n5559, A3 => n5560, A4 => 
                           n5561, ZN => n5557);
   U12066 : OAI21_X1 port map( B1 => n9283, B2 => n61958, A => n5375, ZN => 
                           n9988);
   U12067 : OAI21_X1 port map( B1 => n5376, B2 => n5377, A => n61962, ZN => 
                           n5375);
   U12068 : NAND4_X1 port map( A1 => n5463, A2 => n5464, A3 => n5465, A4 => 
                           n5466, ZN => n5376);
   U12069 : NAND4_X1 port map( A1 => n5378, A2 => n5379, A3 => n5380, A4 => 
                           n5381, ZN => n5377);
   U12070 : OAI21_X1 port map( B1 => n9337, B2 => n61668, A => n9874, ZN => 
                           n9934);
   U12071 : OAI21_X1 port map( B1 => n9875, B2 => n9876, A => n61670, ZN => 
                           n9874);
   U12072 : NAND4_X1 port map( A1 => n9913, A2 => n9914, A3 => n9915, A4 => 
                           n9916, ZN => n9875);
   U12073 : NAND4_X1 port map( A1 => n9877, A2 => n9878, A3 => n9879, A4 => 
                           n9880, ZN => n9876);
   U12074 : OAI21_X1 port map( B1 => n9336, B2 => n61668, A => n9735, ZN => 
                           n9935);
   U12075 : OAI21_X1 port map( B1 => n9736, B2 => n9737, A => n61669, ZN => 
                           n9735);
   U12076 : NAND4_X1 port map( A1 => n9838, A2 => n9839, A3 => n9840, A4 => 
                           n9841, ZN => n9736);
   U12077 : NAND4_X1 port map( A1 => n9738, A2 => n9739, A3 => n9740, A4 => 
                           n9741, ZN => n9737);
   U12078 : OAI21_X1 port map( B1 => n9335, B2 => n61668, A => n9660, ZN => 
                           n9936);
   U12079 : OAI21_X1 port map( B1 => n9661, B2 => n9662, A => n61669, ZN => 
                           n9660);
   U12080 : NAND4_X1 port map( A1 => n9699, A2 => n9700, A3 => n9701, A4 => 
                           n9702, ZN => n9661);
   U12081 : NAND4_X1 port map( A1 => n9663, A2 => n9664, A3 => n9665, A4 => 
                           n9666, ZN => n9662);
   U12082 : OAI21_X1 port map( B1 => n9334, B2 => n61668, A => n9569, ZN => 
                           n9937);
   U12083 : OAI21_X1 port map( B1 => n9570, B2 => n9571, A => n61670, ZN => 
                           n9569);
   U12084 : NAND4_X1 port map( A1 => n9624, A2 => n9625, A3 => n9626, A4 => 
                           n9627, ZN => n9570);
   U12085 : NAND4_X1 port map( A1 => n9572, A2 => n9573, A3 => n9574, A4 => 
                           n9575, ZN => n9571);
   U12086 : OAI21_X1 port map( B1 => n9333, B2 => n61668, A => n9494, ZN => 
                           n9938);
   U12087 : OAI21_X1 port map( B1 => n9495, B2 => n9496, A => n61669, ZN => 
                           n9494);
   U12088 : NAND4_X1 port map( A1 => n9533, A2 => n9534, A3 => n9535, A4 => 
                           n9536, ZN => n9495);
   U12089 : NAND4_X1 port map( A1 => n9497, A2 => n9498, A3 => n9499, A4 => 
                           n9500, ZN => n9496);
   U12090 : OAI21_X1 port map( B1 => n9332, B2 => n61668, A => n9419, ZN => 
                           n9939);
   U12091 : OAI21_X1 port map( B1 => n9420, B2 => n9421, A => n61669, ZN => 
                           n9419);
   U12092 : NAND4_X1 port map( A1 => n9458, A2 => n9459, A3 => n9460, A4 => 
                           n9461, ZN => n9420);
   U12093 : NAND4_X1 port map( A1 => n9422, A2 => n9423, A3 => n9424, A4 => 
                           n9425, ZN => n9421);
   U12094 : OAI21_X1 port map( B1 => n9331, B2 => n61668, A => n9280, ZN => 
                           n9940);
   U12095 : OAI21_X1 port map( B1 => n9281, B2 => n9282, A => n61670, ZN => 
                           n9280);
   U12096 : NAND4_X1 port map( A1 => n9383, A2 => n9384, A3 => n9385, A4 => 
                           n9386, ZN => n9281);
   U12097 : NAND4_X1 port map( A1 => n9347, A2 => n9348, A3 => n9349, A4 => 
                           n9350, ZN => n9282);
   U12098 : OAI21_X1 port map( B1 => n9330, B2 => n61668, A => n9205, ZN => 
                           n9941);
   U12099 : OAI21_X1 port map( B1 => n9206, B2 => n9207, A => n61670, ZN => 
                           n9205);
   U12100 : NAND4_X1 port map( A1 => n9244, A2 => n9245, A3 => n9246, A4 => 
                           n9247, ZN => n9206);
   U12101 : NAND4_X1 port map( A1 => n9208, A2 => n9209, A3 => n9210, A4 => 
                           n9211, ZN => n9207);
   U12102 : OAI21_X1 port map( B1 => n9329, B2 => n61668, A => n9130, ZN => 
                           n9942);
   U12103 : OAI21_X1 port map( B1 => n9131, B2 => n9132, A => n61670, ZN => 
                           n9130);
   U12104 : NAND4_X1 port map( A1 => n9169, A2 => n9170, A3 => n9171, A4 => 
                           n9172, ZN => n9131);
   U12105 : NAND4_X1 port map( A1 => n9133, A2 => n9134, A3 => n9135, A4 => 
                           n9136, ZN => n9132);
   U12106 : OAI21_X1 port map( B1 => n9328, B2 => n61668, A => n9055, ZN => 
                           n9943);
   U12107 : OAI21_X1 port map( B1 => n9056, B2 => n9057, A => n61670, ZN => 
                           n9055);
   U12108 : NAND4_X1 port map( A1 => n9094, A2 => n9095, A3 => n9096, A4 => 
                           n9097, ZN => n9056);
   U12109 : NAND4_X1 port map( A1 => n9058, A2 => n9059, A3 => n9060, A4 => 
                           n9061, ZN => n9057);
   U12110 : OAI21_X1 port map( B1 => n9327, B2 => n61667, A => n8980, ZN => 
                           n9944);
   U12111 : OAI21_X1 port map( B1 => n8981, B2 => n8982, A => n61670, ZN => 
                           n8980);
   U12112 : NAND4_X1 port map( A1 => n9019, A2 => n9020, A3 => n9021, A4 => 
                           n9022, ZN => n8981);
   U12113 : NAND4_X1 port map( A1 => n8983, A2 => n8984, A3 => n8985, A4 => 
                           n8986, ZN => n8982);
   U12114 : OAI21_X1 port map( B1 => n9326, B2 => n61667, A => n8905, ZN => 
                           n9945);
   U12115 : OAI21_X1 port map( B1 => n8906, B2 => n8907, A => n61670, ZN => 
                           n8905);
   U12116 : NAND4_X1 port map( A1 => n8944, A2 => n8945, A3 => n8946, A4 => 
                           n8947, ZN => n8906);
   U12117 : NAND4_X1 port map( A1 => n8908, A2 => n8909, A3 => n8910, A4 => 
                           n8911, ZN => n8907);
   U12118 : OAI21_X1 port map( B1 => n9325, B2 => n61667, A => n8830, ZN => 
                           n9946);
   U12119 : OAI21_X1 port map( B1 => n8831, B2 => n8832, A => n61671, ZN => 
                           n8830);
   U12120 : NAND4_X1 port map( A1 => n8869, A2 => n8870, A3 => n8871, A4 => 
                           n8872, ZN => n8831);
   U12121 : NAND4_X1 port map( A1 => n8833, A2 => n8834, A3 => n8835, A4 => 
                           n8836, ZN => n8832);
   U12122 : OAI21_X1 port map( B1 => n9324, B2 => n61667, A => n8755, ZN => 
                           n9947);
   U12123 : OAI21_X1 port map( B1 => n8756, B2 => n8757, A => n61670, ZN => 
                           n8755);
   U12124 : NAND4_X1 port map( A1 => n8794, A2 => n8795, A3 => n8796, A4 => 
                           n8797, ZN => n8756);
   U12125 : NAND4_X1 port map( A1 => n8758, A2 => n8759, A3 => n8760, A4 => 
                           n8761, ZN => n8757);
   U12126 : OAI21_X1 port map( B1 => n9323, B2 => n61667, A => n8680, ZN => 
                           n9948);
   U12127 : OAI21_X1 port map( B1 => n8681, B2 => n8682, A => n61671, ZN => 
                           n8680);
   U12128 : NAND4_X1 port map( A1 => n8719, A2 => n8720, A3 => n8721, A4 => 
                           n8722, ZN => n8681);
   U12129 : NAND4_X1 port map( A1 => n8683, A2 => n8684, A3 => n8685, A4 => 
                           n8686, ZN => n8682);
   U12130 : OAI21_X1 port map( B1 => n9322, B2 => n61667, A => n8605, ZN => 
                           n9949);
   U12131 : OAI21_X1 port map( B1 => n8606, B2 => n8607, A => n61671, ZN => 
                           n8605);
   U12132 : NAND4_X1 port map( A1 => n8644, A2 => n8645, A3 => n8646, A4 => 
                           n8647, ZN => n8606);
   U12133 : NAND4_X1 port map( A1 => n8608, A2 => n8609, A3 => n8610, A4 => 
                           n8611, ZN => n8607);
   U12134 : OAI21_X1 port map( B1 => n9321, B2 => n61667, A => n8530, ZN => 
                           n9950);
   U12135 : OAI21_X1 port map( B1 => n8531, B2 => n8532, A => n61671, ZN => 
                           n8530);
   U12136 : NAND4_X1 port map( A1 => n8569, A2 => n8570, A3 => n8571, A4 => 
                           n8572, ZN => n8531);
   U12137 : NAND4_X1 port map( A1 => n8533, A2 => n8534, A3 => n8535, A4 => 
                           n8536, ZN => n8532);
   U12138 : OAI21_X1 port map( B1 => n9320, B2 => n61667, A => n8455, ZN => 
                           n9951);
   U12139 : OAI21_X1 port map( B1 => n8456, B2 => n8457, A => n61671, ZN => 
                           n8455);
   U12140 : NAND4_X1 port map( A1 => n8494, A2 => n8495, A3 => n8496, A4 => 
                           n8497, ZN => n8456);
   U12141 : NAND4_X1 port map( A1 => n8458, A2 => n8459, A3 => n8460, A4 => 
                           n8461, ZN => n8457);
   U12142 : OAI21_X1 port map( B1 => n9319, B2 => n61667, A => n8380, ZN => 
                           n9952);
   U12143 : OAI21_X1 port map( B1 => n8381, B2 => n8382, A => n61671, ZN => 
                           n8380);
   U12144 : NAND4_X1 port map( A1 => n8419, A2 => n8420, A3 => n8421, A4 => 
                           n8422, ZN => n8381);
   U12145 : NAND4_X1 port map( A1 => n8383, A2 => n8384, A3 => n8385, A4 => 
                           n8386, ZN => n8382);
   U12146 : OAI21_X1 port map( B1 => n9318, B2 => n61667, A => n8305, ZN => 
                           n9953);
   U12147 : OAI21_X1 port map( B1 => n8306, B2 => n8307, A => n61671, ZN => 
                           n8305);
   U12148 : NAND4_X1 port map( A1 => n8344, A2 => n8345, A3 => n8346, A4 => 
                           n8347, ZN => n8306);
   U12149 : NAND4_X1 port map( A1 => n8308, A2 => n8309, A3 => n8310, A4 => 
                           n8311, ZN => n8307);
   U12150 : OAI21_X1 port map( B1 => n9317, B2 => n61667, A => n8230, ZN => 
                           n9954);
   U12151 : OAI21_X1 port map( B1 => n8231, B2 => n8232, A => n61671, ZN => 
                           n8230);
   U12152 : NAND4_X1 port map( A1 => n8269, A2 => n8270, A3 => n8271, A4 => 
                           n8272, ZN => n8231);
   U12153 : NAND4_X1 port map( A1 => n8233, A2 => n8234, A3 => n8235, A4 => 
                           n8236, ZN => n8232);
   U12154 : OAI21_X1 port map( B1 => n9316, B2 => n61667, A => n8155, ZN => 
                           n9955);
   U12155 : OAI21_X1 port map( B1 => n8156, B2 => n8157, A => n61672, ZN => 
                           n8155);
   U12156 : NAND4_X1 port map( A1 => n8194, A2 => n8195, A3 => n8196, A4 => 
                           n8197, ZN => n8156);
   U12157 : NAND4_X1 port map( A1 => n8158, A2 => n8159, A3 => n8160, A4 => 
                           n8161, ZN => n8157);
   U12158 : OAI21_X1 port map( B1 => n9315, B2 => n61668, A => n7944, ZN => 
                           n9956);
   U12159 : OAI21_X1 port map( B1 => n7945, B2 => n7946, A => n61672, ZN => 
                           n7944);
   U12160 : NAND4_X1 port map( A1 => n8051, A2 => n8052, A3 => n8053, A4 => 
                           n8054, ZN => n7945);
   U12161 : NAND4_X1 port map( A1 => n7947, A2 => n7948, A3 => n7949, A4 => 
                           n7950, ZN => n7946);
   U12162 : OAI21_X1 port map( B1 => n9339, B2 => n61668, A => n14440, ZN => 
                           n9932);
   U12163 : OAI21_X1 port map( B1 => n14441, B2 => n14442, A => n61670, ZN => 
                           n14440);
   U12164 : NAND4_X1 port map( A1 => n14479, A2 => n14480, A3 => n14481, A4 => 
                           n14482, ZN => n14441);
   U12165 : NAND4_X1 port map( A1 => n14443, A2 => n14444, A3 => n14445, A4 => 
                           n14446, ZN => n14442);
   U12166 : INV_X1 port map( A => n7108, ZN => n1525);
   U12167 : OAI222_X1 port map( A1 => n1526, A2 => n59737, B1 => n59740, B2 => 
                           n1578, C1 => n1590, C2 => n59744, ZN => n7108);
   U12168 : INV_X1 port map( A => n7033, ZN => n1523);
   U12169 : OAI222_X1 port map( A1 => n1524, A2 => n59737, B1 => n59741, B2 => 
                           n1577, C1 => n1589, C2 => n59745, ZN => n7033);
   U12170 : INV_X1 port map( A => n6883, ZN => n1519);
   U12171 : OAI222_X1 port map( A1 => n1520, A2 => n59738, B1 => n59743, B2 => 
                           n1575, C1 => n1557, C2 => n59747, ZN => n6883);
   U12172 : INV_X1 port map( A => n7258, ZN => n1529);
   U12173 : OAI222_X1 port map( A1 => n1530, A2 => n59738, B1 => n59740, B2 => 
                           n1580, C1 => n1608, C2 => n59744, ZN => n7258);
   U12174 : INV_X1 port map( A => n7876, ZN => n1545);
   U12175 : OAI222_X1 port map( A1 => n1546, A2 => n59739, B1 => n59740, B2 => 
                           n1588, C1 => n1616, C2 => n59744, ZN => n7876);
   U12176 : INV_X1 port map( A => n7783, ZN => n1543);
   U12177 : OAI222_X1 port map( A1 => n1544, A2 => n59737, B1 => n59741, B2 => 
                           n1587, C1 => n1615, C2 => n59745, ZN => n7783);
   U12178 : INV_X1 port map( A => n7708, ZN => n1541);
   U12179 : OAI222_X1 port map( A1 => n1542, A2 => n59737, B1 => n59740, B2 => 
                           n1586, C1 => n1614, C2 => n59744, ZN => n7708);
   U12180 : INV_X1 port map( A => n7633, ZN => n1539);
   U12181 : OAI222_X1 port map( A1 => n1540, A2 => n59738, B1 => n59741, B2 => 
                           n1585, C1 => n1613, C2 => n59745, ZN => n7633);
   U12182 : INV_X1 port map( A => n7558, ZN => n1537);
   U12183 : OAI222_X1 port map( A1 => n1538, A2 => n59738, B1 => n59742, B2 => 
                           n1584, C1 => n1612, C2 => n59746, ZN => n7558);
   U12184 : INV_X1 port map( A => n7483, ZN => n1535);
   U12185 : OAI222_X1 port map( A1 => n1536, A2 => n59739, B1 => n59743, B2 => 
                           n1583, C1 => n1611, C2 => n59747, ZN => n7483);
   U12186 : INV_X1 port map( A => n7408, ZN => n1533);
   U12187 : OAI222_X1 port map( A1 => n1534, A2 => n59737, B1 => n59742, B2 => 
                           n1582, C1 => n1610, C2 => n59746, ZN => n7408);
   U12188 : INV_X1 port map( A => n7333, ZN => n1531);
   U12189 : OAI222_X1 port map( A1 => n1532, A2 => n59739, B1 => n59743, B2 => 
                           n1581, C1 => n1609, C2 => n59747, ZN => n7333);
   U12190 : INV_X1 port map( A => n7183, ZN => n1527);
   U12191 : OAI222_X1 port map( A1 => n1528, A2 => n59739, B1 => n59741, B2 => 
                           n1579, C1 => n1607, C2 => n59745, ZN => n7183);
   U12192 : INV_X1 port map( A => n6958, ZN => n1521);
   U12193 : OAI222_X1 port map( A1 => n1522, A2 => n59738, B1 => n59742, B2 => 
                           n1576, C1 => n1558, C2 => n59746, ZN => n6958);
   U12194 : NAND2_X1 port map( A1 => DATA_IN(3), A2 => n62186, ZN => n5370);
   U12195 : AND3_X1 port map( A1 => EN, A2 => n62198, A3 => RD1, ZN => n5374);
   U12196 : NAND2_X1 port map( A1 => DATA_IN(0), A2 => n62186, ZN => n5373);
   U12197 : NAND2_X1 port map( A1 => DATA_IN(1), A2 => n62186, ZN => n5372);
   U12198 : NAND2_X1 port map( A1 => DATA_IN(19), A2 => n62185, ZN => n15085);
   U12199 : NAND2_X1 port map( A1 => DATA_IN(20), A2 => n62185, ZN => n15084);
   U12200 : NAND2_X1 port map( A1 => DATA_IN(21), A2 => n62185, ZN => n15083);
   U12201 : NAND2_X1 port map( A1 => DATA_IN(22), A2 => n62186, ZN => n15082);
   U12202 : NAND2_X1 port map( A1 => DATA_IN(23), A2 => n62185, ZN => n15081);
   U12203 : NAND2_X1 port map( A1 => DATA_IN(11), A2 => n62185, ZN => n15093);
   U12204 : NAND2_X1 port map( A1 => DATA_IN(12), A2 => n62185, ZN => n15092);
   U12205 : NAND2_X1 port map( A1 => DATA_IN(13), A2 => n62185, ZN => n15091);
   U12206 : NAND2_X1 port map( A1 => DATA_IN(14), A2 => n62185, ZN => n15090);
   U12207 : NAND2_X1 port map( A1 => DATA_IN(15), A2 => n62185, ZN => n15089);
   U12208 : NAND2_X1 port map( A1 => DATA_IN(16), A2 => n62185, ZN => n15088);
   U12209 : NAND2_X1 port map( A1 => DATA_IN(17), A2 => n62185, ZN => n15087);
   U12210 : NAND2_X1 port map( A1 => DATA_IN(18), A2 => n62185, ZN => n15086);
   U12211 : NAND2_X1 port map( A1 => DATA_IN(4), A2 => n62187, ZN => n5369);
   U12212 : NAND2_X1 port map( A1 => DATA_IN(5), A2 => n62187, ZN => n5368);
   U12213 : NAND2_X1 port map( A1 => DATA_IN(6), A2 => n62187, ZN => n5367);
   U12214 : NAND2_X1 port map( A1 => DATA_IN(7), A2 => n62187, ZN => n5366);
   U12215 : NAND2_X1 port map( A1 => DATA_IN(8), A2 => n62187, ZN => n5365);
   U12216 : NAND2_X1 port map( A1 => DATA_IN(9), A2 => n62187, ZN => n5364);
   U12217 : NAND2_X1 port map( A1 => DATA_IN(10), A2 => n62187, ZN => n5363);
   U12218 : NAND2_X1 port map( A1 => DATA_IN(24), A2 => n62186, ZN => n15080);
   U12219 : NAND2_X1 port map( A1 => DATA_IN(25), A2 => n62186, ZN => n15079);
   U12220 : NAND2_X1 port map( A1 => DATA_IN(26), A2 => n62186, ZN => n15078);
   U12221 : NAND2_X1 port map( A1 => DATA_IN(27), A2 => n62186, ZN => n15077);
   U12222 : NAND2_X1 port map( A1 => DATA_IN(28), A2 => n62186, ZN => n15076);
   U12223 : NAND2_X1 port map( A1 => DATA_IN(29), A2 => n62186, ZN => n15075);
   U12224 : NAND2_X1 port map( A1 => DATA_IN(30), A2 => n62186, ZN => n15074);
   U12225 : NAND2_X1 port map( A1 => DATA_IN(31), A2 => n62186, ZN => n15072);
   U12226 : NAND2_X1 port map( A1 => DATA_IN(2), A2 => n62187, ZN => n5371);
   U12227 : AND3_X1 port map( A1 => EN, A2 => n62198, A3 => RD2, ZN => n7943);
   U12228 : INV_X1 port map( A => RST, ZN => n5276);
   U12229 : NOR3_X4 port map( A1 => ADDR_RD2(0), A2 => ADDR_RD2(1), A3 => n5359
                           , ZN => n14985);
   U12230 : NOR3_X4 port map( A1 => n5361, A2 => ADDR_RD2(1), A3 => n5359, ZN 
                           => n14986);
   U12231 : NOR3_X4 port map( A1 => ADDR_RD2(1), A2 => ADDR_RD2(2), A3 => n5361
                           , ZN => n14981);
   U12232 : NOR3_X4 port map( A1 => ADDR_RD2(1), A2 => ADDR_RD2(2), A3 => 
                           ADDR_RD2(0), ZN => n14980);
   U12233 : NOR3_X4 port map( A1 => n5353, A2 => ADDR_RD1(2), A3 => n5352, ZN 
                           => n7859);
   U12234 : NOR3_X4 port map( A1 => ADDR_RD1(0), A2 => ADDR_RD1(1), A3 => n5351
                           , ZN => n7852);
   U12235 : NOR3_X4 port map( A1 => n5352, A2 => ADDR_RD1(0), A3 => n5351, ZN 
                           => n7850);
   U12236 : NOR3_X4 port map( A1 => n5353, A2 => ADDR_RD1(1), A3 => n5351, ZN 
                           => n7864);
   U12237 : NOR3_X4 port map( A1 => ADDR_RD1(1), A2 => ADDR_RD1(2), A3 => n5353
                           , ZN => n7862);
   U12238 : NOR3_X4 port map( A1 => ADDR_RD1(0), A2 => ADDR_RD1(2), A3 => n5352
                           , ZN => n7860);
   U12239 : NOR3_X4 port map( A1 => ADDR_RD1(1), A2 => ADDR_RD1(2), A3 => 
                           ADDR_RD1(0), ZN => n7856);
   U12240 : CLKBUF_X1 port map( A => n60957, Z => n60969);
   U12241 : CLKBUF_X1 port map( A => n60971, Z => n60983);
   U12242 : CLKBUF_X1 port map( A => n60985, Z => n60997);
   U12243 : CLKBUF_X1 port map( A => n60999, Z => n61011);
   U12244 : CLKBUF_X1 port map( A => n61013, Z => n61025);
   U12245 : CLKBUF_X1 port map( A => n61027, Z => n61039);
   U12246 : CLKBUF_X1 port map( A => n61041, Z => n61053);
   U12247 : CLKBUF_X1 port map( A => n61055, Z => n61067);
   U12248 : CLKBUF_X1 port map( A => n61069, Z => n61081);
   U12249 : CLKBUF_X1 port map( A => n61083, Z => n61095);
   U12250 : CLKBUF_X1 port map( A => n61097, Z => n61109);
   U12251 : CLKBUF_X1 port map( A => n61111, Z => n61123);
   U12252 : CLKBUF_X1 port map( A => n61125, Z => n61137);
   U12253 : CLKBUF_X1 port map( A => n61139, Z => n61151);
   U12254 : CLKBUF_X1 port map( A => n61153, Z => n61165);
   U12255 : CLKBUF_X1 port map( A => n61167, Z => n61179);
   U12256 : CLKBUF_X1 port map( A => n61181, Z => n61193);
   U12257 : CLKBUF_X1 port map( A => n61195, Z => n61207);
   U12258 : CLKBUF_X1 port map( A => n61209, Z => n61221);
   U12259 : CLKBUF_X1 port map( A => n61223, Z => n61235);
   U12260 : CLKBUF_X1 port map( A => n61246, Z => n61258);
   U12261 : CLKBUF_X1 port map( A => n7943, Z => n61672);
   U12262 : INV_X1 port map( A => n6107, ZN => n61674);
   U12263 : INV_X1 port map( A => n6092, ZN => n61678);
   U12264 : INV_X1 port map( A => n6089, ZN => n61682);
   U12265 : INV_X1 port map( A => n6086, ZN => n61686);
   U12266 : INV_X1 port map( A => n6078, ZN => n61690);
   U12267 : INV_X1 port map( A => n6073, ZN => n61694);
   U12268 : INV_X1 port map( A => n6062, ZN => n61698);
   U12269 : INV_X1 port map( A => n6059, ZN => n61702);
   U12270 : INV_X1 port map( A => n6056, ZN => n61706);
   U12271 : INV_X1 port map( A => n6048, ZN => n61710);
   U12272 : INV_X1 port map( A => n6047, ZN => n61712);
   U12273 : INV_X1 port map( A => n6044, ZN => n61714);
   U12274 : INV_X1 port map( A => n6034, ZN => n61720);
   U12275 : INV_X1 port map( A => n6033, ZN => n61722);
   U12276 : INV_X1 port map( A => n6025, ZN => n61724);
   U12277 : INV_X1 port map( A => n6021, ZN => n61728);
   U12278 : INV_X1 port map( A => n6018, ZN => n61732);
   U12279 : CLKBUF_X1 port map( A => n5374, Z => n61962);
   U12280 : CLKBUF_X1 port map( A => n61964, Z => n61976);
   U12281 : CLKBUF_X1 port map( A => n61978, Z => n61990);
   U12282 : CLKBUF_X1 port map( A => n61992, Z => n62004);
   U12283 : CLKBUF_X1 port map( A => n62006, Z => n62018);
   U12284 : CLKBUF_X1 port map( A => n62020, Z => n62032);
   U12285 : CLKBUF_X1 port map( A => n62034, Z => n62046);
   U12286 : CLKBUF_X1 port map( A => n62048, Z => n62060);
   U12287 : CLKBUF_X1 port map( A => n62062, Z => n62074);
   U12288 : CLKBUF_X1 port map( A => n62076, Z => n62088);
   U12289 : CLKBUF_X1 port map( A => n62090, Z => n62102);
   U12290 : CLKBUF_X1 port map( A => n62104, Z => n62116);
   U12291 : CLKBUF_X1 port map( A => n62184, Z => n62198);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_generic_M8_N8_F8_DATA_BIT32.all;

entity MUX21_GENERIC_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32;

architecture SYN_BEH of MUX21_GENERIC_NBIT32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n180, ZN => n170);
   U2 : INV_X1 port map( A => n180, ZN => n171);
   U3 : BUF_X1 port map( A => n169, Z => n178);
   U4 : BUF_X1 port map( A => n168, Z => n177);
   U5 : BUF_X1 port map( A => n168, Z => n176);
   U6 : BUF_X1 port map( A => n168, Z => n175);
   U7 : BUF_X1 port map( A => n167, Z => n174);
   U8 : BUF_X1 port map( A => n167, Z => n173);
   U9 : BUF_X1 port map( A => n167, Z => n172);
   U10 : BUF_X1 port map( A => n169, Z => n180);
   U11 : BUF_X1 port map( A => n169, Z => n179);
   U12 : INV_X1 port map( A => n62, ZN => Y(3));
   U13 : AOI22_X1 port map( A1 => A(3), A2 => n170, B1 => B(3), B2 => n178, ZN 
                           => n62);
   U14 : INV_X1 port map( A => n65, ZN => Y(0));
   U15 : AOI22_X1 port map( A1 => A(0), A2 => n170, B1 => B(0), B2 => n179, ZN 
                           => n65);
   U16 : INV_X1 port map( A => n64, ZN => Y(1));
   U17 : AOI22_X1 port map( A1 => A(1), A2 => n170, B1 => B(1), B2 => n179, ZN 
                           => n64);
   U18 : INV_X1 port map( A => n46, ZN => Y(19));
   U19 : AOI22_X1 port map( A1 => A(19), A2 => n171, B1 => B(19), B2 => n174, 
                           ZN => n46);
   U20 : INV_X1 port map( A => n45, ZN => Y(20));
   U21 : AOI22_X1 port map( A1 => A(20), A2 => n171, B1 => B(20), B2 => n174, 
                           ZN => n45);
   U22 : INV_X1 port map( A => n44, ZN => Y(21));
   U23 : AOI22_X1 port map( A1 => A(21), A2 => n171, B1 => B(21), B2 => n174, 
                           ZN => n44);
   U24 : INV_X1 port map( A => n43, ZN => Y(22));
   U25 : AOI22_X1 port map( A1 => A(22), A2 => n171, B1 => B(22), B2 => n173, 
                           ZN => n43);
   U26 : INV_X1 port map( A => n42, ZN => Y(23));
   U27 : AOI22_X1 port map( A1 => A(23), A2 => n171, B1 => B(23), B2 => n176, 
                           ZN => n42);
   U28 : INV_X1 port map( A => n54, ZN => Y(11));
   U29 : AOI22_X1 port map( A1 => A(11), A2 => n170, B1 => B(11), B2 => n176, 
                           ZN => n54);
   U30 : INV_X1 port map( A => n53, ZN => Y(12));
   U31 : AOI22_X1 port map( A1 => A(12), A2 => n171, B1 => B(12), B2 => n176, 
                           ZN => n53);
   U32 : INV_X1 port map( A => n52, ZN => Y(13));
   U33 : AOI22_X1 port map( A1 => A(13), A2 => n171, B1 => B(13), B2 => n176, 
                           ZN => n52);
   U34 : INV_X1 port map( A => n51, ZN => Y(14));
   U35 : AOI22_X1 port map( A1 => A(14), A2 => n171, B1 => B(14), B2 => n175, 
                           ZN => n51);
   U36 : INV_X1 port map( A => n50, ZN => Y(15));
   U37 : AOI22_X1 port map( A1 => A(15), A2 => n171, B1 => B(15), B2 => n175, 
                           ZN => n50);
   U38 : INV_X1 port map( A => n49, ZN => Y(16));
   U39 : AOI22_X1 port map( A1 => A(16), A2 => n171, B1 => B(16), B2 => n175, 
                           ZN => n49);
   U40 : INV_X1 port map( A => n48, ZN => Y(17));
   U41 : AOI22_X1 port map( A1 => A(17), A2 => n171, B1 => B(17), B2 => n175, 
                           ZN => n48);
   U42 : INV_X1 port map( A => n47, ZN => Y(18));
   U43 : AOI22_X1 port map( A1 => A(18), A2 => n171, B1 => B(18), B2 => n174, 
                           ZN => n47);
   U44 : INV_X1 port map( A => n61, ZN => Y(4));
   U45 : AOI22_X1 port map( A1 => A(4), A2 => n170, B1 => B(4), B2 => n178, ZN 
                           => n61);
   U46 : INV_X1 port map( A => n60, ZN => Y(5));
   U47 : AOI22_X1 port map( A1 => A(5), A2 => n170, B1 => B(5), B2 => n178, ZN 
                           => n60);
   U48 : INV_X1 port map( A => n59, ZN => Y(6));
   U49 : AOI22_X1 port map( A1 => A(6), A2 => n170, B1 => B(6), B2 => n178, ZN 
                           => n59);
   U50 : INV_X1 port map( A => n58, ZN => Y(7));
   U51 : AOI22_X1 port map( A1 => A(7), A2 => n170, B1 => B(7), B2 => n177, ZN 
                           => n58);
   U52 : INV_X1 port map( A => n57, ZN => Y(8));
   U53 : AOI22_X1 port map( A1 => A(8), A2 => n170, B1 => B(8), B2 => n177, ZN 
                           => n57);
   U54 : INV_X1 port map( A => n56, ZN => Y(9));
   U55 : AOI22_X1 port map( A1 => A(9), A2 => n170, B1 => B(9), B2 => n177, ZN 
                           => n56);
   U56 : INV_X1 port map( A => n55, ZN => Y(10));
   U57 : AOI22_X1 port map( A1 => A(10), A2 => n170, B1 => B(10), B2 => n177, 
                           ZN => n55);
   U58 : BUF_X1 port map( A => SEL, Z => n169);
   U59 : BUF_X1 port map( A => SEL, Z => n168);
   U60 : BUF_X1 port map( A => SEL, Z => n167);
   U61 : INV_X1 port map( A => n41, ZN => Y(24));
   U62 : AOI22_X1 port map( A1 => A(24), A2 => n170, B1 => B(24), B2 => n173, 
                           ZN => n41);
   U63 : INV_X1 port map( A => n40, ZN => Y(25));
   U64 : AOI22_X1 port map( A1 => A(25), A2 => n171, B1 => B(25), B2 => n173, 
                           ZN => n40);
   U65 : INV_X1 port map( A => n39, ZN => Y(26));
   U66 : AOI22_X1 port map( A1 => A(26), A2 => n170, B1 => B(26), B2 => n173, 
                           ZN => n39);
   U67 : INV_X1 port map( A => n38, ZN => Y(27));
   U68 : AOI22_X1 port map( A1 => A(27), A2 => n171, B1 => B(27), B2 => n172, 
                           ZN => n38);
   U69 : INV_X1 port map( A => n37, ZN => Y(28));
   U70 : AOI22_X1 port map( A1 => A(28), A2 => n170, B1 => B(28), B2 => n172, 
                           ZN => n37);
   U71 : INV_X1 port map( A => n36, ZN => Y(29));
   U72 : AOI22_X1 port map( A1 => A(29), A2 => n171, B1 => B(29), B2 => n172, 
                           ZN => n36);
   U73 : INV_X1 port map( A => n35, ZN => Y(30));
   U74 : AOI22_X1 port map( A1 => A(30), A2 => n170, B1 => B(30), B2 => n172, 
                           ZN => n35);
   U75 : INV_X1 port map( A => n34, ZN => Y(31));
   U76 : AOI22_X1 port map( A1 => A(31), A2 => n171, B1 => n179, B2 => B(31), 
                           ZN => n34);
   U77 : INV_X1 port map( A => n63, ZN => Y(2));
   U78 : AOI22_X1 port map( A1 => A(2), A2 => n170, B1 => B(2), B2 => n179, ZN 
                           => n63);

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_generic_M8_N8_F8_DATA_BIT32.all;

entity ATU_M8_N8_F8 is

   port( CWP : in std_logic_vector (6 downto 0);  ADDR_WR_i, ADDR_RD1_i, 
         ADDR_RD2_i : in std_logic_vector (4 downto 0);  ADDR_WR_o, ADDR_RD1_o,
         ADDR_RD2_o : out std_logic_vector (7 downto 0));

end ATU_M8_N8_F8;

architecture SYN_beh of ATU_M8_N8_F8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal ADDR_WR_o_6_port, ADDR_WR_o_5_port, ADDR_WR_o_4_port, 
      ADDR_WR_o_3_port, ADDR_RD1_o_6_port, ADDR_RD1_o_5_port, ADDR_RD1_o_4_port
      , ADDR_RD1_o_3_port, ADDR_RD2_o_6_port, ADDR_RD2_o_5_port, 
      ADDR_RD2_o_4_port, ADDR_RD2_o_3_port, N5, N6, N7, N8, N13, N14, N15, N16,
      N21, N22, N23, N24, add_73_n4, add_73_carry_2_port, add_73_carry_3_port, 
      add_73_carry_4_port, add_73_carry_5_port, add_62_n4, add_62_carry_2_port,
      add_62_carry_3_port, add_62_carry_4_port, add_62_carry_5_port, add_51_n4,
      add_51_carry_2_port, add_51_carry_3_port, add_51_carry_4_port, 
      add_51_carry_5_port, ADDR_WR_o_0_port, ADDR_RD1_o_0_port, 
      ADDR_RD2_o_0_port, n1, n2, n3, n4, ADDR_WR_o_2_port, ADDR_RD1_o_2_port, 
      ADDR_RD2_o_2_port, ADDR_WR_o_1_port, ADDR_RD1_o_1_port, ADDR_RD2_o_1_port
      , ADDR_WR_o_7_port, ADDR_RD1_o_7_port, ADDR_RD2_o_7_port, n14_port, 
      n15_port, n16_port, n17, n18, n19, n20, n21_port, n22_port, n23_port, 
      n24_port, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   ADDR_WR_o <= ( ADDR_WR_o_7_port, ADDR_WR_o_6_port, ADDR_WR_o_5_port, 
      ADDR_WR_o_4_port, ADDR_WR_o_3_port, ADDR_WR_o_2_port, ADDR_WR_o_1_port, 
      ADDR_WR_o_0_port );
   ADDR_RD1_o <= ( ADDR_RD1_o_7_port, ADDR_RD1_o_6_port, ADDR_RD1_o_5_port, 
      ADDR_RD1_o_4_port, ADDR_RD1_o_3_port, ADDR_RD1_o_2_port, 
      ADDR_RD1_o_1_port, ADDR_RD1_o_0_port );
   ADDR_RD2_o <= ( ADDR_RD2_o_7_port, ADDR_RD2_o_6_port, ADDR_RD2_o_5_port, 
      ADDR_RD2_o_4_port, ADDR_RD2_o_3_port, ADDR_RD2_o_2_port, 
      ADDR_RD2_o_1_port, ADDR_RD2_o_0_port );
   
   add_73_U1_1 : FA_X1 port map( A => CWP(1), B => ADDR_RD2_i(1), CI => 
                           add_73_n4, CO => add_73_carry_2_port, S => N21);
   add_73_U1_2 : FA_X1 port map( A => CWP(2), B => ADDR_RD2_i(2), CI => 
                           add_73_carry_2_port, CO => add_73_carry_3_port, S =>
                           N22);
   add_73_U1_3 : FA_X1 port map( A => CWP(3), B => ADDR_RD2_i(3), CI => 
                           add_73_carry_3_port, CO => add_73_carry_4_port, S =>
                           N23);
   add_73_U1_4 : FA_X1 port map( A => CWP(4), B => ADDR_RD2_i(4), CI => 
                           add_73_carry_4_port, CO => add_73_carry_5_port, S =>
                           N24);
   add_62_U1_1 : FA_X1 port map( A => CWP(1), B => ADDR_RD1_i(1), CI => 
                           add_62_n4, CO => add_62_carry_2_port, S => N13);
   add_62_U1_2 : FA_X1 port map( A => CWP(2), B => ADDR_RD1_i(2), CI => 
                           add_62_carry_2_port, CO => add_62_carry_3_port, S =>
                           N14);
   add_62_U1_3 : FA_X1 port map( A => CWP(3), B => ADDR_RD1_i(3), CI => 
                           add_62_carry_3_port, CO => add_62_carry_4_port, S =>
                           N15);
   add_62_U1_4 : FA_X1 port map( A => CWP(4), B => ADDR_RD1_i(4), CI => 
                           add_62_carry_4_port, CO => add_62_carry_5_port, S =>
                           N16);
   add_51_U1_1 : FA_X1 port map( A => CWP(1), B => ADDR_WR_i(1), CI => 
                           add_51_n4, CO => add_51_carry_2_port, S => N5);
   add_51_U1_2 : FA_X1 port map( A => CWP(2), B => ADDR_WR_i(2), CI => 
                           add_51_carry_2_port, CO => add_51_carry_3_port, S =>
                           N6);
   add_51_U1_3 : FA_X1 port map( A => CWP(3), B => ADDR_WR_i(3), CI => 
                           add_51_carry_3_port, CO => add_51_carry_4_port, S =>
                           N7);
   add_51_U1_4 : FA_X1 port map( A => CWP(4), B => ADDR_WR_i(4), CI => 
                           add_51_carry_4_port, CO => add_51_carry_5_port, S =>
                           N8);
   U34 : XNOR2_X2 port map( A => ADDR_RD1_i(0), B => n33, ZN => 
                           ADDR_RD1_o_0_port);
   U50 : XOR2_X1 port map( A => n2, B => CWP(5), Z => n26);
   U51 : XOR2_X1 port map( A => n4, B => CWP(5), Z => n29);
   U52 : XOR2_X1 port map( A => n3, B => CWP(5), Z => n32);
   U2 : XNOR2_X1 port map( A => ADDR_RD2_i(0), B => n30, ZN => 
                           ADDR_RD2_o_0_port);
   U3 : NOR2_X1 port map( A1 => ADDR_WR_o_7_port, A2 => n23_port, ZN => 
                           ADDR_WR_o_6_port);
   U4 : AOI221_X1 port map( B1 => CWP(6), B2 => n2, C1 => add_51_carry_5_port, 
                           C2 => n24_port, A => n25, ZN => n23_port);
   U5 : NOR2_X1 port map( A1 => ADDR_WR_o_7_port, A2 => n26, ZN => 
                           ADDR_WR_o_5_port);
   U6 : NOR2_X1 port map( A1 => n1, A2 => CWP(6), ZN => n24_port);
   U7 : NOR2_X1 port map( A1 => ADDR_RD1_o_7_port, A2 => n31, ZN => 
                           ADDR_RD1_o_6_port);
   U8 : AOI221_X1 port map( B1 => CWP(6), B2 => n3, C1 => add_62_carry_5_port, 
                           C2 => n24_port, A => n25, ZN => n31);
   U9 : NOR2_X1 port map( A1 => ADDR_RD2_o_7_port, A2 => n28, ZN => 
                           ADDR_RD2_o_6_port);
   U10 : AOI221_X1 port map( B1 => CWP(6), B2 => n4, C1 => add_73_carry_5_port,
                           C2 => n24_port, A => n25, ZN => n28);
   U11 : NOR2_X1 port map( A1 => ADDR_RD1_o_7_port, A2 => n32, ZN => 
                           ADDR_RD1_o_5_port);
   U12 : NOR2_X1 port map( A1 => ADDR_RD2_o_7_port, A2 => n29, ZN => 
                           ADDR_RD2_o_5_port);
   U13 : AND2_X1 port map( A1 => CWP(6), A2 => n1, ZN => n25);
   U14 : AND2_X1 port map( A1 => N7, A2 => n15_port, ZN => ADDR_WR_o_3_port);
   U15 : AND2_X1 port map( A1 => N24, A2 => n19, ZN => ADDR_RD2_o_4_port);
   U16 : AND2_X1 port map( A1 => N16, A2 => n17, ZN => ADDR_RD1_o_4_port);
   U17 : AND2_X1 port map( A1 => N23, A2 => n19, ZN => ADDR_RD2_o_3_port);
   U18 : AND2_X1 port map( A1 => N15, A2 => n17, ZN => ADDR_RD1_o_3_port);
   U19 : INV_X1 port map( A => CWP(5), ZN => n1);
   U20 : AND2_X1 port map( A1 => N8, A2 => n15_port, ZN => ADDR_WR_o_4_port);
   U21 : INV_X1 port map( A => add_62_carry_5_port, ZN => n3);
   U22 : INV_X1 port map( A => add_73_carry_5_port, ZN => n4);
   U23 : INV_X1 port map( A => add_51_carry_5_port, ZN => n2);
   U24 : INV_X1 port map( A => n19, ZN => ADDR_RD2_o_7_port);
   U25 : INV_X1 port map( A => n17, ZN => ADDR_RD1_o_7_port);
   U26 : INV_X1 port map( A => n15_port, ZN => ADDR_WR_o_7_port);
   U27 : NAND2_X1 port map( A1 => CWP(0), A2 => n19, ZN => n30);
   U28 : INV_X1 port map( A => n18, ZN => ADDR_RD2_o_2_port);
   U29 : AOI22_X1 port map( A1 => ADDR_RD2_i(2), A2 => ADDR_RD2_o_7_port, B1 =>
                           N22, B2 => n19, ZN => n18);
   U30 : INV_X1 port map( A => n16_port, ZN => ADDR_RD1_o_2_port);
   U31 : AOI22_X1 port map( A1 => ADDR_RD1_i(2), A2 => ADDR_RD1_o_7_port, B1 =>
                           N14, B2 => n17, ZN => n16_port);
   U32 : XNOR2_X1 port map( A => ADDR_WR_i(0), B => n27, ZN => ADDR_WR_o_0_port
                           );
   U33 : NAND2_X1 port map( A1 => CWP(0), A2 => n15_port, ZN => n27);
   U35 : INV_X1 port map( A => n22_port, ZN => ADDR_RD2_o_1_port);
   U36 : AOI22_X1 port map( A1 => ADDR_RD2_i(1), A2 => ADDR_RD2_o_7_port, B1 =>
                           N21, B2 => n19, ZN => n22_port);
   U37 : INV_X1 port map( A => n21_port, ZN => ADDR_RD1_o_1_port);
   U38 : AOI22_X1 port map( A1 => ADDR_RD1_i(1), A2 => ADDR_RD1_o_7_port, B1 =>
                           N13, B2 => n17, ZN => n21_port);
   U39 : NAND2_X1 port map( A1 => CWP(0), A2 => n17, ZN => n33);
   U40 : INV_X1 port map( A => n20, ZN => ADDR_WR_o_1_port);
   U41 : AOI22_X1 port map( A1 => ADDR_WR_i(1), A2 => ADDR_WR_o_7_port, B1 => 
                           N5, B2 => n15_port, ZN => n20);
   U42 : AND2_X1 port map( A1 => CWP(0), A2 => ADDR_RD1_i(0), ZN => add_62_n4);
   U43 : AND2_X1 port map( A1 => ADDR_RD2_i(0), A2 => CWP(0), ZN => add_73_n4);
   U44 : AND2_X1 port map( A1 => CWP(0), A2 => ADDR_WR_i(0), ZN => add_51_n4);
   U45 : INV_X1 port map( A => n14_port, ZN => ADDR_WR_o_2_port);
   U46 : AOI22_X1 port map( A1 => ADDR_WR_i(2), A2 => ADDR_WR_o_7_port, B1 => 
                           N6, B2 => n15_port, ZN => n14_port);
   U47 : NAND2_X1 port map( A1 => ADDR_RD2_i(4), A2 => ADDR_RD2_i(3), ZN => n19
                           );
   U48 : NAND2_X1 port map( A1 => ADDR_RD1_i(4), A2 => ADDR_RD1_i(3), ZN => n17
                           );
   U49 : NAND2_X1 port map( A1 => ADDR_WR_i(4), A2 => ADDR_WR_i(3), ZN => 
                           n15_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_generic_M8_N8_F8_DATA_BIT32.all;

entity RML_M8_N8_F8 is

   port( CLK, RST, EN, CALL, RET : in std_logic;  BASE_ADDR : out 
         std_logic_vector (6 downto 0);  SPILL, FILL : out std_logic);

end RML_M8_N8_F8;

architecture SYN_beh of RML_M8_N8_F8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal FILL_port, N64, U3_U1_Z_4, n48, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, r126_carry_5_port, n13, SPILL_port, n141, n418, 
      n419, n422, n425, n426, n26, n29, n142, n17, n21, n22, n28, n33, n155, n1
      , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n18, n19,
      n20, n23, n24, n25, n27, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40
      , n42, n43, n44, n46, n47, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64_port, n65, n66, n67, n68, n69, n70, n71
      , n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, 
      n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n135, n136, n137, n138, n139, n140, n143, n144, n145, n146, n147, 
      n148, n151, n152, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287 : 
      std_logic;

begin
   SPILL <= SPILL_port;
   FILL <= FILL_port;
   
   r126_U1_4 : FA_X1 port map( A => U3_U1_Z_4, B => n43, CI => n13, CO => 
                           r126_carry_5_port, S => N64);
   U139 : NAND3_X1 port map( A1 => n17, A2 => n16, A3 => n63, ZN => n62);
   U140 : NAND3_X1 port map( A1 => n46, A2 => n35, A3 => n64_port, ZN => n72);
   U141 : XOR2_X1 port map( A => n34, B => n19, Z => n78);
   U142 : NAND3_X1 port map( A1 => n28, A2 => n90, A3 => n425, ZN => n89);
   U143 : NAND3_X1 port map( A1 => n97, A2 => n9, A3 => n22, ZN => n107);
   U144 : NAND3_X1 port map( A1 => n46, A2 => SPILL_port, A3 => n100, ZN => n94
                           );
   U145 : XOR2_X1 port map( A => r126_carry_5_port, B => n136, Z => n108);
   U146 : NAND3_X1 port map( A1 => n49, A2 => n46, A3 => n147, ZN => n88);
   U147 : NAND3_X1 port map( A1 => n147, A2 => n46, A3 => RET, ZN => n92);
   U148 : NAND3_X1 port map( A1 => EN, A2 => n44, A3 => RET, ZN => n148);
   CWP_reg_3_inst : DFF_X1 port map( D => n115, CK => CLK, Q => n155, QN => n11
                           );
   CWP_reg_0_inst : DFF_X1 port map( D => n118, CK => CLK, Q => n_2282, QN => 
                           n12);
   CWP_reg_1_inst : DFF_X1 port map( D => n117, CK => CLK, Q => n_2283, QN => 
                           n14);
   CANRESTORE_reg_1_inst : DFF_X1 port map( D => n130, CK => CLK, Q => n17, QN 
                           => n36);
   SWP_reg_0_inst : DFF_X1 port map( D => n124, CK => CLK, Q => n418, QN => n10
                           );
   CANSAVE_reg_1_inst : DFF_X1 port map( D => n128, CK => CLK, Q => n33, QN => 
                           n38);
   CANRESTORE_reg_2_inst : DFF_X1 port map( D => n132, CK => CLK, Q => n26, QN 
                           => n15);
   CWP_reg_2_inst : DFF_X1 port map( D => n116, CK => CLK, Q => n_2284, QN => 
                           n20);
   SWP_reg_3_inst : DFF_X1 port map( D => n125, CK => CLK, Q => n_2285, QN => 
                           n24);
   CWP_reg_4_inst : DFF_X1 port map( D => n114, CK => CLK, Q => n152, QN => n30
                           );
   SWP_reg_5_inst : DFF_X1 port map( D => n120, CK => CLK, Q => n29, QN => n31)
                           ;
   SWP_reg_6_inst : DFF_X1 port map( D => n119, CK => CLK, Q => n151, QN => n32
                           );
   CANSAVE_reg_0_inst : DFF_X1 port map( D => n129, CK => CLK, Q => n34, QN => 
                           n426);
   CANRESTORE_reg_0_inst : DFF_X1 port map( D => n131, CK => CLK, Q => n35, QN 
                           => n142);
   SWP_reg_1_inst : DFF_X1 port map( D => n123, CK => CLK, Q => n37, QN => n422
                           );
   CANSAVE_reg_2_inst : DFF_X1 port map( D => n127, CK => CLK, Q => n39, QN => 
                           n419);
   SWP_reg_2_inst : DFF_X1 port map( D => n122, CK => CLK, Q => n23, QN => n21)
                           ;
   SWP_reg_4_inst : DFF_X1 port map( D => n121, CK => CLK, Q => n_2286, QN => 
                           n22);
   CWP_reg_5_inst : DFF_X1 port map( D => n113, CK => CLK, Q => n40, QN => n425
                           );
   CWP_reg_6_inst : DFF_X1 port map( D => n126, CK => CLK, Q => n_2287, QN => 
                           n28);
   regFILL_reg : DFF_X1 port map( D => n134, CK => CLK, Q => FILL_port, QN => 
                           n141);
   regSPILL_reg : DFF_X1 port map( D => n133, CK => CLK, Q => SPILL_port, QN =>
                           n48);
   U3 : NAND2_X1 port map( A1 => n48, A2 => n141, ZN => n85);
   U4 : NOR3_X1 port map( A1 => n8, A2 => RST, A3 => SPILL_port, ZN => n97);
   U5 : INV_X1 port map( A => n143, ZN => n5);
   U6 : INV_X1 port map( A => n145, ZN => n4);
   U7 : INV_X1 port map( A => n64_port, ZN => n19);
   U8 : INV_X1 port map( A => n65, ZN => n16);
   U9 : OAI22_X1 port map( A1 => n85, A2 => n12, B1 => n44, B2 => n10, ZN => 
                           BASE_ADDR(0));
   U10 : OAI22_X1 port map( A1 => n85, A2 => n11, B1 => n44, B2 => n24, ZN => 
                           BASE_ADDR(3));
   U11 : INV_X1 port map( A => n85, ZN => n44);
   U12 : OAI221_X1 port map( B1 => n88, B2 => n3, C1 => n30, C2 => n147, A => 
                           n25, ZN => n114);
   U13 : NAND2_X1 port map( A1 => n4, A2 => n146, ZN => n74);
   U14 : NAND2_X1 port map( A1 => n5, A2 => n144, ZN => n145);
   U15 : NAND2_X1 port map( A1 => SPILL_port, A2 => n140, ZN => n143);
   U16 : INV_X1 port map( A => N64, ZN => n3);
   U17 : OAI21_X1 port map( B1 => n47, B2 => n84, A => n53, ZN => n147);
   U18 : OAI221_X1 port map( B1 => n94, B2 => n99, C1 => n10, C2 => n100, A => 
                           n101, ZN => n124);
   U19 : NOR2_X1 port map( A1 => n49, A2 => n52, ZN => n64_port);
   U20 : OAI22_X1 port map( A1 => n139, A2 => n20, B1 => n88, B2 => n104, ZN =>
                           n116);
   U21 : OAI22_X1 port map( A1 => n139, A2 => n14, B1 => n88, B2 => n103, ZN =>
                           n117);
   U22 : OAI22_X1 port map( A1 => n139, A2 => n12, B1 => n88, B2 => n99, ZN => 
                           n118);
   U23 : OAI22_X1 port map( A1 => n139, A2 => n11, B1 => n73, B2 => n88, ZN => 
                           n115);
   U24 : NAND2_X1 port map( A1 => n97, A2 => n10, ZN => n101);
   U25 : AOI21_X1 port map( B1 => n96, B2 => n97, A => n8, ZN => n106);
   U26 : OAI21_X1 port map( B1 => n92, B2 => n30, A => n147, ZN => n91);
   U27 : OAI21_X1 port map( B1 => n34, B2 => n19, A => n18, ZN => n79);
   U28 : INV_X1 port map( A => n76, ZN => n18);
   U29 : OAI21_X1 port map( B1 => n4, B2 => n146, A => n74, ZN => n104);
   U30 : OAI21_X1 port map( B1 => SPILL_port, B2 => n140, A => n143, ZN => n99)
                           ;
   U31 : OAI21_X1 port map( B1 => n5, B2 => n144, A => n145, ZN => n103);
   U32 : INV_X1 port map( A => n97, ZN => n7);
   U33 : NAND2_X1 port map( A1 => n18, A2 => n46, ZN => n65);
   U34 : INV_X1 port map( A => n84, ZN => n43);
   U35 : AND2_X1 port map( A1 => n92, A2 => n147, ZN => n139);
   U36 : OAI222_X1 port map( A1 => n93, A2 => n24, B1 => n94, B2 => n95, C1 => 
                           n96, C2 => n7, ZN => n125);
   U37 : AOI21_X1 port map( B1 => n97, B2 => n23, A => n98, ZN => n93);
   U38 : XNOR2_X1 port map( A => n73, B => n74, ZN => n95);
   U39 : INV_X1 port map( A => n100, ZN => n8);
   U40 : INV_X1 port map( A => n96, ZN => n9);
   U41 : NAND2_X1 port map( A1 => n18, A2 => n72, ZN => n67);
   U42 : INV_X1 port map( A => n90, ZN => n25);
   U43 : OAI22_X1 port map( A1 => n28, A2 => n85, B1 => n44, B2 => n32, ZN => 
                           BASE_ADDR(6));
   U44 : OAI22_X1 port map( A1 => n85, A2 => n14, B1 => n422, B2 => n44, ZN => 
                           BASE_ADDR(1));
   U45 : OAI22_X1 port map( A1 => n85, A2 => n20, B1 => n21, B2 => n44, ZN => 
                           BASE_ADDR(2));
   U46 : OAI22_X1 port map( A1 => n85, A2 => n30, B1 => n22, B2 => n44, ZN => 
                           BASE_ADDR(4));
   U47 : OAI22_X1 port map( A1 => n425, A2 => n85, B1 => n44, B2 => n31, ZN => 
                           BASE_ADDR(5));
   U48 : OAI222_X1 port map( A1 => n425, A2 => n27, B1 => n25, B2 => n40, C1 =>
                           n88, C2 => n108, ZN => n113);
   U49 : INV_X1 port map( A => n91, ZN => n27);
   U50 : OAI222_X1 port map( A1 => n94, A2 => n108, B1 => n29, B2 => n107, C1 
                           => n6, C2 => n31, ZN => n120);
   U51 : INV_X1 port map( A => n109, ZN => n6);
   U52 : OAI22_X1 port map( A1 => n48, A2 => n10, B1 => n84, B2 => n12, ZN => 
                           n140);
   U53 : OAI22_X1 port map( A1 => n48, A2 => n422, B1 => n84, B2 => n14, ZN => 
                           n144);
   U54 : NAND2_X1 port map( A1 => CALL, A2 => n44, ZN => n84);
   U55 : OAI221_X1 port map( B1 => n22, B2 => n106, C1 => n94, C2 => n3, A => 
                           n107, ZN => n121);
   U56 : OAI221_X1 port map( B1 => n110, B2 => n32, C1 => n87, C2 => n94, A => 
                           n111, ZN => n119);
   U57 : AOI21_X1 port map( B1 => n97, B2 => n29, A => n109, ZN => n110);
   U58 : OR3_X1 port map( A1 => n29, A2 => n151, A3 => n107, ZN => n111);
   U59 : OAI221_X1 port map( B1 => n28, B2 => n86, C1 => n87, C2 => n88, A => 
                           n89, ZN => n126);
   U60 : AOI21_X1 port map( B1 => n42, B2 => n40, A => n91, ZN => n86);
   U61 : INV_X1 port map( A => n92, ZN => n42);
   U62 : XNOR2_X1 port map( A => n112, B => n135, ZN => n87);
   U63 : OAI22_X1 port map( A1 => n48, A2 => n32, B1 => n28, B2 => n84, ZN => 
                           n112);
   U64 : NOR2_X1 port map( A1 => n136, A2 => n2, ZN => n135);
   U65 : INV_X1 port map( A => r126_carry_5_port, ZN => n2);
   U66 : OAI22_X1 port map( A1 => n48, A2 => n22, B1 => n84, B2 => n30, ZN => 
                           U3_U1_Z_4);
   U67 : NOR2_X1 port map( A1 => n73, A2 => n74, ZN => n13);
   U68 : OAI222_X1 port map( A1 => n422, A2 => n102, B1 => n37, B2 => n101, C1 
                           => n94, C2 => n103, ZN => n123);
   U69 : NOR3_X1 port map( A1 => n17, A2 => n26, A3 => n35, ZN => n52);
   U70 : AOI21_X1 port map( B1 => n43, B2 => n155, A => n60, ZN => n73);
   U71 : OAI22_X1 port map( A1 => n48, A2 => n21, B1 => n84, B2 => n20, ZN => 
                           n146);
   U72 : NOR3_X1 port map( A1 => n39, A2 => n33, A3 => n34, ZN => n57);
   U73 : NAND4_X1 port map( A1 => n422, A2 => n21, A3 => n10, A4 => n24, ZN => 
                           n96);
   U74 : OAI221_X1 port map( B1 => n21, B2 => n1, C1 => n94, C2 => n104, A => 
                           n105, ZN => n122);
   U75 : OR3_X1 port map( A1 => n37, A2 => n23, A3 => n101, ZN => n105);
   U76 : INV_X1 port map( A => n98, ZN => n1);
   U77 : OAI21_X1 port map( B1 => n137, B2 => n47, A => n46, ZN => n100);
   U78 : AOI211_X1 port map( C1 => n96, C2 => FILL_port, A => SPILL_port, B => 
                           n138, ZN => n137);
   U79 : AND3_X1 port map( A1 => n52, A2 => n141, A3 => RET, ZN => n138);
   U80 : AOI22_X1 port map( A1 => SPILL_port, A2 => n29, B1 => n40, B2 => n43, 
                           ZN => n136);
   U81 : AOI21_X1 port map( B1 => n83, B2 => EN, A => RST, ZN => n76);
   U82 : OAI22_X1 port map( A1 => n84, A2 => n57, B1 => n19, B2 => n85, ZN => 
                           n83);
   U83 : OAI22_X1 port map( A1 => n35, A2 => n36, B1 => n17, B2 => n64_port, ZN
                           => n66);
   U84 : AOI21_X1 port map( B1 => n418, B2 => n97, A => n8, ZN => n102);
   U85 : OAI21_X1 port map( B1 => n422, B2 => n7, A => n102, ZN => n98);
   U86 : NOR3_X1 port map( A1 => n35, A2 => RST, A3 => RET, ZN => n71);
   U87 : OAI21_X1 port map( B1 => n22, B2 => n7, A => n106, ZN => n109);
   U88 : NOR2_X1 port map( A1 => n24, A2 => n48, ZN => n60);
   U89 : OAI22_X1 port map( A1 => n68, A2 => n36, B1 => n65, B2 => n69, ZN => 
                           n130);
   U90 : NAND2_X1 port map( A1 => n70, A2 => n36, ZN => n69);
   U91 : NOR2_X1 port map( A1 => n71, A2 => n67, ZN => n68);
   U92 : OAI22_X1 port map( A1 => n142, A2 => RET, B1 => n35, B2 => n19, ZN => 
                           n70);
   U93 : OAI22_X1 port map( A1 => n142, A2 => n18, B1 => n35, B2 => n65, ZN => 
                           n131);
   U94 : OAI22_X1 port map( A1 => n426, A2 => n18, B1 => n34, B2 => n65, ZN => 
                           n129);
   U95 : OAI22_X1 port map( A1 => n75, A2 => n38, B1 => n76, B2 => n77, ZN => 
                           n128);
   U96 : AOI21_X1 port map( B1 => n78, B2 => n38, A => RST, ZN => n77);
   U97 : AOI21_X1 port map( B1 => n19, B2 => n34, A => n79, ZN => n75);
   U98 : NOR2_X1 port map( A1 => n92, A2 => n152, ZN => n90);
   U99 : NOR3_X1 port map( A1 => n64_port, A2 => n26, A3 => n142, ZN => n63);
   U100 : OAI21_X1 port map( B1 => n48, B2 => n55, A => n56, ZN => n133);
   U101 : NAND4_X1 port map( A1 => n57, A2 => n48, A3 => n55, A4 => n46, ZN => 
                           n56);
   U102 : NAND2_X1 port map( A1 => n46, A2 => n58, ZN => n55);
   U103 : OAI21_X1 port map( B1 => n59, B2 => n43, A => EN, ZN => n58);
   U104 : OAI21_X1 port map( B1 => n141, B2 => n50, A => n51, ZN => n134);
   U105 : NAND4_X1 port map( A1 => n52, A2 => n141, A3 => n50, A4 => n46, ZN =>
                           n51);
   U106 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => n50);
   U107 : NAND4_X1 port map( A1 => n9, A2 => EN, A3 => n48, A4 => FILL_port, ZN
                           => n54);
   U108 : OAI21_X1 port map( B1 => n419, B2 => n80, A => n81, ZN => n127);
   U109 : OAI21_X1 port map( B1 => n82, B2 => RST, A => n18, ZN => n81);
   U110 : AOI221_X1 port map( B1 => n33, B2 => n19, C1 => n38, C2 => n34, A => 
                           n79, ZN => n80);
   U111 : NOR4_X1 port map( A1 => n426, A2 => n39, A3 => n19, A4 => n38, ZN => 
                           n82);
   U112 : OAI21_X1 port map( B1 => n61, B2 => n15, A => n62, ZN => n132);
   U113 : AOI21_X1 port map( B1 => n66, B2 => n46, A => n67, ZN => n61);
   U114 : AND2_X1 port map( A1 => n46, A2 => n148, ZN => n53);
   U115 : AND4_X1 port map( A1 => n37, A2 => n23, A3 => n60, A4 => n418, ZN => 
                           n59);
   U116 : INV_X1 port map( A => RST, ZN => n46);
   U117 : INV_X1 port map( A => EN, ZN => n47);
   U118 : INV_X1 port map( A => RET, ZN => n49);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_generic_M8_N8_F8_DATA_BIT32.all;

entity WRF_generic_M8_N8_F8_DATA_BIT32 is

   port( CLK, RST, EN, RD1, RD2, WR, CALL, RET : in std_logic;  ADDR_WR, 
         ADDR_RD1, ADDR_RD2 : in std_logic_vector (4 downto 0);  DATA_IN_MEM, 
         DATA_IN : in std_logic_vector (31 downto 0);  SPILL, FILL : out 
         std_logic;  OUT_MEM, OUT1, OUT2 : out std_logic_vector (31 downto 0));

end WRF_generic_M8_N8_F8_DATA_BIT32;

architecture SYN_struct of WRF_generic_M8_N8_F8_DATA_BIT32 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component physicalRF_M8_N8_F8_DATA_BIT32
      port( CLK, RST, EN, RD1, RD2, WR : in std_logic;  ADDR_WR, ADDR_RD1, 
            ADDR_RD2 : in std_logic_vector (7 downto 0);  DATA_IN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component ATU_M8_N8_F8
      port( CWP : in std_logic_vector (6 downto 0);  ADDR_WR_i, ADDR_RD1_i, 
            ADDR_RD2_i : in std_logic_vector (4 downto 0);  ADDR_WR_o, 
            ADDR_RD1_o, ADDR_RD2_o : out std_logic_vector (7 downto 0));
   end component;
   
   component RML_M8_N8_F8
      port( CLK, RST, EN, CALL, RET : in std_logic;  BASE_ADDR : out 
            std_logic_vector (6 downto 0);  SPILL, FILL : out std_logic);
   end component;
   
   signal SPILL_port, FILL_port, OUT1_31_port, OUT1_30_port, OUT1_29_port, 
      OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, 
      OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, 
      OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, 
      OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, 
      OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, 
      OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port, intermediate_WR, 
      intermediate_RD1, intermediate_CWP_6_port, intermediate_CWP_5_port, 
      intermediate_CWP_4_port, intermediate_CWP_3_port, intermediate_CWP_2_port
      , intermediate_CWP_1_port, intermediate_CWP_0_port, 
      intermediate_ADDR_WR_o_7_port, intermediate_ADDR_WR_o_6_port, 
      intermediate_ADDR_WR_o_5_port, intermediate_ADDR_WR_o_4_port, 
      intermediate_ADDR_WR_o_3_port, intermediate_ADDR_WR_o_2_port, 
      intermediate_ADDR_WR_o_1_port, intermediate_ADDR_WR_o_0_port, 
      intermediate_ADDR_RD1_o_7_port, intermediate_ADDR_RD1_o_6_port, 
      intermediate_ADDR_RD1_o_5_port, intermediate_ADDR_RD1_o_4_port, 
      intermediate_ADDR_RD1_o_3_port, intermediate_ADDR_RD1_o_2_port, 
      intermediate_ADDR_RD1_o_1_port, intermediate_ADDR_RD1_o_0_port, 
      intermediate_ADDR_RD2_o_7_port, intermediate_ADDR_RD2_o_6_port, 
      intermediate_ADDR_RD2_o_5_port, intermediate_ADDR_RD2_o_4_port, 
      intermediate_ADDR_RD2_o_3_port, intermediate_ADDR_RD2_o_2_port, 
      intermediate_ADDR_RD2_o_1_port, intermediate_ADDR_RD2_o_0_port, 
      intermediate_DATA_IN_31_port, intermediate_DATA_IN_30_port, 
      intermediate_DATA_IN_29_port, intermediate_DATA_IN_28_port, 
      intermediate_DATA_IN_27_port, intermediate_DATA_IN_26_port, 
      intermediate_DATA_IN_25_port, intermediate_DATA_IN_24_port, 
      intermediate_DATA_IN_23_port, intermediate_DATA_IN_22_port, 
      intermediate_DATA_IN_21_port, intermediate_DATA_IN_20_port, 
      intermediate_DATA_IN_19_port, intermediate_DATA_IN_18_port, 
      intermediate_DATA_IN_17_port, intermediate_DATA_IN_16_port, 
      intermediate_DATA_IN_15_port, intermediate_DATA_IN_14_port, 
      intermediate_DATA_IN_13_port, intermediate_DATA_IN_12_port, 
      intermediate_DATA_IN_11_port, intermediate_DATA_IN_10_port, 
      intermediate_DATA_IN_9_port, intermediate_DATA_IN_8_port, 
      intermediate_DATA_IN_7_port, intermediate_DATA_IN_6_port, 
      intermediate_DATA_IN_5_port, intermediate_DATA_IN_4_port, 
      intermediate_DATA_IN_3_port, intermediate_DATA_IN_2_port, 
      intermediate_DATA_IN_1_port, intermediate_DATA_IN_0_port, n5 : std_logic;

begin
   SPILL <= SPILL_port;
   FILL <= FILL_port;
   OUT_MEM <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   
   REG_MGMT_LOGIC : RML_M8_N8_F8 port map( CLK => CLK, RST => RST, EN => EN, 
                           CALL => CALL, RET => RET, BASE_ADDR(6) => 
                           intermediate_CWP_6_port, BASE_ADDR(5) => 
                           intermediate_CWP_5_port, BASE_ADDR(4) => 
                           intermediate_CWP_4_port, BASE_ADDR(3) => 
                           intermediate_CWP_3_port, BASE_ADDR(2) => 
                           intermediate_CWP_2_port, BASE_ADDR(1) => 
                           intermediate_CWP_1_port, BASE_ADDR(0) => 
                           intermediate_CWP_0_port, SPILL => SPILL_port, FILL 
                           => FILL_port);
   ADDR_TRANSLATION_UNIT : ATU_M8_N8_F8 port map( CWP(6) => 
                           intermediate_CWP_6_port, CWP(5) => 
                           intermediate_CWP_5_port, CWP(4) => 
                           intermediate_CWP_4_port, CWP(3) => 
                           intermediate_CWP_3_port, CWP(2) => 
                           intermediate_CWP_2_port, CWP(1) => 
                           intermediate_CWP_1_port, CWP(0) => 
                           intermediate_CWP_0_port, ADDR_WR_i(4) => ADDR_WR(4),
                           ADDR_WR_i(3) => ADDR_WR(3), ADDR_WR_i(2) => 
                           ADDR_WR(2), ADDR_WR_i(1) => ADDR_WR(1), ADDR_WR_i(0)
                           => ADDR_WR(0), ADDR_RD1_i(4) => ADDR_RD1(4), 
                           ADDR_RD1_i(3) => ADDR_RD1(3), ADDR_RD1_i(2) => 
                           ADDR_RD1(2), ADDR_RD1_i(1) => ADDR_RD1(1), 
                           ADDR_RD1_i(0) => ADDR_RD1(0), ADDR_RD2_i(4) => 
                           ADDR_RD2(4), ADDR_RD2_i(3) => ADDR_RD2(3), 
                           ADDR_RD2_i(2) => ADDR_RD2(2), ADDR_RD2_i(1) => 
                           ADDR_RD2(1), ADDR_RD2_i(0) => ADDR_RD2(0), 
                           ADDR_WR_o(7) => intermediate_ADDR_WR_o_7_port, 
                           ADDR_WR_o(6) => intermediate_ADDR_WR_o_6_port, 
                           ADDR_WR_o(5) => intermediate_ADDR_WR_o_5_port, 
                           ADDR_WR_o(4) => intermediate_ADDR_WR_o_4_port, 
                           ADDR_WR_o(3) => intermediate_ADDR_WR_o_3_port, 
                           ADDR_WR_o(2) => intermediate_ADDR_WR_o_2_port, 
                           ADDR_WR_o(1) => intermediate_ADDR_WR_o_1_port, 
                           ADDR_WR_o(0) => intermediate_ADDR_WR_o_0_port, 
                           ADDR_RD1_o(7) => intermediate_ADDR_RD1_o_7_port, 
                           ADDR_RD1_o(6) => intermediate_ADDR_RD1_o_6_port, 
                           ADDR_RD1_o(5) => intermediate_ADDR_RD1_o_5_port, 
                           ADDR_RD1_o(4) => intermediate_ADDR_RD1_o_4_port, 
                           ADDR_RD1_o(3) => intermediate_ADDR_RD1_o_3_port, 
                           ADDR_RD1_o(2) => intermediate_ADDR_RD1_o_2_port, 
                           ADDR_RD1_o(1) => intermediate_ADDR_RD1_o_1_port, 
                           ADDR_RD1_o(0) => intermediate_ADDR_RD1_o_0_port, 
                           ADDR_RD2_o(7) => intermediate_ADDR_RD2_o_7_port, 
                           ADDR_RD2_o(6) => intermediate_ADDR_RD2_o_6_port, 
                           ADDR_RD2_o(5) => intermediate_ADDR_RD2_o_5_port, 
                           ADDR_RD2_o(4) => intermediate_ADDR_RD2_o_4_port, 
                           ADDR_RD2_o(3) => intermediate_ADDR_RD2_o_3_port, 
                           ADDR_RD2_o(2) => intermediate_ADDR_RD2_o_2_port, 
                           ADDR_RD2_o(1) => intermediate_ADDR_RD2_o_1_port, 
                           ADDR_RD2_o(0) => intermediate_ADDR_RD2_o_0_port);
   MUX21 : MUX21_GENERIC_NBIT32 port map( A(31) => DATA_IN(31), A(30) => 
                           DATA_IN(30), A(29) => DATA_IN(29), A(28) => 
                           DATA_IN(28), A(27) => DATA_IN(27), A(26) => 
                           DATA_IN(26), A(25) => DATA_IN(25), A(24) => 
                           DATA_IN(24), A(23) => DATA_IN(23), A(22) => 
                           DATA_IN(22), A(21) => DATA_IN(21), A(20) => 
                           DATA_IN(20), A(19) => DATA_IN(19), A(18) => 
                           DATA_IN(18), A(17) => DATA_IN(17), A(16) => 
                           DATA_IN(16), A(15) => DATA_IN(15), A(14) => 
                           DATA_IN(14), A(13) => DATA_IN(13), A(12) => 
                           DATA_IN(12), A(11) => DATA_IN(11), A(10) => 
                           DATA_IN(10), A(9) => DATA_IN(9), A(8) => DATA_IN(8),
                           A(7) => DATA_IN(7), A(6) => DATA_IN(6), A(5) => 
                           DATA_IN(5), A(4) => DATA_IN(4), A(3) => DATA_IN(3), 
                           A(2) => DATA_IN(2), A(1) => DATA_IN(1), A(0) => 
                           DATA_IN(0), B(31) => DATA_IN_MEM(31), B(30) => 
                           DATA_IN_MEM(30), B(29) => DATA_IN_MEM(29), B(28) => 
                           DATA_IN_MEM(28), B(27) => DATA_IN_MEM(27), B(26) => 
                           DATA_IN_MEM(26), B(25) => DATA_IN_MEM(25), B(24) => 
                           DATA_IN_MEM(24), B(23) => DATA_IN_MEM(23), B(22) => 
                           DATA_IN_MEM(22), B(21) => DATA_IN_MEM(21), B(20) => 
                           DATA_IN_MEM(20), B(19) => DATA_IN_MEM(19), B(18) => 
                           DATA_IN_MEM(18), B(17) => DATA_IN_MEM(17), B(16) => 
                           DATA_IN_MEM(16), B(15) => DATA_IN_MEM(15), B(14) => 
                           DATA_IN_MEM(14), B(13) => DATA_IN_MEM(13), B(12) => 
                           DATA_IN_MEM(12), B(11) => DATA_IN_MEM(11), B(10) => 
                           DATA_IN_MEM(10), B(9) => DATA_IN_MEM(9), B(8) => 
                           DATA_IN_MEM(8), B(7) => DATA_IN_MEM(7), B(6) => 
                           DATA_IN_MEM(6), B(5) => DATA_IN_MEM(5), B(4) => 
                           DATA_IN_MEM(4), B(3) => DATA_IN_MEM(3), B(2) => 
                           DATA_IN_MEM(2), B(1) => DATA_IN_MEM(1), B(0) => 
                           DATA_IN_MEM(0), SEL => FILL_port, Y(31) => 
                           intermediate_DATA_IN_31_port, Y(30) => 
                           intermediate_DATA_IN_30_port, Y(29) => 
                           intermediate_DATA_IN_29_port, Y(28) => 
                           intermediate_DATA_IN_28_port, Y(27) => 
                           intermediate_DATA_IN_27_port, Y(26) => 
                           intermediate_DATA_IN_26_port, Y(25) => 
                           intermediate_DATA_IN_25_port, Y(24) => 
                           intermediate_DATA_IN_24_port, Y(23) => 
                           intermediate_DATA_IN_23_port, Y(22) => 
                           intermediate_DATA_IN_22_port, Y(21) => 
                           intermediate_DATA_IN_21_port, Y(20) => 
                           intermediate_DATA_IN_20_port, Y(19) => 
                           intermediate_DATA_IN_19_port, Y(18) => 
                           intermediate_DATA_IN_18_port, Y(17) => 
                           intermediate_DATA_IN_17_port, Y(16) => 
                           intermediate_DATA_IN_16_port, Y(15) => 
                           intermediate_DATA_IN_15_port, Y(14) => 
                           intermediate_DATA_IN_14_port, Y(13) => 
                           intermediate_DATA_IN_13_port, Y(12) => 
                           intermediate_DATA_IN_12_port, Y(11) => 
                           intermediate_DATA_IN_11_port, Y(10) => 
                           intermediate_DATA_IN_10_port, Y(9) => 
                           intermediate_DATA_IN_9_port, Y(8) => 
                           intermediate_DATA_IN_8_port, Y(7) => 
                           intermediate_DATA_IN_7_port, Y(6) => 
                           intermediate_DATA_IN_6_port, Y(5) => 
                           intermediate_DATA_IN_5_port, Y(4) => 
                           intermediate_DATA_IN_4_port, Y(3) => 
                           intermediate_DATA_IN_3_port, Y(2) => 
                           intermediate_DATA_IN_2_port, Y(1) => 
                           intermediate_DATA_IN_1_port, Y(0) => 
                           intermediate_DATA_IN_0_port);
   PHYSICAL_REGFILE : physicalRF_M8_N8_F8_DATA_BIT32 port map( CLK => CLK, RST 
                           => RST, EN => EN, RD1 => intermediate_RD1, RD2 => 
                           RD2, WR => intermediate_WR, ADDR_WR(7) => 
                           intermediate_ADDR_WR_o_7_port, ADDR_WR(6) => 
                           intermediate_ADDR_WR_o_6_port, ADDR_WR(5) => 
                           intermediate_ADDR_WR_o_5_port, ADDR_WR(4) => 
                           intermediate_ADDR_WR_o_4_port, ADDR_WR(3) => 
                           intermediate_ADDR_WR_o_3_port, ADDR_WR(2) => 
                           intermediate_ADDR_WR_o_2_port, ADDR_WR(1) => 
                           intermediate_ADDR_WR_o_1_port, ADDR_WR(0) => 
                           intermediate_ADDR_WR_o_0_port, ADDR_RD1(7) => 
                           intermediate_ADDR_RD1_o_7_port, ADDR_RD1(6) => 
                           intermediate_ADDR_RD1_o_6_port, ADDR_RD1(5) => 
                           intermediate_ADDR_RD1_o_5_port, ADDR_RD1(4) => 
                           intermediate_ADDR_RD1_o_4_port, ADDR_RD1(3) => 
                           intermediate_ADDR_RD1_o_3_port, ADDR_RD1(2) => 
                           intermediate_ADDR_RD1_o_2_port, ADDR_RD1(1) => 
                           intermediate_ADDR_RD1_o_1_port, ADDR_RD1(0) => 
                           intermediate_ADDR_RD1_o_0_port, ADDR_RD2(7) => 
                           intermediate_ADDR_RD2_o_7_port, ADDR_RD2(6) => 
                           intermediate_ADDR_RD2_o_6_port, ADDR_RD2(5) => 
                           intermediate_ADDR_RD2_o_5_port, ADDR_RD2(4) => 
                           intermediate_ADDR_RD2_o_4_port, ADDR_RD2(3) => 
                           intermediate_ADDR_RD2_o_3_port, ADDR_RD2(2) => 
                           intermediate_ADDR_RD2_o_2_port, ADDR_RD2(1) => 
                           intermediate_ADDR_RD2_o_1_port, ADDR_RD2(0) => 
                           intermediate_ADDR_RD2_o_0_port, DATA_IN(31) => 
                           intermediate_DATA_IN_31_port, DATA_IN(30) => 
                           intermediate_DATA_IN_30_port, DATA_IN(29) => 
                           intermediate_DATA_IN_29_port, DATA_IN(28) => 
                           intermediate_DATA_IN_28_port, DATA_IN(27) => 
                           intermediate_DATA_IN_27_port, DATA_IN(26) => 
                           intermediate_DATA_IN_26_port, DATA_IN(25) => 
                           intermediate_DATA_IN_25_port, DATA_IN(24) => 
                           intermediate_DATA_IN_24_port, DATA_IN(23) => 
                           intermediate_DATA_IN_23_port, DATA_IN(22) => 
                           intermediate_DATA_IN_22_port, DATA_IN(21) => 
                           intermediate_DATA_IN_21_port, DATA_IN(20) => 
                           intermediate_DATA_IN_20_port, DATA_IN(19) => 
                           intermediate_DATA_IN_19_port, DATA_IN(18) => 
                           intermediate_DATA_IN_18_port, DATA_IN(17) => 
                           intermediate_DATA_IN_17_port, DATA_IN(16) => 
                           intermediate_DATA_IN_16_port, DATA_IN(15) => 
                           intermediate_DATA_IN_15_port, DATA_IN(14) => 
                           intermediate_DATA_IN_14_port, DATA_IN(13) => 
                           intermediate_DATA_IN_13_port, DATA_IN(12) => 
                           intermediate_DATA_IN_12_port, DATA_IN(11) => 
                           intermediate_DATA_IN_11_port, DATA_IN(10) => 
                           intermediate_DATA_IN_10_port, DATA_IN(9) => 
                           intermediate_DATA_IN_9_port, DATA_IN(8) => 
                           intermediate_DATA_IN_8_port, DATA_IN(7) => 
                           intermediate_DATA_IN_7_port, DATA_IN(6) => 
                           intermediate_DATA_IN_6_port, DATA_IN(5) => 
                           intermediate_DATA_IN_5_port, DATA_IN(4) => 
                           intermediate_DATA_IN_4_port, DATA_IN(3) => 
                           intermediate_DATA_IN_3_port, DATA_IN(2) => 
                           intermediate_DATA_IN_2_port, DATA_IN(1) => 
                           intermediate_DATA_IN_1_port, DATA_IN(0) => 
                           intermediate_DATA_IN_0_port, OUT1(31) => 
                           OUT1_31_port, OUT1(30) => OUT1_30_port, OUT1(29) => 
                           OUT1_29_port, OUT1(28) => OUT1_28_port, OUT1(27) => 
                           OUT1_27_port, OUT1(26) => OUT1_26_port, OUT1(25) => 
                           OUT1_25_port, OUT1(24) => OUT1_24_port, OUT1(23) => 
                           OUT1_23_port, OUT1(22) => OUT1_22_port, OUT1(21) => 
                           OUT1_21_port, OUT1(20) => OUT1_20_port, OUT1(19) => 
                           OUT1_19_port, OUT1(18) => OUT1_18_port, OUT1(17) => 
                           OUT1_17_port, OUT1(16) => OUT1_16_port, OUT1(15) => 
                           OUT1_15_port, OUT1(14) => OUT1_14_port, OUT1(13) => 
                           OUT1_13_port, OUT1(12) => OUT1_12_port, OUT1(11) => 
                           OUT1_11_port, OUT1(10) => OUT1_10_port, OUT1(9) => 
                           OUT1_9_port, OUT1(8) => OUT1_8_port, OUT1(7) => 
                           OUT1_7_port, OUT1(6) => OUT1_6_port, OUT1(5) => 
                           OUT1_5_port, OUT1(4) => OUT1_4_port, OUT1(3) => 
                           OUT1_3_port, OUT1(2) => OUT1_2_port, OUT1(1) => 
                           OUT1_1_port, OUT1(0) => OUT1_0_port, OUT2(31) => 
                           OUT2(31), OUT2(30) => OUT2(30), OUT2(29) => OUT2(29)
                           , OUT2(28) => OUT2(28), OUT2(27) => OUT2(27), 
                           OUT2(26) => OUT2(26), OUT2(25) => OUT2(25), OUT2(24)
                           => OUT2(24), OUT2(23) => OUT2(23), OUT2(22) => 
                           OUT2(22), OUT2(21) => OUT2(21), OUT2(20) => OUT2(20)
                           , OUT2(19) => OUT2(19), OUT2(18) => OUT2(18), 
                           OUT2(17) => OUT2(17), OUT2(16) => OUT2(16), OUT2(15)
                           => OUT2(15), OUT2(14) => OUT2(14), OUT2(13) => 
                           OUT2(13), OUT2(12) => OUT2(12), OUT2(11) => OUT2(11)
                           , OUT2(10) => OUT2(10), OUT2(9) => OUT2(9), OUT2(8) 
                           => OUT2(8), OUT2(7) => OUT2(7), OUT2(6) => OUT2(6), 
                           OUT2(5) => OUT2(5), OUT2(4) => OUT2(4), OUT2(3) => 
                           OUT2(3), OUT2(2) => OUT2(2), OUT2(1) => OUT2(1), 
                           OUT2(0) => OUT2(0));
   U13 : NOR2_X1 port map( A1 => SPILL_port, A2 => n5, ZN => intermediate_WR);
   U14 : NOR2_X1 port map( A1 => FILL_port, A2 => WR, ZN => n5);
   U15 : OR2_X1 port map( A1 => RD1, A2 => SPILL_port, ZN => intermediate_RD1);

end SYN_struct;
